PK   �n�X���e"  ��    cirkitFile.json�]ێ�F��C�y���_�m<�쌍��,����(�v��zU�i{���~�F�R��*���c?�.1��0�dd3����P���_m����q�p?{��|��8l?�_�|�i�:>�~8�>����/�?}*�CYl�Tg����u.����Y�7v�X���RJ��_����y�~��Z��VZ�A��VF�A��VV�A��VN�A��V^�A��VA�A��VQ�A��VI�A��VY�A�@>J�(+������aq(�w�V������~�	��v��m>~z�/�7J�]����vᲊ�T�r�+�ή��_�(}�Ӯ D A�r�/� r�/� r�/�PܤbA*+#��|�C��!� �DA3L�"� r�/� ��|�m�WA,�WA,�WA,�WA,�SA,�SA,侳1v�V7_ �}��Nc�i,;����X�A�i,;R?�vk;(;�e�Vk;����ƲS+������Nc٩����cme����*`m�����Xvj���X�A�i,;�JX�%���4��Ze��2�vPv�N�ި#� ��?���������px���(X~̏�^��)X~̏W���*X~̏׻��+X~̏W���,X~̏	��-X~̏�7��.X~̏f��/X~̏�����������p��������e|���$�p�a���X~̏�N���?��4�o� �`�i0?ޮ�8����`~��l?p�����x��~���Ow𻠍�|nE��yc���إ���me��/?�H6�{`GV�ݼ:���ӑ�o���m	Y���#���Y�vK���{GV�݄8V6R�	u���el}��Z_w��/�^료����k}�0��P���c�K��P���c���ڜ>��P��c���ڄ=v���
�g��PV�?+ԟ��
�g���B�9���P��CQ�|\��J���Q.�~���]iy��sa��EX�����`9j��۵��6���[G�~,��=�	{��H/�^8"x����P�^8"x�����B����PA�� �_�/H����B����PQ��(�_�/
������QB�E���PI��$�_�/	����KB�%����}�PI��,�_�/�����B�e���PY��,}!/~#/}%����������W���J�^^I_�+�y%}5��J�/I�(^����+D�%"��x�H�J���DZ�N��EZ�R��KEZ�V���E���"U���jQ�C �-���[X���2d��>ir�KQ��Vrȝ�N�,����.ԮL����&,��F�mܭ#o�����=[\��ܹ�Y���yP���>���dWP�0��5*h�>�l/���d�m4�(֋X���Nѝ��^l\��슭s/4�����}P���ަ�Jj���K�(�!���"������^�����'�o���g���f�/�(��t#Pu*:��:#�T���a��O�0U��c�����1�@@�I�F ���u#P}
;�EVH�|��s���_J9�7
�>��	�5�y���C�A�`�[�8
�>��	��5̉�����A�`~���8
�>�	7��M�a~���8
�>C�	��̏�����A�`~���8
�>{�	��̏�!��h��|8j�� �}J;Ƶ}f;h�)��r�X��<8*ЮSpm���9!pT�]���> c���C�@�N��}8<����Q�v��k��x�n����:����ܞCG�u
���1�=��
��\ۇ�c,p{�h�)�����	�Z纃��m��,Ҷ]E]�]��]����H�NzM¶�{<,Ҷӄ_���8����4!�$l;���"m;M6	ێ���H�N�M¶��|<,Ҷӄc���8P���4!�$l;���"m;MX6	ێ���ȕ�i��&a�qH?i�i�I�v���E�v�%�i����xX�m���&a�q�?i�i�I�v$��"m;M\6	ێ�xX�m���&aۑL ���4q�$l;�a���&.�`�S���Nh�i�֙� #��"�t���r�����CPzv_�=D�ҳ�y����]�c�R�����{�Fu �b����X�~�>��Qp�Mca0��lh,F�}猅�`����Z�Qq߷!ca0*��c,F�}�9�u1*�[�T�b�Q�Ũ�bTl1*�[��F��bg�#��0�;
�Q�è�U*v�TZS��}��X��F��b�Q���b����aT�1��c|�Ǩ�cT0*��F��� z?�Qq��8`T0*�G��#F���QqĨ8�^�aT1*�'��F�	��Qq¨8aT�0*N���'��3F���Qqƨ8cT�1*�g��3h���Z�P�uZ�P��Z�P��Z�P��Z�P =Ö�@zF-�V�PKy��<�bj5��Z�Ӡ=Z�Ӡ%=Z�ӠE=Z�Ӡe==`]o`Z
 J���eh� J�e����i^���l//M� ��j�k�e�͛�2��� (�Zwh2 J�.��ű�V�/�������R+ ���
F �:���N� a�S+@����
F �:���N� a�S+@����
F �Sj���ym�ۆ�ms�(�Sj'���0�B:�V�p��os�(�Sj'��0'�B:�V�p��q��(�Sj'��7��q��(�Sj'�70?�B:�V�p��q��(�Sj'�70?އH��F�?��v�V@�¸v�V@��:׎�
��fA��:׎�
��eA��:׎�
��dA��:׎�
��cA��:׎�
��bA��:׎�
��aA��:׎�
��`A��:׎�
��_A��:׎�
��4W;Yf?M�5	ۮ�
pX�m'
������
�H�NzM¶+�i�i¯I�v�V��"m;M6	ۮ�
pX�m�	�&aەZ���4��$l�R+�a���&��mWj8,Ҷӄd���J� �E�v��l�]��ȕ�i�I�v�V��"m;M\6	ۮ�
pX�m'Z�&.k'+��"m;M\6	ۮ�
pX�m���&aەZ���4q�$l�R+�a���&.��mWj8,Ҷ��e���J� �E�v��l�]��H�N�b;���c?+����{�.�g���S&!(=��Ǟ�A�٩;��!��@�Ũ��#��0��}j5�����`4����X���>����}�2��oC��`T���X����s;�bTl1*���F��b�Q�Ũ�bTl1*�;��F��b�cT�0*v;��F��b�Q�Ǩ�cT�1*����b�Q�Ǩ�cT�1*��F���Qq ����8`T0*G��#F���QqĨ8bTA��0*�G��F�	��Qq¨8aT�0*N'��b��F���Qqƨ8cT�1*�g��3F���Z� -{(к�-|(�ʇ-}(�ڇ-~(��-(��a�x =��P+y��<�Zj1���Z���iЂ���iВ���iТ���iв���74���U�N� Gy����
r�W{���
r�W{���
r�W�;8�(�S+�Q�O�˜����j�p�pX�?�ބ����P>�>��r��߯��0{���dݯAX|�������Q��=T�"�7���~*��g�"�pu�/:�]���'�H�\��/:T["����X-}x������n��?�ݞ���فʏ� ^�o���[b�����ر������/�5ܼ�Bo&0����A��aK䂓)SHG���o�5vJ�=�I����#��b�I�O����u�?�v��8���~Hl��91D��N�BQ'��C�I�,�u�:!1D��N�BQ'��C�I�,�u�9!1D�lN�BqJ0'u[�����BZo�۴����V7������1N��< .W|��EN�#��p�r�S�8)�'� W,�8%��N� 3Yp�r�S28)�l� ܫ��M��^���1N�ݤ< �Z�r�S7)�?5 ��"L��G^}d��#A��#)b?,��l��m�ވÃ�˯#՚�y['4�� ����H�&|��)�8<����:R�	��u�"b?,��i��m���Ã�˯#��y['&�� ����Hy&|�֩�8<����:R�	��u�!b?,��f��.: i'��x[_z�/�ǘ���xT�K�پ���#0îd@@���	�aW�1  Ɔ�̰+�cCt�fؕ;��!:R3������v�bl��X��r~16DG-`�]�������0î^@@��q
�aW�.  Ɔ�t���r����v��bl��S��rl16D�)`�]������0î�Y@@��q
�aWn,  Ɔ�8����=�Z ���KI-�bxcᷣ��9[k�����[�NG�om�9��~ks�����[�!�2*���|8�<=)�T��/U�H5���c,�T���/�Hu��:a,�T�����}�T���c�JloV Ub{{�X ���ǎiR%Z��xX�*�J�h�J�R%Z��T�V�D'U��*�u|�wf���^I��Iu�:u�=F	^l�%	�T�N�b/U����K����S/t�:�R���K��JR%��T�A�� Ub��R%��T�A��(Ub�*1J��J�R%F�����T�Q��(Ub�*1I���JLR%&��T�I��$~)Ub�*1K���J�R%f��T�Y��,Ub�*1�_��ߊ�_�+�{q%~1��oƕ�ո�W��J�v\�_�+�&K5bM�k�5���z�|�F�b#_���h���h���h���h�ҍ~q�fh��W����;�E4�p��
�:عn����zl?8�а�Ѓ�I�t�����|CÌ=8�P��N9$���u��ԯ��2�]��|�5>�!�C�������w$n_n��~d���E�2UA.Y������Kk.����
�k�a*l�a����k�a����kX�a����p�5,װ\�r�5,�p\�q�����lq�5�p\�q�5��\�s�5<���Cs�5<��\�s��5�\#p��5Be'��F��kD��F��kD��F�L�5"׈\#q��5�H\#q��5�HUkp��52��\#s��52��\#s��5rՀuVMX����q�G�#��|]��+ǣ�U+��r���_խP+��@��Z�
jT:Е���Sխ��+1�J���_���-�R�!�������9޳d^�ו�s��ީ�c?����<rw^�E�i�~o�y��ڣC7�_%YV{lXF�?�}�ś�V��� e�Ȳ՞�%N��^��H�������>C���4�N���"���r�GN�xW��;v�m�:�sy�����o�%۾�N�\��?]��K�t)�/�ӥؾ�N�R��:]R�K�tI󜱸�[5���=����Gn�A��|B��O�*ۼ�+jťˍ���Y��}������X�~�~����<�%O���I�����
䤗9��b������*fK�,�o�d6S�i�[�2�+��E�Q�н޹T��{� ����X�A�g4?��hД|>{8�	��Y��>~�ܕ�g{��Y��K���m2n���ϑ�w�T1e��6-�a.��R{.p2��b4%����x��ʅer���g����24j^�K&�lu]�eP�����2���iQť�R�&���n}a݉��gTj�h�\��b�p9X�r6��֌�m6�6ВvK[ݵ�nɄ��,G��meCEC'RM�{��U���u��j��u�j�#�e
d�x�{6�,&*߰Q\Ҵ=����$��k��b�l��2{�%���~i����O~��~�|��[>%�0��l
�����	�z*Gd�s��ߪ��]ڤSn�/����+��м����n�DŏF����4Ԗ�5�����vv��u���.-#y�l�(�,�L����)�\�$�C�:�.��|�l��2jj�SEj3}�|����U:y՚�b�;���*���v>4��������8,���_U,8�T��O���^�������Y+4
ў�U�y\ +���47J�[��.����2Y8���O�M2o�7��PI"'�]1(�z�S�7�2�{�J��(����s��z~���I&����'��\_/U ���$zvz��놟�<�u��䅔�:�L��Ϸo^V���Tpv�_S�_��!g�sW���;x��iG}�֧!�$CgN�4�R
�@MI�tϊ��4�����s�:V61���$�29K׸޸"7�n<����CK<MO*��e䮘/�ȿ��J�RdҰ�e���| �h|���Ԃd��f�EOR��P<���x<��+�v�~I��ף. O���<�c�O�����!��\�W�cN�3��L*{6y����S�B�&=��Ȕ���c��g��Z�k��Ix��ZbJ��6�YnP���}�ZZC}�T+�#��1j��ӝ��,#�g��i�Ι��S3�Р��A��ԍ,��ΟP����y�>4�3�6�C0Vl2�bA�k�b��"E�>��i�C�*{�Oh��f���OO��gS�Ԭ�F�xn���Z������ ��xv/g��!_{�Ց�����G���C�ݎ���4��g�T�m&�5�D�fIb}nr�.���ץ�	�?/��3%z���%'��m����y:�OC�uD��UCe�8C�J���(E^��h�EB43���խ���m^���yq�M@|��Q*��j܊zW ��F�ш����ۑ�x[���hx'��]Ӥ�Vu���scUw1�f@�F�K���Rdz�.��{$��z�}��,�-O�oh�|��Ul�4�Z=�e&�u+���V�Kst�"}��}��n���
���gք\���������L��à���4�e���/�i�f��^[�r9�\���f�D�������Ő���I����.���]_�M�!�i�k��r���udR۬mha�eh�Ǥ'��
�U��6�Ǩ����j�Ir><���A��{�`�y�scpE���<��WHW�tG��W�^E�M�l��W�z*�6��i�Kcb�Fh�䨡}�z��S�:��#�}�|�\�4&�G��{;�T��ZB5b��gE��"39BIW �8g��݋�]d�|���R4���mb�ޑ{Y f[�5�yRM��͛��濍�4q�<�k>����N�NJj�@�{�u�J��ˤ�lM=ä1�RS/��	*��j>)yc�j��<'>��SӐ���n�����z|���߲�H8K;�e���!=�֜�=?'�S ���+�X�4�Y��7��P����Ҥ�L�va3�ϐ���W>O�Z�{4���yv�Y��4��7�q [�x��<�im4h�n��Ȼ.=���.<On�K�9�:F�K3����MΝ94�Sn׮4�.|\�.m5=�:/v;�^�슲Z�|�<��*�'86ς|�X��.���%�ۗ<�h�_ɺ˥v�/i���O��6-�|<��?����o�:����{���O���?臧������{������?��ͮ�{,��cy���q��+�;����?�d��ᩤf�X�?����P^��؅����ǯ���<<}��� N7�-Y��� 4g���v��)d+�Z����ba�IM�Zl���\���VR⠅�J�)��1��E����L}�\O�/��_��}�h���><�����Q�Ұ��ԥ-��oZ������_��᭚g�h2�3�ȁ��թ�=ܕ�[B�y����B�R���������X�!����Ȥ�O�W����U��~��&Blu�??}\�����}�uq�}|��m��+�n��a��o�p���H���\���F)��i9�uQ���H�U�4�윋���� ���1l����p��W�r4��|U����tn���lAq?�����j��~�4�s�N?}�o������\}(�g!CT/rm���Ǜ�?]���b��~�����<�������ĕZ~Gֿ{8���y7���F�w��;r��������mu鋷�T`���E�a;f*�C���Hj���8v������
��w���x�����|����ȿ�y���	dCP+��r�yU*��l�,UM�Ɩ�Y�M������B�����:P>j�|��q�G��v#�s���m+�;
-�=rG1���?���ۍPư]b8e���A��%ʸ��V�vv�p�͇��ԍ0��Z�a��o^�ϗ��{AB�m~�i��w���^��#n�^V��H�Uqťisg���q�K6M���_��r�7+�r���	{ls���Ԧ��o&�ź[��R��3�a�Jq�1��5b�/i�˾��g^�64ۓb���;��|��ʵ�ڥ���wƗpg0l:1p����@�w�!;��۫����u�2�Tc��u��R_<q�s:k��ȍv,��c��{��>伻�J7�lOpcԕ8��)��kU�Ū�z�=Z=��������}/��T�k�Ӑ�!�b������}��Sq,���'A=V�������*�~������O��E���������qs�:������PK   �m�X�l����	 ��	 /   images/50cc3d53-9c96-4f8d-a7da-648aea826718.pngl�g4^��u!J��]�Dt3J�!�ѻ����^"D�]���$���e����w�u?�g����k�o{�ki�H�鉱��HU���`a�aaa�<!�O�3֘������êc���l��屰~�?������\��<���{���^�����he�k�	v�wU���d�i����n�d��b����.e���.%�������?$!*��ea����?6R1����z�Py/��k�}O��i�U�{���y�*r>Z	HgT�bN|���M[�g��A7	`B.`�l5 8~�I�泭7E4ou8�����>������(]����4�Y<��8ķ�-_ �n���!�c�;;!����_]�}����oB��z����ׅ��a�w.�wǑ�[,�	5Y]^�Y��/Wn�>��u��<`�E�;>L���U��F�p=�y���ߦ]��혎��~����(8��kr�������<�A��އ�&��o��o�ܮ1�C���d�w� ��5��(p�J��l��P��ڼ��}o��Ǆ������>*4�� ��.r#�6�>n�Av��H�6�����I(�j2\�4�x��<�k
A^�Ս�c��!�Mۏ�R�0s��+�v���sEs��RR6���	���wk�k�%ߙ۝�BUq���H���Y����>|8��6�� �9�],���.�2=�ʳ?�X9����5"� 0U���Y3���e: �R��;0
���9��G��ŻȪ͊N��B�p���P!�B$3��JP28���Q]��l�Q����6�g��0Ӯ�]�xNaB�!��m�X�?�0�0�c�D��V6�<����R|b���ƪ�oq2��2(6~5��|�}MF�h\�����=�.����ɿ!KhR�#x	C�j��;:��ÒB��d#we+�X��d��i[�nW��,����q3iRa��=��G�+>è��Ȩ`�%���[�~�d'����i��і��r���;,!;`nN�1�j49�V5�1Ts'��W=s.�9ʲn����<H@��:s[{7���6����
 #A�i��I�5nN><��:�[eV"�*l
�Z;(R�I�A���g+-��"��!�?>0��s�,l|�C,3ː�/%ᑮ�?��t�c��|D�<�"E�'��!����7ϧ�
9�~c���S1N��i_��cb$l.�Rރ(���TN����W��j��fm��t8VT�{�vDA#lMFBل�K���D����~|�5���4j�s���N���͠��&QAe��д��G�����V(@��&�~"��T8�* ��ɽ��K�Z��(:���X�qHM����3��?i��\F��Ÿ�o�X��y	gՃ7I����2Xw�$��
�A��42Eå�RN�%0٢�Ea{U���M`HsL&n�aK/|�����k"n���Km�Y��2�HY��$0��Z��n�.T�?^s�V��8��f+��Y�M �݉ �c`C���ć��E~��{+��`���"���8ɲ�f�v�U���!���Q=�ӯ��ͯk5(��]��1-�������
�7�CZ[��^�>��7��1$��q�N�Z��ĝ�[���Ҹ������~M�n�כܩo���~�����q���"f̊�K�eg���#+�5�B7m�䁯��)i{��M�
�Mq�ތ��ے��ǃ�'F�A15��M�jװx�b|�{I�h���)]��_Z�����v��#�r؎L��Kɥݣ�Kt�mv_߭~�ߍy��M*��\���ʚBM�~<c��I��Ge�y�JvU��v�'�ZR����[��m��ea�o������	aH��߶t4�<Ȍ�w:�SG3~`,�ʻ�1��'gi�-�����h{8��r��5RL@{
Dk^��L;_|�*��p�����D5��ON�6�JD4��ЅYT�]ME����`�)kԠ����Dժ���72���x�]�M��v����vb���3I�k��D�\3�{zo�I�(��c�I�=1��N#nFZst�u$�"�N���lMss�J/��\7Ȫm�R�X;�7�M��wL��n��!�6�}�GD
|�G��*��%����5r@ �Kuq�Uvf�"t��O�.���4�=+�NGH8YL���1:���#�P��g�NMa��KsR^�4m�I���a@�[��4�6R��*S�C�uW�>���Z���A+�Ӥ��VB��}<ٻ��i��SH��A>��3���"�?�vp��6�6(�HW}�-�ID�{�O�G��H��$�oI�3[��t�a���)���&4%�t񔯜a�(bt����M��������Ql����yQ��
��
����#����#|����OC�ɒveO�;��&��i] �"��8��y�bk1����ʿ=tn�y��"�I-���m����y�e�q�ʜY;�����AShө)����\
O� .��Ǻ�V��_�j1���S�`Т�y5?/`� 9o*�Р��y��ު���b�M�#46�/ڜm[�~�b�U0��oc�ƻ�d�#���	����m���e��)9�\���ㆽ	v�m�a��������t&���7P�Pk/E��J�|iz�8�|�>Xz�^�;��c�a�_�{�BP#���!ZW�y@�7�t*��ʅ�v(�q斥���VN)��̋D1{܂��5=Y��k:��	�k��k���P��X�fbb��U)��7���e�B5�1[3���:y��I�#��sOX�ZĪ�{���Y��TL�KO}��6�upb5�D���/m!/�M��Q�w�v�@/��)�ھ�n߆]!�Uo�9�va���
S��H5���Lh�����p��R��(��/����8��hrė'��/��~�������oO�ߔ�Ęm8>ߵ:� ��P������8�=w6��m��� >(�����t�ې�/94~f�L�qE� e3����x
+ǖ2��i���!���,�;h����f;���I�a}��Կ&�<Uf���s�VX���c��.�L3��u��
ú(�'�cT~*c�ƶ26Z�-��W� ��g�^����'�d��6z��_�z��\�8 �\7�C��
�^f�scPQ�Ez��@�o���� r��? 2^�����H�UwZ8M6W���%�O*y���n�.��s	����*�����q˴���q/�uj��Ѳ����1ۋ��~^3��y)�>��6UXNI`�}7���J�Ě4��f5�Ov�eE��K,�1gg�G�y"��tw|� b�u��`�~${��Y�����c�&��ګk����/���
��Z��-*0�8W�����K���xv�SvE<��}�Q4���S�s!�OV�e0(o.i{�������Y���#c1�Z��̃�b��#:�)�R��X2�c�o��tɣ5���Uy�)��H�F
Z��5#)�tq�|��`\eq3��s��Mns��o8]��[OV���n#�F���{#���2T�����?xԪp�S���F� ��'���R�u����C� :�T�<w�{��lm���e���$G{����Û�*�/1ƾ�Mbï�RLs>�#�w\X@L�>�.42�xd?-fm�,�A�3��é��A|�Q�jv���5D4̂qx�
gH�T���n���h��F�;�j����φt�ٍ2��<ʷ�A���:痰���r�Mau��f�O��Ny,\\\�ϫ`����D�u��Ś�T���9���;"��v�f%jp���̀�i�uZ�4�'u)o�3މ&F��'�U�e].9kx��W-���ۅ���n%�<z��q�jH�{�i���3���Y>GF픘}����� &��2dC��� U��vQ���B����K����9��Hz��P|k1���~.:��,R�=B�q
R0�:�[i"�r�՗e��7�͌�t�����%m9�4�y��0�d�	�A�m��+��e؟����U��J��#�Sr/�������M�U�B��s��<�15ft�Wa�"���縷v�2��X�aT����� �z�W*��dG����ۋ��H
��א��E�ޡ�1û����2�C�Q�`8�����I�\��pZܦ�o�h?�Y��
GU
G��$���~*u��h08gvFJB�yS�����!\�v"��r|����}٧����%��f{y�+���ց�x��%b������0a	d��F�"9Z��^"OJ���xL�B��"��9�H��Ll�9�xP|5�8:p,�L��zZc8N�����S�#.$��?&'����V�-5ej�x�� �{h��@����T�Ѯ�Jc�+u�X����-����HM����8�!ɳ=�&6�#�HS1�f�hX)��?h��zM��?�jw~'bET��fB�z=h��,�F�������Sܴ4F�@X%,��ǋΙodZ�c�n"M��8߹ɧ\qGE�͒�o�$��w��M��[�OXߙT'Z��ǳ�LY�y��H��~Q�E��Tw!>���fb 8�?*o
��L'I�lO��l�����L�pX�q�D`f�/u<��2������+���>� *�����Ǚ�aZ�H ���w�0��"�� vq\n�~�^3���.��g��_��Ү��M�%EF��㶐+*lbBث���j��Wgϭ�駄W�J��:Ädo64#~̒����W}z4��������^��R� /���bL��H�)�+i�^���1|�����z���*�{���k?��ޒB)�/ ��l�_������dEſ=KN�5	��j�:�Q�l�y���/F��o�BĪįԮ��㸶�&E��3F�gBm�`�"l�1�-R?��,E��h�	ؼb:%����n�ʪ��^ӕ��[CfGea����e������I8�[uV���q�4���$^� ��6M�fxR(�|yj��28���TOME��^�Q�E�ܬi�*G؝�+-v��-��S��@����JF�jJ�'e:����eln�c�&[3�퓂 �8~�%g�0�޿D�k�+c�S�+;�	l&ׂf�� t��b�7��2��`�
�b;W�?|ɪ�2{��L��A=���u�_�3J�uU���9j|Ϙ�1�5O11�F?D4�1���'�����:j}�������_���@W4��5܎>b���l�3]&-L��Dg�y��mAluG�9���z�Y1nfuɗNG���7\�o
	RO�_��U��6W:c�e'2�?5�, �"�Ke0ЩJ�e������9[�MS���|7wg�g�����+f��ieJ=MF�c�3+#n�,�;|�N�%s�����b�Zg֭l�=��.b�?�Ty���,aj������^�	�ɸ�]2��y87�!�a6�\�B��$�I��N�z�Z���N{R��V}?�<~�����=�Ӣ��da��N�b���+n�TA\/������|���<���X��_)E���z!=�tvp�!��h���Ɓ/'�N�;�s*XW_ i����/E1ؓ��C�E"��yw�o)6+"n�+A��<�;��Ԛ�7d���j��M�p\R� t�|��u���֍�F!�����w[��MG��ŉu`��	^��\�����������@��VL�AU��2���ܯ�c�B&�*Pd�OQb���K�T�­ʦ,�MNo�"ީ'v�l��ַ���K����Ub�y���Z�$6���0�xSv������SoL�|��Y��zѤ�A��<�S6Sp���e��WbAKukq�cves���`�U��U-�� %)�<9���?��^���-����k�ZD;[��J�����}��0}���ga:��DfX郎�j��,df���n�8����ñ4وi������V���KBL������Bݯʃrf2)ȗ�]�V/F�,N�@&�&iWS-i�	z?�4������Z���F9P�/O��Q�3��g?�����:W�F<&]
�/����6�๡�5
(��&{����Y	ۜ[?h�v�h�9Q%�p4󒩤'�PXDȔ�k��ӑa��;znq� I�գwq�J���o�n��}J`^�C��|�b�B������4�J�������2��͉�Ҍ��c������])�[ՔJ�$�Jfe��^ʃ���k@b���j6İ��K�-�`�}�c4�Fa#;�^��Z�&,|�ru*x����<���ұ���ӑ���V��-AŜ	̱��T5Jv<�7O�!����iJ�V!�VbH�w}���[=�b��3���FD'k�	wpb����HZ���?L�1��W9��Dj~�Q����o��
���/'tdg�ݽ��f�<E� �F۰�E�~�&�-��8Fv��A.���bĂf2&Q�ڞ9����Qդ9􋤮i�L� �h�����2s92����l�"�p��@ ˚}���A�AQf;[dpQ�3�}b�U���k/G)�0��<�̩��%B�H��9�{s�¦_R�����Y�cM����������ɋd
����i�U��4�*B�#���tt��S~��-g���pr�a�W6���|I�Z}~LZ�8{�F�rǯi@�;�;�"=4T�~� ���h�������^3��3cH�)k�!��������ݛM��@&�B��l�����V�0�CC}	
wm�GE0��E%���Z|z�P<,H��vj�&Ͱһ1����{�����P�dɍҌl��������������G$��<!Q�K!��n��3}x�;�(�T}2R� d�)� U@6c�Bh�U}��|x�k'�Ҥ��kM�����I���qWuK��	�wH�6��J̛S�En��)4A�*f�QI�������J�Ef�g/�h8�Wl��[�.�w�%����r)eXYl8e*��G���'�|�.d��8Fa[���]zV`=����|�K�$<�.Ň]�7�*�*��ޤ��a*n��w�`go��������	w��+��~\L�q:v�O�5Ŏ�����c>���s�P���O_z7x��U���-U��>����Ϲy\?W��,x�a#�ݱ���%���Y+��;ط���h&>��dUޘ4�k/T�	8Q�]�I���䴓F��w)p�u�<QC����"�A��5d��q���7X��z6�b�2�O>L#�	}�&53�"x&�[
,��s�(�		+Q�iJ�^�K;K�Q��`W�EѺ�9bE�o�Y�԰Ǻ��*`ᔿ+�^k��e���Yi�G	�fk�x�|䬣K[�e#I�zܡ�B�.�&�Pl$�}��c2�Q�PdK����\T�b�65�����@���Tr;k����2����_?�Bo}B��9Up|���c�7�urD>����Լ�o�]���i��RiƔ�k��&�}�Qݠ]���'����oh	��^u�[����9Pd]��c��?���/]~X�Œ
OmdI�����!�����_1�55VM���"~V��rQ��A�)i�?����CS7&�v\EJ�({��^�H٦Yn؆;F�O����z�&�Ӕ0hȓ�sr�FI%�����`N����Ա{-I#�������Ń1�P�T ?㯼��q2 ��ɬ#;;AH��&��C�1ܫ�N���UqE6(^����(�˽?����xމ2�w�!�˨B�g$�z�s9i݆qEP�A�U��7S/��/{�kipY�[{���y�zb����w�6��R���eLh���v��-��vJ�!B�!�oO��MCǚP{a�a���S`/�XQ�TsK�F>�k}��NE��>�geW2�f��PR��Y�K֘�uS'{G��ߨeG��p;�@��r{X����_��O����� {J�a���-.�RGGU��Ⰹ�����`|�	X��ӻ�V��ɭS�3��^�9.K�����6�D_ߏ�Ӏa�MC(��Ti�n��Y�ʳvJK���^^^�1Yϲ�,����&Ы�%!�|������s�������@d��ˣ�^�G�����(��iRe�險\2���A�B�q�B������0�i���	�K���4_�24�2��\�´)�L��vhDuE#��G���! 2h��v�u�M��Cg��k���S�Ut�)��\�y�<�����w�c���~o^���K��?Q8W09fn���\,�=�\��)io.%7���'dpϚ?��t)�t�����cd�k�*���T4}���	��C��&��-xbiz�f{���Q\�iWP���-?LVc��ڧ�0h'��ڜ���g�����J���a`�|UY����NU#�YD�!{5��B�\��;�sc1V�N����֊Aֵ��:�����'������L�@;�BJ�ƾ>3#0"M+�z֙ܽ|@�ԊW�{���=%zO�H�]^Y�[r~���� �^�����*��J�kʢ��'�l�o e�绉�XZklf�_��.�"#Xc8���J��X�=�PpE,Ӓ ����N'�t�I�G&�W��9����x�Ω �����&9$���_vpB��塺|kc�c��c8e�Ʉ~�:j�3�������(�%�����v�-�WOǇ�kOrù-0�u���FG�M/G�g��F
̀�%�������W� ��ǆ�7Q$�۸�^��~�oV�{����|=0��^�Q�H7��3DD�p�5��C
��:�q�m��0�����`�&�4�M>�F4|sg����*�G*J L��Q�	:E���FI�|��*���K`�$�7� 7f4nANjlP����
cZ�t�ˠ�q�PO�����5Ӳ4�"Ǖ��q�J�D~}��_�1�_���t�'��L!��Ĺs�E
��-d�+���	��ː�])����x�v�T�ڐ��~$���|�5����uc�u��Ҝ�Kwy�>ݧ"|�{zth��%�n����p���b�y[!B�׹7���������/���ײ����n.�䦻MM��k�'���ut��]�;b��Ǝ?�{�1=C�ٔ�p%���P_Ao�O�ז>
���P�*��JPҜDPnݯ��m��O�5�CΦ�o��(i�m�d�)�$���A9��z����O��])�poÚ�<�M�7�y�+חuV&dl'>�GDA��&�2P"K7W�D�w!D��U�;Mhq����ʔ��I]�����)	&��òr���8�������ʭ;��) ��
������h2��$z�MD�4�_�ј�p��9���U�%w����<��n�s�M������ߗ��{=�e��YKF�,G��s����e-�����U=�T� �D!���ٵ�K�iΥR�Ź>��c 9l�����ٔ�'��ˏ-��?�}>y�Qh�r�FIB(�\v����o�leeu*�9��n�E(�c'dX[�,L���q���?��FV�q�����`��?e�{�lԜa��UBu!���:�-��v:5Ѡr>�,A�P��s_tS�~�$r>��A�C�-�d�*3h+��A�i�Pk�J��B�X�V��ʏ.��ա����mY�l��U�,��9�!���	��z������%yG���3�\U|k��&3:`֑yjr`�-��f��Vگ�����0yE��B�����{��K,!����h�2���%Sj!���gW�Ej<��P�����+�"��y'H2����Ձ� ���� ���hU�%������F�?)_��,����'?K���x�ڣwN�F�HpB��*��E�]|�'M�*_/�J��5V"�f�
bb
>��9�#��Z�����%HmcJ�����V��=ƙ�eA��2j����ɬ�A8�9n�r޼�*�	��/q��oK�e���{ZhQy,��S�Bn�o�F�_�޴�T����dQ�[|�4�%�N����[A�����␬yj̼+�+8u!�M����K�ڋ#H2��dsq��խ����$kmtrv��G=;[�7�͎$���ԑw�Tĩn���f��:��QҬ�N䵉*�8O=�����7dFRm��"�GE�7&�-I�h#ç�Q�������n3�7�D�� ���V���$�D]qX�x;;�h�3���r�!(��N@&�3S��Z���3Bq)���,~������R�+�X��`$R3{�Ar(+^q�Q��z�f��b�����Z ���e����6眖�}��ȟif���:4~����Ψq�iN�u��g��g,�k�A�̵�c���ڙ�x�X62E�j�=ԕ���U�����	  �����M�%:T,ٰ����U��
�"~K���b$&m�T���B�ӹ������������f�Wى;�_M�-Pʦf=����"��s,�#�Cӝ�20ỉv��z!K��:�{>�Ji�*��R��������h?�$��*Y���k5� �(��J6�Pc�ͩ�"wP#UQ
���gh�3����|�!{��������9d��m��:k��O�p���w��=gN��\U`i/�T/?z�8��|֏��Z��V=]"r�Y%1�g_ըj��^��~)ŉ1�=�Q�D�߄4����#�Fabj^@�����k�ɧ����ET�k�U ��.��*��G)Y{.�Ow�m�G=�*A��Pw*���nS�F6�����{.��l�)���3,��i_��:,eG9K��/� ��7#Hu�E��9�'����i�~ntM��#=��"�q1���,�������T/��7R��e�������5M�4U��T�]���2���j4�bY7�K8,bmq��
����oc李����4f[���8f#�[ݯ�m��{���&4F���~�K�N����Γt7� ��S��y���G[���e_���7j�H�� zT�����c^)ct �]8!���u�ɝ~�ӎ���G`i_7h�Y09D�|�rg8�J�=�o������b��C�G�:9�F�7!��Ƶa7z�x��9$<	���Q���YW2藙��y9��J/�n� �#�U�׻��z!C�;���>M�8 �%�`���o�7�g��0I�V���i
@sn#�j���[�n䀛��C���-R��'����K �jM�J�B��IЗ�Z@��"sҫ�Oa�u(-_lڗZK��'���Xk��-����L+3!B���eK�e������2ݗx#VR�!�RCE*ŪH�5=��7��mD��ė��[W;N��\�;	'U�A�L����2^�����%�tҀk�k��]�7�1��㝱���B���U�>?	̦��0�N��2�[����|�_ͭd0V��S[����s�<p
�Ș������r�7jL*H:^J#_�4��;nf��<d=��f�)����-m��ڋ�q�����*hZ����R�Y��JZ�1@9�PN��w~��=*79�ծ"��B��ɗck�ZdwJy��Ks�S�r��t�|�1�7�@V+@[��f�ȠЧ��i�+��S�Վ�R �t��X�c~�����7�Q�|��q�����|�~��Ýߠ$6��~[{:
���qb�нd|��b�0�/� ����t�^y�����Z#%F�dS��5�DF���ގ/]-����EYN	d�E.*ѧ��<�5dy*�.�'N}�[���-yw9X8(����K*�� N>1��݌�"#�C��Pt�%o�̃Y�ŧ*���Z�rd���<�@��Bj�&�&~t��a˗��>�׌�bf�~?ܙw���qi0^�`c\�>k+��O$�G���dX���d�\�(t�<u�V����{�i�{�r�w�) �D�����S���"殢�"�Pxq�cc�H��H���/���b��X�)�&�^�I�zq�����}!�.��J�H�I*�1GYV�v�?�
�����r�]fQ3vy�c��Tn���҄e�t:on�0{W��2����[�EN�}P���N�%���C0�F���KP	�{�3�4�3Ǒ�x�����dӸ���/�^���_��l�$b�<]�G�!pJ���^J[�)��s�)�n{j���	�J=����BBK�O�E���ǀ�D�Xl�jj���w���Xul0j~�s���5Qg�g��=���s���N���D�[��_/6���m��|�Xz�N��~-�	j���t�iw�Z��zeʘ�;c&~H�����d�{3�aʚ��rW"����i��[�q�!��D"~a�M�_�FH����82>e�Oh0��W���Y�=�o��ffJ��Q ,MLV�+6��A���am��H(Є� ������
��#0Z�^�g���QǬ�"���E���T�;�O3��,��	 P��h*�ު����]�Y�!�N���]1�����ck}��Yڞ��=�����QX��홨]3�^7s�,�Ԇ���� ��E&?��%$?i}m�st�q��!L�\���wԌ�����M��e�X[�Q�{f���91��VC��c��-���*�,�N�OQ�5��ߍ�;O�Tg�$��;*x�ݍ�����*�M�Duw։���Ul��*Tb�7�y��&��[�"7,IAT�o�{g\$�TY�cO<&(�;QP��qF��U�G�u�����+JU���r�2�4;��<�>Fo�o����<�R��$�Ʀ=*а�Қ�٪�"K�{n��h["D�Hg�x��Q*�Cø���bIS������rx]L�f�kC�ƻ�������,���1{>���ə�[��ME8W=:��O��T�����z7���4�8<�����O�m�� )xK��k�{�$A{����_Su|{�,�����x��`4u̺�;k �*D�H��.����I$�$���(]�ǖE�NC����mz#�%y��w d1vp�a����(��������C�24�+}/K�}�t����*����A^�z���g��V�<���ޏ�&���;��FsGa�%����y�:�u�#�R���S���G�_H6a���?�RYp�I�
w7��DW#ϟ�ˎ˰�����q��#��7�~v�\)'����#���������-�Wk��·2��_��v	Q1��������b�ℵyWski>��_�i�my$)��I�����z}i:��3�R��oW�rBI2���nf�G�i���0��I-��~�q�!�Od&�aenUs���1�^*^ol���$b�&����Ŗ�戳���#����[���Ĥ���1}^{w&��C_!�u�ڬ�)�m��W��	eL���7{��#><hI�3��t��B��޸5����c�S¿����ߚ���賫a��{�� �Ď�c�j�8������h�f��1�LX��a�@5���X�8���t��Tk�r_��CN���ޛ��0u^����cѩW�{�=�^i�T�@������'��B.۩�p��%�r��Gf�4s��8'�M3��������|�Rx�J�E���Kz�v��X�;ȎipL�"���*H��N9drv{�b�:�Ӳ G�S��/$b"�r�?�HzYb�m�J����*��k�e��}zʮ��I϶��@F	P�ݘ��k>�p�%� $h�i�}��r:UBͩ�}�r���������%����ZF����`�A�Vs�*��͊m�h���9AO��+ö��l�s�O�6���SmD���T,�ù��qU�k��(�!��~*���³
/KEToyIz� ���ǬK�,�c�d���d�6/���m��"���5FnqgSAه��ēiX|��/����uc�%�
o�_|5}�M����_V�Y7�������6��I~H�S�n���Zp��W�mޯ��������A�;��&b�>O���k:A$�Ek�>�(���������4���v��sE��E)>���&x� �"��D�s����l\�r�E/d�in��3�l���z�e�?)�b�39�Zi!=��KÊ8TN\+IQ�۩A�I�9�F^>mz�*����*8�]�Hè�f�^
A������q"��6dՍg��s�j�X �]��UP��Q��<d!_qU�Y���`�_��ݣ��d,�� ��Ǽ d�w�7&0�ڋj�]<�K����#q��?oN.V�h�e���̤��t݌�h����[7����T�>��rih�M����l����m����t�t���������|ٽ���Ug�4B	;ut��g~�a��
ڍμ_�zq,�Z�7�"H�Շ\ާDx/ͪ"�*l�[��-B��-�.V�0��q�Kȣ_�ϣJ��WГH���ܩ	bvHl>aޠ�+��~[ñ��<�ә���7v�2%�3y�M�D���'�����@*���V�T�J�֋N�e��qɣ�M��*�3���! s������٩���娢C���p��cr-x�M�_�X^�n��� 4�����e�ג`�ܻFt��4��M~�՞��������qL�?�?z�5�/��i� �H�V�z�9�Y�����WI����E	��e��>l)u��ڰd��ı�.���k�{̀hB]mF�K�Z���J�L�Bx�0�0-n�Nr#�Q�=�X%$^4�<[W5~�ܭ�1`��ae�nc����Yj���̋����Y]���J��C����?��ˢK�:c>�LJ:g>�lTJTK�O!�ษ��G����>5z��jo~8.aRIY�ǸgU��$7�2��{3:�>:Q�L�ٞ�3nW�U�_:�ٕ+��k���8��l?���4��pp
�Y�m�_O���$t�g�	y�/��5��,�/�LM�A􂖧ֳ�P�����A{�0Z��kWEϬ�=&� 5m���|ğz\x�� ��|�}����J!�o��>����PC��5	�M�͈ͭXV�ޫI��`�2H�y�����wQlkJ����7��p���gu2x�Y�dj����xJ�f:���9�~w�K��f�.��.��3f6�"����"�j�`��@�wjX��}����<	W��r�/�$z��׾����zU�<�#)Oi��mǒ�� ����WG��ǫ}uM�o��\��cju�׉�8�v�{��F�Ek)Ry�e=��ȑ,]߾��{*���5����Mi�,<38I6b�M�Kϲ�f$Rn|�tAU�Rf�I(�0�5��0M�X�۷2b����� ���¤����,{�s�Ll௮�f�R}��N43�8-�g�r�̶zW���q�M�*8ܶ���f�!Gv���c"4����٫M}�7qKb����T M��ӕ浢��h���4�IUoS��s��=�Cӿ���q�\�������.�s�t"|{h��C`#���xW𿩫�8Q��L��1ZE�s�}���HX�J��i�=�h�B�XA�j�[�[�=Q����q�e�����C�I���g�a�6
y^�FRQE@P�A�J���ۜGcT|���������B�|6��h�f����C��sĲa�a���֧7R�;o�Af{��	� �Ozq���6��ud�j�.l�'c�X]�Bl����ą���c͉��d�-,���i����h+�����f�D|�{}�l�:W s�V3��*�*���7>���9|�Cɩ]�^�4��M��"d~1��0���|����[ ��[X1N��~4q�jm$�Hy~iT�P�{S�Y%��a�i>~dr%>���^�ڣ��'���`x̝��k�R/�D'̬�K�u�m]m�����T�BT���!��{�c�mT_椣��ܗ�]=�bC���e-������v`��a�W�o��=5� ��>������XM��ޛ)σ�g�e��&�y���0�}D�U>�<��U<Vh�~so?,(sW~w9�2��Yoc�UqNJu�}{�q0�cKN���ۧ������}�ߓy��	9�ϵfM܏�^C[e��_u���e)e��}�g�z�*���d7	�;���-|"��9sQ�RMl�m��ʲ�������ޛv�,
���ld����ї���U�	��y,��5�+�喣��QM�4��)���W�Sm�w\��6�����R��/K����u1٢�����G�}��+6	�+��N�~1rDA[�1���r\�>�S�lG\�|�劉C�͟Ր�[�H�d�`��i��#�	�z�z�I�U:"E��%zZ�I���y�����&�'��U��Z�=,��ηw�Ƒ� �o͓�Mp\��k��Bic�|D�/�6��ӑ28�#{���y�D��͞�ӻV���=m)��m]��̵g�M������� (@׿ �U�PS��	���nGI�Ly��>J5��Z~{�-���m�8xT{���c�,/L{���� �:%��)K��!��8-cw�~��ȑ����7�������Y����a���|���\��?�_>�ݧ���yt�#6c�G0�g�F�����(�Xy�rz�_�Ż�o���7o�S'���`wYUK˥ܺ���O��/���?�cy��%p�`�\#��������Z&�,iXm����]����țߔr�9�!/��	�á%���Nl<(C}8R���H��X9�Ty��+��wo��'&ॊĽ��͖�>�W�����7���|w�qYZ�.�GJw�0���C�
����-�oF'��N�Ƒ�E�	:)�Ϟ%�^�z��2E��ć��O~�M��o>+� +e��\:rnXP?<,���9�������d�k��6ɝ�䟺-1t��f$�x�B�I'Qr�w�$hO�~�\��h�86_u�����ɳʨuk'�o��ߝ8�4���jn�O�P���T�����|N�����rn�<�2ku^�i���G'ݼNI����5��]�A���.�Ў��Ք�;N��$}`�9'�B����S�� ��o�y�\����K��IO7��<t#<H�ԋ���UoY�x�ڐځX�x{�,x�}uu��O�%�:���.��}p|���7��?���P.�?Z�aA�jH����l~�|s�V�쳯�_�*O�Υ��\C�C���#��ƍk�G?y/ב1�ڐ�������_T������/?+/^�D��m�A��Q_f�[A�W�
G+ݐ&6���2,_���,@o��l�x����?������JEFz�f
��I��ֵ�Y��c���l�ײ��Mr��3���B��_ �RϩG\����q:���MX�s�SG�����a����t��k�q�t�%�!��8P�)�C�e�0e��AmC6n����Q^e����c7�.��銎�����L!�μ٦>g�h�+�8y�o��V�,,�ԛ,�lG��A]��u`����C޺����Z�Y'p��❣��pG������ʝ2f��Ω��x�N	���dޡ�MG�7�W����!�8=����7I��hP% XW�z�2�����?о�P�ٹ(n}������#�[O��6�O T{�P+��CYmZ�@�5@4�AU�A���fͬ,NN�T}V�߁��pzO��ɶ��ȣ<hw�y�]v�8�w��-/����2e�u�xy�ƕ�8�r�X��b��I�����?��|����ŰH��K�U0>����%n*� �v�!"����/�E1��<��F�t�A���|b	�o���Vd��j�E�ġ���E�:x R�<N���h�/}�E��^g���(+̯�yTX��&����a�W��_�Lܶ��� ��^s4D���̎�0I��8H�:/gˠ2��q���ayiO���H��	s7���'�塸n�H������8���8��p�+��=-�0|�=�*hq"�u|n��L�O�wQ���?�/:�*��M�tT�^]\��F@�7�s�����@�mj��{an����[g��8~M�T.L�gMצm��Ѽo�,�}�s�:�5����u��m��ܚ��NN������Q���pr$p�}�戱 �΍�4Z,��Y����,��(��s�����r�@�T9i�k�;,���{lkN�s���Ҁ��!��*F���7�-����{�罧�*/�Gi�^�1-ϒ��8�ʡ۩/�q����o]+�������,SL�@���/~�e���� �Y[���qଢ଼X;;ԇ��9�ư����U�(��o����w��7.���#e���̭�$��o�}X~���?��ay�l���0�	�tV$!��H���M[=���S�{1!�5j&��I�IQ��i���d��Ca䵳k9�>���R�*gϜ(�s��5A�ի���pŋ�[�_.~�]y����G}^��d���'����r_���D�a�-��L�K�v�i��6��g�[o�Q~�w���^�G�p>���~�ɭ����ᇟ��]�گS�����G��7M���;��C[��g1y1���R���Ӆ�N���z��r�{�ܽ]����j��8�Ϫ�Ө�/ͶGZ5���6�Y�no.���%{Z�֎�N	�/�^n�0~d��f����<��S(ݼ�ά��qT#�����'��d=
iw�4^�4u5p9�����ӹ�������U�\:�O�u�7��fd��2z�å�������K���h��H} �d�z�)�]�!j��!��\�<�\f�|nӪ�=;5����>�3�����������KO�!�\ ��7JY_�,�Kk������)��u���o˓'�U���z��]���F3������7o���O���-����vY�����w���~_n}�My�r� b;ۺ;��9�-���\�W��Ñ}}�����[De
��nn�����N��dR��J&(Q����U�)�� �Q�!|<ʾS���?��{ߵ;o:��h���celt�g�eaq]�$mr��{q���QO����'@ ��m����F��v��[�3��n��t��MvHGyyߴNY�]�$:?7_V�W�G�KR^�� �N���!qnv��F�ڎ6�U*�� ����a��}n�>�U��uV�!��np�T�up���g?(o���j���d�H'�n�4��6���ʈ/�v�:U�v�oA�I?>.�j�O�������,�;�a	8��	7�ӯ������`� k����=����\�>G���>����١�p孌����Eu`֐�3:h�����Cy�H>�Dd��rvȗ��nv�؏�Ǉϼ�]�%�F�i��ӖP��/��}�d���-�I|Е�2��U��4A��+���L� k�Z�[���A�Ed=|6_ֶK��eÐ�����N����d���� S E.v�8{H��I���K�U�uI(2&��W��@{���.ɛ���G7�p���V���������F�[Te���
�����n/���l��iy�m`i�M��k��? �k�&��v�� ?0�<5��vԛW��A�Ar�ס���:��^���2�YL�ѫ�V�V�T�y�����\����X�m�r��y��*�:|YD.mI����C�h:��[����T�u��[�
�|Q˭������?��-4<ka��H�Cf����c35m��?[u��6��.�g�n��
��|\qnol�G�������3j��	Px:4��_걽�/L�Q,��p����g)�;�9�X��p��մ<����m扣b�����iҷ��,<�R	� ��m=�6��Iٔ���W1���2���z-ۂ��y�ԟu}����2|��m�Z�͏&��u�Ml%Ϸ6���сr�ƅ�7���c���ǎ���80����n�������� k��/#Y�4�SI�:����vo�����_����g?y�\�t������Jy�r��{�G�N��_�/>�Cе�!/𦽛N}���j��3\��v���-ꚁ!�nԝ�iYYY�t�r�R�huh��Iw�FT�cmP��]�����,�v˱����7�����?'}�LM�����[+����?��|���B8�k:f��I��OL���G���7��S�ʶ��ރC�ճN�v��Sg�;o�Q���;���sq�鲰�[���n�O��/�?��/����E���ګ,u#����!h�Sj��8��4U��Y�W�tgr� fx��)���m����]q�`���AH�S��ȾN�<K�q ��&�XݰÏ|;��H�:���T��?��;C8�c��e� ���Y]uKo�%D:������rY^^.~�� ��<G���٪𮻽�k��G�]#���s'Ӳ�9apd�N��Ñ�,��Vgǡ��av̮�����ٲ��<�D7q�.�S4k)bK��K��A���1�R~���ى� _�EhRu��~l��[�7��G�k�q�@c�]�?����:R�%�g&˛o^'�z�\�v�u�%YV�����/ˣ�O˝��ʷw����+<+�s+T�%`��`��0�����r�̩[g�������fYZ^%�#�+��/�	H���#�C�ñ��SNA�/r�2�v�~3hdx��o����\����|��t��I�K�evq�,��Ć��͍Ͳ�.��D�[D�0�WN+��\��@F��ۺFF���]/:lRV������p��:QF�G�'��������<T�`<�f�5�~@��[9��c�v`NsC
"_�@z[��Po����@�'�L�700�+_4A�
����,����@i/r��[h��x6��env%�uu"�u�"<�i�C�(����2~d,�?�.�<8����ɥŕ������"���"�^�)+��`�s�$<緧��E/8�1<�j��߃�����ANv������zY[_ˌM�zc�������t9zt"�}vv��n=-^�1Fh8��\L��w{���@p��qض���K�E���lA�̆�޼	��Κ&�v�����ʀ��@w�+�g��f�I��r��F��C��5Ȋ�D�;�}eu�,.,H��NGl�=Ny�~ڠ.���`ቮ�j��4��v�!#=����这���A���/���`�&�t�U05��_~���da�>�/�D�=D�{(C�,G�2|Ke:=���J6 'Oⲁe�{� �� *�T�B��ml-�:���:���:~ְ��?�>,Ox�[Us-H�/�$~u��O�»���U8��.�>��k�N�x枃,���<�5o�E{Z4���W���>�L�+��oX��t�Ѧi�=|���4:�2�
�uSG��{�Z�#�+���<�^�Vxęt3�N���o]mFw>�J[�8k~�Y�=/
E�7x6]��W+�W�B'#����[�A�i�	.�۟�߇KrQ{���,���W�(!�H8�2�UT�6�PD9������ ��cf����N9Ig"q[if�Z���54�"q�
������s�W���I#����-�����(�������Cx<iu�Հ�)�*���*B����D�+O�ߑ�w�|�ʤW3x��8���iCsX���P�4�[�ҎW��S��#y�R��▧>�v�Ĭa@�˹s��O�{����o��N��#����ć��*�����	A�S���-���駭u���e�C�C3�$�sgf�����O�Z9�(�|�)��,�Ͽ�]~����O�-Ϟa�q]3�6���uع`0ֲ���#f3�I��թH�8�ϟ���-�W�G��k����8E@�!38~�˫���Z��8W���H�O~�n9u�xq�;j��j�����?��|��we~^�BGt�6�{�A 4�����׽�u��e�� l��.���25ӏs�[��̔+�.��W/�S��D��#_pz_�_��w���MY�ѴC�ssk�@h�DGZ��Q�m���5T:�5�
B� �~rtGr���*��G�VÀb~~� o1��t�4vz���v6GX���C�2Xu
���n���`�N����.Q���/�G'����p�>˄����)s�s/���jt���� �W�h�#��� ��_�C�"��"غS�\�,�(;_��.�˩Q��7<�_N���h��f�e�]$�ew�5Fena�<y��z	:��:�z���/�s.س�X����K:�uM.���*���C����?�� Kd�g���mG���u4Hنޮ�"�B�S�$Nԕ+�ʻ��,o�y���iu�pi~����^���[���+��?��_B�Mڣ\� 6�w��v�"wSӓ���cy������7�:���Z_]�+��D�Pm�@��+i���1h~��n�����du���!`���-��8ҫ����� k�iv���unv�<z� ��@�:�S��F��S+�k��hT����I�M�����qq~ Fy7Lp7qd2������g�ˋϳK���nh1;;O@��3��,���"�}���P������l���#��ɩr���9R&&G��a����M;�n��KW�׎�����FG��=��%�_,�/�M_}u�<��{�>�&&�����ip�¹r���2c����kD݁R|ɻۛ�Կ�n]�g,�����J� �zj���yy.��ч�J�2M��[������K���1�Y}}N�(�K��<|�0��d�t'O�*�/_�z�ɩ����\��Z��0����,_|}�|��Cp�?�Ӄ\ԥ�f����_������m���Փ*P�r���=G�7���[_Ь�{D���k�U���5�>�s�6:~��	���R���m�Y���OX�6<��Y��ם��'
���� y�9~	�΁[;�֗�v���X�t�Df�\>�\8	�Q��ή������|L���J��3���u$�^ �Ù}�i��\tO@�Cp���u���Z̽=#^Efuu���Og� ˼����@������4��I�H����8��R������+���͖��Wa%�
q�0��uY�u7g0����?�h�@�eg����)2�L�/��z�;�[���	��&�>�m*G�v������|�	l��NL��u�����K^�գʶ�Zv-��X�+���ִ*f�k���z���v�~83�u�G�ba������Y�a8y�<��w5O�/���3��60e�7�铓S| \5�O�XO� ,F�I+�����s�n���GUZ���� ��S�SiX�U��S8Z\���uZJ�<����񩳅�|M`�ƽ4��-������[�2X��i��_pgs|@[4��Uhã����|��O#�MzUu�m�^N�ᾀ^'����W�4���Qy��8ep�U��q����}��;�٣:бUv7WH���-�ݼ���7��;QE�/��o~����D_d͖�u�>�	�=����82���Q�+�Δ��w?+?���r��H����F��p������_�}A���ide��m�����wm�(�;�� ��Gǲu�;c�:��4�!G,t���H��a�Wpf6vp´Y�w	n�g��Ht=��F�4���ղ����RN��)?�ɻ��������X#~k��3�O��u��?*�ܺO��U]\�=u�23U�ѓu޻�Y%8:1V�];[�x�|9s�h9>1����N9��� ��޿��ܾ�,Ӧ%�'8qlp�7h�|l���&��3�	�G���թ_�]=[�〟��:u�8����Z�Z�G�8�$Q�&����R�s�~�s�>u��f��u�6t�"�d�4��4�k�EP������3'���7�����q.w���x=��ݯ?~\?��s��7��[������W��+Ν۷��{�����5��Lk;���m'xk3����A������ezj��:���]����%��㲆�����1�3v˽{��a?q�#��%���d��8YN't��Ә���{u���ի2�=A^�S'��SqV��)
���U�-{��:�c�ֿ��4ȂI	�]���5N�x����6�O~�f�|�l��s���WߕO~�y���˭����%��@i�,ꡎ�!��s
b���;�4Dn�l9�:Ӗ]?��H2��Q�%���&��/&&&���r��)h1��1�i+�i�n:V��������bY�DG�~�a�޻s�|��WyK	F�t. ��Q�E�vy����;솇��g f�:�3��'��c��s��:eR���m'k>GF��F�A2p��;��on����G.�-�x?���I�_�Ug��e�X)W.�+W�]�>'	X'p3���M��?��s?���`Ն:�ie��@��&G\�Z>����/~[��yT��%�@�v��`�Tp<�G s��������*3ǎж�&��"uH�N��G��Jp��#u��Oʭ[w�w����K�G潽udٝ)^����T����q�r�t�\ں��Z<x\�����矗�d����u3��7�E-�⽝Ͳ����'��7s����/~�;t����2��R@`)����F�LyY]��T�M�x�}s�2��ʀ�[}�O�mm��� K�Nr�=�i�N��r�\�P�c�����V���*�E�N���3�R�~�p�p5�e	�0Z^4�&�st� +��uM-2j�e�m���>1=Npu��q�r��H։�2�~���w�1��ey�l䮗5����E��)@Y �[*��m\榣8����� ���O�`c���*y8�:�6�ź"����2�S�$D&�j?N�Q���o�y5Xa[G^����qa�=����ք WF�N6���.t��"��|U�S���u���s�-[��n�i<�H�<���z�=os�rlK��Dy�:kYչ��M���C������Hb�^~w8��G��P�0�FP#Dm�;دo���_\��<�Ļ����;�eO��~�����R@�Ly��-�)~�{�6alyó��"9�5��w����ysXys&M�>g��������W�@=(�
S���ؚ�|�i;6�ц�����<�f����)��4x�tU�񯅳�Wp�1���k����Ӓ+	�ԍ#���	�ű�S=���:xVۘ&�Rj�l�R}}΍��:%L��"�?q�C��sc�pQث�֝��uR�ROK�^�i��>{2��D�^��2�#���&��p$GxF�5��n}Q�c �={����ǡ��ܐN�4X�t�S8�o'嘛L���l������X��'8��<z�J7q+�1���Ѱ��t^�v�������(��v�\$x�at��;w�tzE�	t�\�ഒ�ǎqΤ'|lt�ʻp6��p��P:��(��p��m`�]� ���tt�(���@��'O���w�;8��^��8uR'F�t���f�
��,��n��48{�/^<W�~�r� ��a"[a�ІG����:�N�]�}�Գ_�	��3mǅ��h�L���텶�����L���<y����孷.�g�:L[ul�ho?��d����Sq�*�'	lq���'fm�8t��=�֥���l����� �&0u�������,�u�\�z��95�F����&��^?j����SǲN�����9`={�g'	�&���p���~��w�����.0t'9� n�ca���ˉ�G��_+�߼Z�_�@�G)k4���9G	�ƀ��qp�	�ϝ9��?��M���n�Yu��)-�3��qF^X�Cf(�����M�;2��h�9ѻ��G�Ӊ̽�M���c�WeR�j����`'OgG�Ѐ�lw�Y-���](�Xkk��^�^G	�SN;�p��t��W��J�֔� �q���d��ˁ�n��nǑG?zꇑ_�~5���@ߙit������w�l7trD���<��щ��NL�t6}�/��������岼8GP�5�rD���3����th���Q�1xG�s�� �~bpK��(��0���n~w�$�訠:�v�Sp�>���[����/�l�z����7��w޾^^�20�.�O���f�H-�=)6���pG�ƀ�������/�_oF�;�E+K������<u�����+[ä���gOf���>>s$S�G\�V�U�� ���'eeZ�"8<
��L^<��m��UxuZ�������;����]*gN��C��Vn��np�'��u�^�|���_FFz��͉����ɱ�B����8�?|R�V�����U�2��톦u�D�D:i���)��F���F���;[�����08 ���\Zn�I�LmG޴�8����au�~��6ѓ�"ehiq����5����5+4m�5Uc��w�^��v��7	[����-���������=��6;D��yt=<�����2�nDE����A|���b���ey�|�,��/Q[�@]pV�}R���*�� K��X���A.H��h�T��@���]�܊�ܖ��dR.iZ´�uH�8�£Bu��|[%�:Hk�;[�����M]%���؊Sy��*� ��i��i����!���/�<�&鸷�)�6�U�WFH�ܶ u�*{�[b'�|.F�Wم���̦Kq����Wgu��.���0��;��4]���PF�8��)�SX���I���C~��Wq��0���--�i�S�꺆�����:�)7�\k�k�*�[Z+`\\�O�癏ȧB���8�yana�5�=���O0��ѵ�}�|�
�-��Z��8��`L�&?e�Gm;ď��ʫ>7�6��Օ�:�ee;Sq�#�|Tީ���5�b���_��<����y�K���Y��ͨ���|���xv�=��6Z^�gw���9��B��\>���{^�7�>3��uyZf�mO�;� �$N@�Ӷx�μ>�L �*V%<�NS/��vv��x��|��q������	,�Oˣ'Oʃ�/��GOʋ�semy��n�l/���D�� ��Y��z���N�؍��`��淴�]?}Y��xE���mw�.��LM������-����.JE'؞��~	�A���~�o��N�q� �,�'q$IՀ-�x9�L�'���MqRş<�����1;�3ﺀ1�����\y�܎=w�s�m�f�\����,��^�b9%Qzmo�W���U�38�.4vZ�����:6ݴ�3�%��)�.��?,���]=z�)<�M����t��Q���H���`�@���[o�^*./G&�éu���)q�FǇygY���7T��������;e]��<�SK=���YK .7	Zu��&p"�(����r���֡L���u$��z���Y;3�SM�l^��C��n��q��0G<u���e'����b�x�\�[�t�~�vz���0d���魘Ƒ�g�d�|�6�#�:L�i/2�Ƨp=�|280X�V�u3��E���2�i��n����Lt�HxQ#k�W2/骜�?R������ |�C�����;5� ٩r�0�k%�_X4`rp��.m@^{܆�鹽��N �n��)� ��f�<�-ph�99�ڄ������U'�M���~�����yv���"���u�v��Y��� ;�P�3�x���##�7�YW�g_�a�?��w��u�K�+;r,��*<\���|n?.-�Ⱥ�ć���`g�5��5G�m�A��#�	�ea��j�������K�3k�w_K�ѵ�g�~��ް 4u�=__���u4V�ĽκS�9���p��θ�A2�]f��,�{vn���8ڝ��g����3�:rp��r��f��x&��#@��z8Z���!;��Ĺ*v�J塿�74t����U8*첒u���C����O�k�`w�,� ����Η'�N�>o\*�.]��?5�#ش."
�{�KFk�W�ʓ�����'ea	�h{�);[b��[�Ȩ?�]��&�V9��ں��O���
�`7`r72�?#~dX����'�g�\��M}��ߨk]W��S�~e��G�R��p�1�nhdؙp��lul|n�Qzm�G��=.��A�P4z!�4v�h��z~� �$A�$<p$�i�K����z� �ɫ k���`݀�&�[P�,������ �C#���"l�D�Nwr3�۩�*O��hR!it�t�$�:��}�̂���o:��.	���_7�����:"�d�d���%z�%�,w_d�q*����^-
Ji�%Ad�h� �@Ķcu���IL���WA��_����Q��������.I*Cg�9x�v�J���%x&Sj���
ʄ9�.mR~���Y�"ӫPU�"i*����6��zZ�U�+]Z��N.���2���	���C��)퐦M�l�N�ֆ;��8*4���/ ��#c��+t�,ߐO��ն�^ǿ�՘i\��C��Xt;O\��\�;g��&�=[�e��N`��!\�5Mp������M���<�m (�T5���Q��6m�m������G9�s� _omP��T���7�|g�\�^�2���k;�\���$%��L [K{��̬/�X���ς����U�bͩ*�jv23�OI+>�������/2�.X�{y�:��w&�ȣ�C�`9M����l]��:Y��L:��y��og��ӥA�z�J9v�Ƥ�,/�����>)/g�`�}n�P^G��S����l�C� ~���� �G���;��F]/����9��dN���38�n��ڵr���L������׍l�����Zu�l�Bq��#�. �t�#8��l��jaa6A�ƫ"N��Z��U�W���1�gΜ��mɚ%����Jy1�P�4��IтC�tM�4ȂB���ݢm�S�S��z${h��Ȧ��N��Qr��[mg�u,.��b_}u+A~	.Ap�ʩ��>�a��m����zQ�����5�i��B���wA���{Tn��i0�-�)�����)E	���N�fu���.t�I�>��%�$�8�	�^'h~������'��D|�=���1Wλ�(��(<��W6�� #���Gp~I���G9�њ-/^J�l=����:vb�\�q� ��r�5x�@��m���9���I���^ڮC�:�[�ǥ� �>pq�ZGp`h0����
��Tdb�).�\!}=��z�;dp�+�sz�pp�I�m�N�>���t dt�lw���Μ�ߎ��:�n��M�!O��;w�q�����ab� x8R�(O��Fy�١�[-������(u��������K�˵+�7���>yl�D���9�l�ܼj`��L`�x�!�P�K�t�K]?����tW�!�#+�G�l�#�gN�`]�v� ��FqN{ph	��u�+\�$���&��>��t�L_���n��TX;���M=J�2	���ssea~.0�:q���ֵ��^�x�Z���A"�_d��Y�_�7_�ZZ\n�; �f���r�����Fy9��>}�]77��֋<��]cgG̳gO��rF��������_<w�LM:UV�A|���Q�^e� ŝW��%�WE�a��0v��	6A��i�d笛��H�?s
ڟ�z��O���g� zڑ1t�ɓ'������!;�����#"<�䮬m�g��{���ۜ���C���}��8��N+�^w���𻁖AG�?��y�yܴ�|�6�mK6�'��?h\P���e�{:�G键��#ʑ�U����v|��+E?�xy�N �%�W���7�E���9�"�bث��&#��wD(T��řN<������'f�"��Nt)�P�,��<�]&Ț%Ț�H��Eػ���y2I<N#r�3�
�ڲ:+5"��� ���T$�����Xb~�X�H�-n9��B�#[��%�J�֓@Dv�-#i���;a��n%GyQ��������e�Οe
�x�6��.	3@[̛���M��)��*�8�$�P�׀0��.Μ�չ�9h�
�Uq@ִ_��ob�Kj���lOb5]œ���:�ǫ�X�x�iܩd��}�/�)�D���e۫�_:�>w�%�4X)��Q�5Μ�!(l��6Op@>ӊ�,ٛQidy`l���%�.��,o~����x�~��
� 8���u��vԀ:�>e����8�Q��Ex��<1F/D�76ʮAil���4V6Y'���A�T�T�$]u4��0�~�/��7��Q����Ļ�T�
=U ���se~�)�G���N�3 �V,q��8��H/l��4-��:M�L:�-
�rt��������leQC���欼�s����λ6��h�u�t��;�&uJk��_�TOp�y_�B�W:�(x=��ۼKe�>1�xv(퓼n�kUX��t��|��:��y�\���Qk Y�ڣ�wd=�;jIS���ܧ]45��Է4)u
�#�g&���Х��n� ����?��_[]K�hbfz��>}�\�����r�����uѽN�Fj�,/.��y9�'f�@g��]0O�=]�H	��4V{�Y���M�lLr�ғA'� K�p���0�<u����r����Y����:]oi�n��������@���:C� Ў��aR"�N�k̺@\Pŧ���<nq�'���ly��E��������������5u�������~Wv��Y��."����}q�#t#��E4 y��q���P���h}c/S�i���\~S���a^������u�گ�!��;�d�k�o��f�t�L����s�cҢ����4�`u����Y��u軼��U'e5��$�#��{��^��G����i��v�	���1���-��o<�S�cȥGG7�c�<Z}a��#�XC'i����#$Z�t?y�x1K[6(S甄�~> ]�{�AV=��4��Z�iq� ������T�/"���z�N��\kX'���骓��G	�Fy��I�'��l~4whp��8~��r$g��I�^��'2����t�ȹ�I���qd�v�(�6)��l��� p�����.%�r���x�G���<�?~�$��EN��`9���$���=�5���C�0-��z��Lm�]BOlq+���`y�ojg�zJ[�{��t���S�H���s�����FX�2Ȓ�}�.��d�Lp���|��{ʵ���&�w�g��|Z�M��6��+�!��_��G�a5���0�F���k���Q��ַ�˯��;*�1O��R��37�9�O�k`���o��o^�&g	f&2��@W���dp��"���s���2��C��{�wj�
���E7P��P�C��T7����}������3����#7���;MЩ��﮻t �_[N���R�힮�}�r�ܹξ}P�d�����	�z�)��'u�<cǰe���i�!��7 ��N\Ƿ����^�ۙ6�v}�|ۋ�t�;���C��3��t��gIQ}%�j���ӦS���G��>�H�>$��A<D��{�:#Y<�:K��� ��̧�������4�c�n>4>���#Y��tv�<p$��\Yr��6�8�&��aC��cd�e��U���k�PP L� @�2��WgK't��ε�	�Bxn��0�(�vx�o��@Fbkl+�.��uP)W�%X?�4"Qd{�YG	���3C�k� ���Õy����B���V{�`dwF�h��!H���P%yZ��o�U�TG�����[�?�O\��uF�!6ޛ$�O2���l�����)LՎb�N�)���:��xKPJ����i8.�_^\�B �,Gj�'��(f����'��4��P &�yt��ϴN��S&0�~�c����7(1�k:�uu�=�W�`P�= -�.�1��cp&���߄�t��N�S<�åbI ��f
xJ/��Q9yR�t�����������N��W�� �v
�48�)��_�u�g�y����:'ټ�.�h�t���O:
���n�x%"�
�0f4�r"s�e�i��Yws�=Ҏ(�	�.��9sZ���/4�8r4<j=Qz�%���������,�>�R�`�ě;���q��2�Gʈ��r�W�!��o5�4�x�������Nv���|מ�G~O�U�O����D����rd'�,ո�cߩS'���W�E��1�Ņ�l�|��{�>A�;�՝��z2z�&h����^�q��)w�:�4�����Y�܉
�����lT�S�n^'qڜx����.��+����o�8�iC���� ������ݻq�t~�eJ�p=�N�����lP��s�����75p�c�s��|H�`Ze�@���'g�����8��u�tie;[$?����.Q��ұ=�!�X�W��@k���ґו���]u���n{iɄL�&;�t�YXX �}D{�o��[�/����Χ:��D^�)�L�t��0��8Ig�#P:AO)�~�}�^>��&:�8����ϭx-�(>�t#7���::�=�&��S�ޮ!x��[�ն:��H�k+^'��N�|t�٫�0�q�FY�!ӑ}�Sf��ӿ���рG���8�Ϟ=ˆ:on��-�Ǚra��#;{n5�[�݁�>�	����f"U��Zy�Y��U������:������L�qt��X���:=狠���?h 7@ȿx7m�(�pr�d����oe�:�6*󀦭��~K6d���g:-���=�ò����g�l{�ԓ��yl{}�]7\����z��f�6���!�v��#G���sA5�:s�TΓ�c33Y;u���Lu=C�>��Q��󜁯�dv	�P?g�� �䱙r���L���_���%���e�`�1�w��.���/��ݝ�ҷ�`��n�k��]��6�s/_�%�#Iv�i�]��
L��'p<K�5=5#�isD���^�~��������mt����u��{�">���8�urr<v��?������6z	���V���gݸq����k���3��lr��;w�ʳ��囯o��8=yGߎI�v������6wH�|��7壏~_>�s�n���?�	<���t�)�|�b�^�VΟs[�Q�^�]��2��7@�ޤN;�?~^���#\�����	^�@U��\B�7W�8]Y_% Z$�t����ų�O����1xБIy2Kp"�a
�����1v6�_���)������������v���h�3�� 9|�U^�Y�`�琯��w�_�w�}<������~�z����kY���{����*��v�Йl�p�/�A����X]�M��R�A��������c�eX�|�X��>�#�=����+j]NG_[�����R:#��� �d�ut���Q�##��n���T����˜n7��q���0�ȟ�r.��a[�;(�~�۞I��L��{���ͩ���8iu+Z SG_pTA�H	��^B:���罍��~ ��!�d	��j��q3 ������ ���g:J ��v��^G.t��Q>�0`�B�`���P�(�^�o>�)R`�N�܅Q?��5�tǖ��e�b�A�ԅ�r��>��on�������m �D6RnN�	/�c���F{�8�2.&uT �]_)+K(e�_�д���]I����O�ŹO���-�5���:Y#}���;wً���=)�~��&_C��Й�,�3�s������/�v݆�1�: |��i�C�&�^oO?��<.huB��!x
�y��RyD8�W廑Q�=��^�00P��될D�����Ac�^ozX�ݢ���9�N	Q\�6Q�,��hx���w��r��Bow�:J.~�-*W;���AՔ��iO�������)mo�Ҧ:�����ֆS(�zH��s��
���������`�UU�ɱ��J>G1�Mċ�W������)�!t�Np�έc��<�+bpU@8<���� ��̣�i�\Y�>�O8� ;��݉ąۘ��C�l�`������3|ե*��l�*xX��|8Mb�s���e�S���;�7��
8X.;\i�S����Lۀ&�p�����5箻�K~R����xbB�e���ڔt�۶q��&�Fn�)�y��Iz��I#�o� �����ܙKC3ȑ�<7�b�ܹ��<~�>߀&���ckNw���Q^ԁ�)�^_������p913VΜ�(�O-��ҭ}ݚ��Ç���enn6S�.a�_�f����r��29s��YV04G�ܽ��|������z��c��G82O)k�`��iy���Q�!C0ƶ�������\f_�`��`V���S�#z7����S�g�?S���,���lo��O�ʓ'8�؝5�#{5����YGv�]�Wh�����H��<}��,��o��%����';��]�~��q��w_�O��Un�}�ӷ��x�P$4��~񟐥�v8��Z(�>рk���t��^C��>��<x�s�c{�ν��ዲ8�Y�_��G�^�/>��|��oʭ���|Y_A��uoO�4�@ꡱ{�'��pj'A���,�m��'�ʵʛ�\/o�}���1�A���=���S柭��?�[~�����/��/�������[���]����q�^�'O���=�{�R}| W+h����	_ �����;o��s�\9�L�a/�q��s�f���]����rK���5��ww�g�}^>������$8^�e� ��:�N9��;-��ĩ�NM�׽і�!�?t)������g�_�1�����7jI��d�m�<�.P��(B^��!��ʓ�ɡ#exl�-ݽ�Jo�Q 'GP��Ogbx|��.G����T;ҋ���#�=�v�� ����N>��Ͳ���C����vn?h��E�L��cC�`݄^�~>#X�s���E�uy�G��,/������"��<N�,�;�d;	ֱs܏/G�ж��ϒώ�^�;�F�$Y1����+eq��k�aV���=�]~q�v�u�^�#����͉�Y���W;�ķ��v�w���mxy6<z���r�Ƶr��>� 'd���w���~�I��/���ei��C���X�>y�.~N���3G@�"��_}G ��=���~��(/_�797Jg��v�\�x�����ҥ�e��A�������NW�D~ܽqay�<��,)�k���'��}��4��i�� �l��x�ƮWG�9���U'!��8]�Sl� ������ezz:#Cj8Lo���+G!�N�]X+/���ťM��Ot�[��]��yp��|�)r��=���/|���T�e�`���i�����y�����Vjx*d��?I̑u}~g_�����U�� ��?BfT��)ԭo���n�����>����=q!��r$>�����Î�t�R�=Ϊ������ f]�"v럈����������ѱ1G��gG'	���R�,���bv�z�ܑ�����[Kʴp�����KF@p���Ec��iV���pO�*\� I՚���J�4��d��;8Ju�|$0�pI ���̣�����s͍H˨��ރ�3G���z�>���8�"eMT0k��N4S(��#c�W�����c-�#�Q�:�:�ٶ�X:�~� ���I/��<�׉����{�v^���k�T�:̊����"3;r!�l����3.�T�}0�۟:�)���3L-|�C{��]�j`�_W#����:��)�rYYù6�i�`�9�k`E�M�GA�W0`�ǅ�fP��V�n�-~ċp٫k����m�x���V�aϾ��a�Gb\X�e�ŰSp�+���ǐH#G����+�>����yΎ^9�P��5^���1��ڝ8��((�/o�̠�K���*Ѧ�
D>�'��y$ȲL�GFh�����
�<��wq�!k+�I�ԡb�yz�U�b�'|.<6k+n�!?Z�=vʰ�-�ΈA?�3�����1on�!���L�*�g�k�'��yv���U�.�� Hybu �����S9��lc�k�)���:�!`>�v�+���tI�Co�"��ya���jj�	�t`�He�����m���!^q�h�c'��yJ]�YV���'�	&���^�U��ػf&��	��t�(S�_׌� ������r���rlfڠ;��V�O�>�ax����#�w]عs��̱qʱ���t�b�<+_�m�/����Ɓy���r�x�b�@l�z1��p�!���qpD{�����H9"�����
�ȣ����AB�3��h��:�gG�Aޣ��a�@��z�#�0x�fʾzB��vZ���R�Q7��3dn'r�%����&�Ǧ2j60<���?n���'��{D.��v�u��r�x\� ;�r͈�t�o�K��+j��ndcey�=�:��y�Mڱ��^V�p�:�#��u����~F���<���Z���O��2:2
_��Cv2�knv6:�5 W�^(ׯ_��;�n3��E��p g��ۯ�O�%�җ�֭;����'8h�˷8vn����'����X�B�C#Ù�!]D���r�G��'O3ri/�S#�x��l��HN�q]Z\���%�}���q�m�ìG|D����_��ch����J�Led_F��@3���u��i�vP�{��f{x�w͡Jࢎ��W��z��VOܣ��U���֎���Mc ��N񹝸鍇_�h����)��%:�;ȊvJ>v��>���~��8vHD�غ�����}�;-J��eʁ��]o��ϣ�N���9-wz- O��]������evn<��������l���4G��<l��9���ZLN�`�����Kxx�,#�Yg�<���v�����9R977\w��t8�����r���r�;A��0�t�ɟ�M ,S�ի��h��#)n����́�Rsz����ezf��|<��G�CTrJ����	�o����sx�~oyi5�iNOV�=F�ݿ��<x��`�9�L|i��-g�8��ݽ�U��\�Ȁ#I�ex�>p[��u;�6�]�g/^�{�[�=(_~}�|��7�Swb��>�0kG�� ��v �}�ӻ;	PW���-�'��B��rd[33��e�6�rj ��?��Bȏ���<u�ӧ/��~���' ����苻w�^k� ��~{Q^mgu�!�Y�Ax�w�v�[�I�gD�3�=�-����
׸�'�3�����U��wf�Y��^噲��N�f]��l�7&�jg�#i[͈�>�2[er7��y.�-y\/m��Hg��+��b�� ���v�;��L�wDkr��wuw�Y/�d�f�AV��P+�4TKg�-�H?���V�u� �+��a�#��"�"�2��bC��$*f2�ߤ�CqLo0f��H�ßm��N�'��* �a�e=�
ru�ܐ֏Of7�����:��l�p�J���5����O��84SS:>
$�?y6^,��1��t���7N�;�34��*(�Td�@������� B&P�Yp�ju�%����5�0XPa:t���i����-b	;�~��>35]���2T��3�t���WZ�=�]{���P]t�4:�;M�)N)P!�����}JŻ�O�i��}�Y�C���]$m�a[2��ѯ�s�yub{{�8�k.Y�xqu.{n|�;�_O�rt�̧��y&�8u$�)����G�s��N�w���J�/o5B�h��3�gą����#��x����@�z��?���h��4����Q��q��Q��ɑE�H�%���Z�|Y�8B�"i�K3{�L�;������=9�D��|7GZ�v{����J�jl3%?������;yh2�Tg��Q����`^��6..�����7���AJ���I8B�g&����Qd �g�0����Ѩ��!�$;?��:�ʏ���N��}�Ϊ�6�4xrJ���.^����3�9���[[{/���N�����>|���"I�_9�9�	���83��9RF���҃��Ř�-�?�د��)���g����Nu�F�N��[�d���o\�q�?�t���C�GE����s8��c�q�g�M��5�}��n����8�_���p����\���p>~���Ӯ�pݖ83�r*l:��S:�_� ��g݌��65r�ȟ2��w�E7�8M�u�ı�K����m��;���>�^�r�Үn�qA|��&p��#��<�����}��]$�܄�1v�ױ�3����G���i�_��O?��{��U��QE��|Iĩ��?ڣ�ӐWXc�	w�Z[_ɹ�f��ѯ���^�q�\�`�ܖ�k�t� o^k��#���iQ��2��1Ο�5�?v|�\�x� �|9yl$x�"0�� ����~U���v�ҧ~.`y�`܀y�̻�`)��"�j�T\��r-�]�娟<���|�4?m�i�]�p50R�`����@�6��[���%�|�ӽ��)ڦ��∀�������jK�U�cc�|��;�qg�QG��-�R�}=����!��W���=Y���Uxί�K)��M��4>�>B��Y��*Ӫ�j��d������)��ٕ� gqq[Eb�)e�ઓ��w�Y�Ux�޵L@#�2+��٩�-��Y��]�Y�T�y\��g
O8��)�l��w]�Q`L��i�C'S��F����<ڽ�	rn#/�����7�u���wuDġ��+.�1K !���a�����*�`�R����}��V��	�r@~��`�@����_̺�	�\Αu٤����t�N��U[��	�����V3�usGC��/w}T�lm�anp�h]�ϒY-�. G�F~��OV�G� ��H�C�SSv~�v�N�M�j=����/�}���l�*��!E[-�{N~҃J�06g�]G�����r��kʸ�2�L���2�t���	��=t�����/���ʝ��c��}C �?>����w�
I l��j��S����
�o۩�ª��l�J�������K�cZ}se��ٱ�����i؎jE&u@9�_�T�COy�gԅ��>�Lԑ��z8s�����((�Yc�W�E9^�� ��|�2^0�V�TO�+pҞ��Q�����55���s��CA֓03�tM�_�_7��1b����E\�����8BR7�p��(<�� ��& �;=;4���"L�`��Cen���P�=��D��%��S�!����2w%��|D\&��&���8e�L�g��SG"j6��� mA�E�N��޸�ſ~ߡ��T�{r���v�ݑqN{���}���r�̙��GF���p9R��#=�#���~;�����X��Ӏ�m>]D�r]��y�:��z��j̝8::HY#8bG˕K��{����A����Uc��O��3Ǧ����S崻���0�|m�,�l�=:�8p�밻���:\�q��I��
�@:
%�2լߞ4iS��vz�8y�Ζ�5~_���{�̑a�6:A	f��w�50�)��(��1���Y�`���p��8O�v}	�>h[t�g���z\�x���,�z^Vr8������Sm�j���3�����i���`�]'N^�Gb����?�s��l:��љ��onu;�s�u��]|���`6�18;�A�GJ�����5<B �|����w�)�G��Y�NV��<r� ���ܹ���������,2�_7���p�s����O�����Y�p���tP����a�� ����҉�a�3��hL\$.�=����,\����Aw�x�����"p�h����Dh��q��o�(#T��`v��G��8��ݱ��]載��	�;}�`t�OO�FS�K@��եm�[�ѣeei)���F��b����Yv��|׍'9��#���G=�q�C���6�(��ɵ?NC��ޓ�4�ʫ|�b�a~��i���oʧ�|��ƞ�M�=�/f�Ή��N���NI�E0{�@��{w64�p���fl�`��鬪WU�n,$/��ԃG�ٳ����S)q6�C�����t�����8mM�O#�=�,�I'8	n�R�ȋ[u���Ny��wZ�<O@W�Q��5�+�����Ͼ*_|�5��
vK�i >D=M�7jo��?�Şف�Y�6�P�S(߷r�m��w�426����ŏ������4��	{�ʙ�/��h�kM�Kg�����N��؝��w��q��gO��ɑL�q�������W�K��M�B��-�#8�Ξ��J!Om\?0��)�����?E��Do��P^�&pz
��|� Gk/]tM��m�>/d��AuM_]��������]��35=U�a;Na�N��i��?�B�� ��u�R�w;�W�[ƾ��F���⪽�w}�3�%Mns/�$����T���j1e��=�o�tt̝��(����8�R�ܩ�n�ﮙ��:����%Pvڥ�/�ծ3%��5p��Qmg#��K6HX]!@A&�_l�q�Z?�_�Ee�e���B��:It�#��vz�w��'�r�q���k���B>���T��(Ҏt~{�;��o���8��5ОD��ݾA%.SF��1n��f<��g�e�op���V���}��&N�ՏsY��\�9�n�w;�l���0�?�:˩�|_N��2�sY��t�1��.�!�7�w:����H��kv�$`2����YU���::��nv.q��S[O����äz���[�u9뷾��;�+O�:�1���b��|�:Ft�<�D ��J�j ;��qD���Ԧ�������o��W��:�)l��MP�8Ŏ�~�������)Knv$ݾ�(ڷ�SGќ"}�t�f4�BwNtO�;�ʣ����k@�)Z�G�iD��`ɷҢ��:���0��(������ď�����Q5X�����[��ik�@~I���}��d�M���K H�m h6}w�,۔%?��!�kp�Ω1C��0G��w�� >�I�G�� �c���J���{���|Q>��V��d�̮c0�Q�Ώ�9�gD���ysmƙ-[kek��`��=�z1`=B�U`m�D
�h�P�I	�i3*��6B噴 $۵sc��o�!ړm��[�Q�����r�����W��0��xߛ�� ߩYN�q��;o�V��/��������L�x��qy�bz��t��`(8:����c#]��o���0���YCbtBZ���}���}֟�[ө��F�!�!͡�V��K�S<�D5�=M���"�Ĝ9y!�#_+++�������0d�e�hA�J��S�#�(�	�(ewf������G�ǩ��@��n1��a�Q���:
*.?��c�fG�[�X)��b^�O�vaW�@uҮ�G����Q(q^�ʡt�p�����kО^-�Q��ٶ�ťe�%
o�O��K�N6� ��s��\�V��ɓ�\�y�iiw��#���L���A�/�b�f3gܶt6�pǍ+0�n�1���=���;�r��� ��4��5�^��n>8T�\j�����������0�V� x�/�bR�xs$�)~��Ѓ d�h������3O<�&`h˞�l����k���IG��N�葉�:�Ϟ>�����S����r!?A;�Ng�My\`�=M�aU�z�g�'��GY9�V�Q�"U��{��1��|-��j�+S�-S"�w=��\���7�p&b���h�Z;G��E�?����������������Η�����,���/�ln���"3���޲���q�.]}8`]�h��נGg9�x��;7ʟ�ٻ��w_ǉ�h;��A���_�~�!��#�W�^*?��;��Y.^:��bD�"��_}T>��S���u�4�p�db���s�no��i��'���o�,?�ɻ�ʕ
�^��e�կ?.���,_{�E�앧L[�"=�� ��t9�Ly��1��뛯�,���)������>����_t�4�:��n�����m�~�v�~-&��`�6�1��K�ϗ�޸��N�;����\��߿_~���ƪ����vH�����Gm�L��7����t*�=����&!)��>X5ʶ3i���L0����W��|+�:�v|<o�6����ezf��:����Y;<V�������_�����GE�]g���Ӝo�u9:dum�<�Y���/��򻏾��Gn�)[&�'��ؑ���<��E�����r�ƕ|������铘��� w���w�d�ߋ�/�{g�����ߖ�߸��b��@�	*��S��u�����@�3,E@�	8G	С�v7�XW7@cğ9{�0Mzl=஀��~�q����3��a#�R�Οk��	�Ɏl5�0l��v�2<x�ܽ:=ۇ2���	Q~��y��ԯ�GvͭSϝ�b���\�v������G���Q\���ۦi���ʱ�S��h�:z���b��	�'_"�����(�ّ��I|�!l�L�p�T9wz�̸.�s7:�uQNכ3����c��`k [�>tFA:%]�=�]r���Z\'`;�z	�7�w�n�_��W���?���r���r���r���2s���8zw�|�|�ɧ�朻ځ�Q����(��?�ya[�7�6�]W�ZƇ���~���^��6=},�ʽ{���������y�F���S3��'*��ך�<���溣k��'�զr�C���J���(֣L]~��%��}�+<��p�Q�(
����iCϜ:Z��߽[��^�t<vB�r����ǟ�����n�{W� ���I�[dg������c�L������o������r� N����vy��/����m��o?�~���י�ؚS�_�Y��{o�s����|~i=3��s?�̾��6�3K�]�q�j�.i�2��ʔ4�A�|�l��G��ř>��bG��R0�#�1���Q:��ZV9�C�b��[9�J_U����m�Q[�jL��ʢ�n�f���	��K�0���i�f0� �?��p�S�����V����Ҁt^�����cr��U+�*�O�`�3>�_N�)�.�.�q�\�f_;���|%Ț��>��ny�ן��~�my� k`{p�1Y�;B5�P�=�4�������j�� C.���`��he�;�:�A���� Dk!�!��f���,����"���(�M��L��m]��}����<���Hl,�m�-� ����C�^9A���[o������8\����kD�*7GdTNuF�2�`�0��;Ѹ�ZWy>�<C�N+p}���JH�ϠL����O���e���U8��[�Ѻy�}tn|p�t�s�c�Թ�S��OO��u��JGOG&5f3����YNm�A=	�ܙ�ު�%迒��&��]x(�ێ�JЩAY�~�s'��J� F�*(���N�rJ������y�	�Bw�Y�i�$G�K5 ����("ʑ�Pܒڹ�~�f5S���0��y� ƞq���	wRtj�J� ��UԮ'�bif`�?iq�47����4�쎆cC���F�Ky���%�18���U��0u��'W�+(/��	�"R���D
��08�1��/��^�2R��?�/*!�0���u�	Fm�m�m�eue/SA�=����������N�@ցC|&H&��<��t���sq���f������$�w�tvנ��-3SU�@*}�k�%��� �;�VEN��G|�l�(�^Tvų��T��L������#2N�tM����A�/������8��ԣå>u�4��ߔ��?-7^;Y��KO��;�Y�������k��ڪ���������9�βݱ�"MV�?A���ြS~�1�x�lt���B�{����w�����	�~F@v�+о���G8����	0^<��l�0�8c�ow�S��n�#���v�긟���r��e��qx��-�H|V��~Y>��+��Y����FZ(�N)s�����~#��v����w�� '����?/���g��;h���Ȼ!�~�Sj�PH� ggu�����S�3�N8\+o����Uh0�iN��=,���~��mt��@=��m���=��t٣������㨣W��u � ���$�F�{鈍zҩ؎�_��-���;�9:agd�@W��]���ä�kB>�=�����M����«Y�g?*�?�oDO�� ��O�,����_>��g�`	���>vڎ�Mt�;�eJ,���+��A��{oC��ֹ҇��0� m��	~���[w��A�dy����>;[2B}����]�Ӻ��~FŲ�Փ��k�M�d� 'H�!���3�0I��n��Ï�?�����o�á6��!h��o�,�c-t�A��1�� ��E����l	� ��S�9p��=P�b��:`��`Š�Q��8�NO��X+��/���R�y��SX��.�9z��d96=].�p���W��\X._~�u��7�.w���+�/GTϜ<��4'�;b��s�s��#���'i�No�{LS��Q���<�3��n8���~���)���W�$x���v���Ε��|�\�r9�B�C���Ͼ ���ܾ{7�5G�\�.�w����z��#��mxpsm�\Ɔz�_��Oʿ�?)o�u^;�~�*��/�_}�A֯�̾X��u-���(�N�;����˟��W/b��^��e�_��Ns��T��O C]���G������
�?,���ߔ~�qqM��p��>�4�&HV�A�?��7���������5��}�����D�/��myH𶵃/�맄��3�� 7Q�Z}k��ѣ�GM����Y���'ꇥ�W�˯?����?~�>�M�M�e���+W���~��wʍ붛�}�4�ٹ�lG��ǟ�_�i�����}�凅�G�-�{��l;.2�O���W�������'�l�~����ܫ6�S�m����'��J}ByN)�Y�і_� }y��4��*�՟�ttҒ%�����z�k��9�#\��w�g+<�6��tn�d�����M5f�9�A�0�a;62����r����7���玕�'��1g(�w�w��K�;_�=z^�0e�`>F"�����%���ػ���ei��3�	W�X.9y%���ۛ�Ek ��l�"��W��kEW��kK�68�6=BU�:jU{�`�����:�����\�+��P�l�@�5E��$����x9�T��m��Ӊ\{�:��#~��lә��.#~ΩZ�N�2@%�ʖՃ]���Ȓ_��8����2��P��S�4fGG�ĄS�,[V�HG,�`���5=5��X������D�u=�y�}I ���T>�e�-��9Lp���ͲW��\�>���ǩg�p����\�n;ăC�Nw�cxNtz��N�A�S�\k��&�q9�ѮI�?���V��c��� NApZ�1�=��|�u_N9����)W�L�۫l�Vw��QqZ�e;�pf��V�x��2�����g��S�����LmsZ�$�5���%��W�a�uw�����Ŭ������)�pJ$4�ݼw�H;S@�ad��#�3h��&�!r*�����̯3��'w[;BZq�z�>�<�v�S��#��
�m���<ly�Jcc�l �`�x��͝,���cGʱ���1��Ld]P֟�{�t��j~G t6	�{�qhw�2�N�<�l����Ɯ�%쁴����N/��v��MO;�zÓ���ظ��.����S`GŃ��#K޷W�<�vcCerb$�Y�Rwr�G�e.�;�����N���������A���mn`L7H����d���#:M���I���1�^Z#oW�`ݼq� �fFN#�C�{t�)����e��K�]�KyO����S�!G��~U;ug��~�Ι��(u3�E���p�\ݻ�F3��ѡ��f�����?J���ؿ�܅���1�Y��V(~�����Р�t�����ŕ���Kk8�N���U��|S"z@�Q%��9���{h���Q=z��i�X�\��>��W�x����h�<qra!�ĳ�0E��NP:�G{��k;|�ͅG7ח���:r�_.��w�z'����kר�l9s�:p:�S�u���#vR�s�[�]��R�dZ,�X������Y��������3�؛i��qR7�?���۲~����e�ږ~�F�2Wl�������U�j� �D�t�LF�zx� �`F�����{8���� 6�\�(n��Ў}�O�i��P�Mtg��O �ȑ�<Ќ�����q��p�q�)C��)��ё]eqq1m��9훇g�}�FT;�����l�;?DLN�U;��}��{���#߅��U�۸Wn����dw?n�d/,�e����l�,�Ļ8�Nv�)'�Kn���3�I;m�Y��Bv ��f��2�n� @{�U��;3�m@/��]�>;�ҹI~�,�������G�B�#�:Ե��L��k��cNv�tE)}i���Jq�GO��s}Δu�Lݚ�ϼ�#���TA�c- ǎ� �x=	�����lGo���p;�ک�N'wʷ��W�]�L�[�'�C�=x���>��)�o�\;()���|�G���<�ѩOc�!�Z�3��C��Y�Kz:����f;Cő0u�3j��'���\+��`;��[ڌ3����1�@X�N��;�a�n6�YX\��Ki�����d�wD���Э�n\-7�],'���<�/�s
�˫kn� �������l��n�-�~N��6�e~����Xz���O~�^�fY�k���Z�h���NM (�/�ā�@Vf�qo`��qt���L�3`��*�����LУ�s�)�?���<�&��-Kޖ�kPXˑ�Ų;0v��'p����Ά�֐!J�a����XR-/��B����ڱ�!�*�qF�RW�⿌�ק���������v����w���� �>
���ٲ���;�1"�H�z���\����F�4L�gD% "dg=��8kУ�����%V��zJ�R��m��1VQ�y�3���5�=���(��H� ���%��%�� n��<(|{K4~�5k50W.��W��\R�L!lug={�5:����t���u㊆X��i�:������s����{K�PY(@:����;��a��aP)��:6��m�(���^�^� ~���+������\/���:���D:�8��t����P�Ʀ:�:��g g�ie��(V�T4Re0����SOG]�[ �![�	�`o�=v���C�+�ψ�T�o�t�&4���f��t�B�@�m?iŷg�x�X믰�;�E�Y����\󥃮��:��-C�z��)픋�iÃD~��H8`8���;�C���>�s�D졜�]h��i�:��JZ���;�Սl��m0��1u���S�@�hd�
�oҁ��[32i������r�)�����·�N��n�w*�VfO�D-�d,b�t
{z����h.{�C��buP��1z������no���V��~��:�!?#ZR��nyт�cz�#�խ����!`@���08T�\��t�wz���������WN�8���Y.^:�3".�G��\���YN��Jp`À�]$�By{w5A���y��k��?~����լ�'ش�8ξ\*w��W����Y�ĺ!��K�5��A��/Aa����u8���V~O��fwt47b�T.4T��7�8�q��%>N����LJ�}��Z�L���k��х�&�:�ng�k7�d�#��:�!�������mZ,[k[�A��N`�S��s�ܸ��o���B�|�-�/�/�q�.���G�# �]`�g�����\�SJ�k'L�(���v��ʏM���o�GƯ^:[~�����^y��7�yh#��R��*�Y��2�P�^ʓO2ҫ���9
I�~�T�����<}�N`O2�Վ(��u��5�\��s%�Y��B�N=|���+S[�\�t��CZm�r���ZK���g�u��F`���1�Ti��:����t8ݼy���+�Iw
�62z[]���~�V������vp�ϟ������@2-�Fw��3��!�WWw���2����<�۰FN
�Y}����:Q�
#��������Iۜꄃ��L]oh�͓�\�`Ge*յ~
%�oA�+W�g�ʖ0K��y�I������t9s� �)�ΤqV��~��EY^Z�=��>��q����[t68T�����keYE���h�N�m���i�ڼ���v�=����/a][�J�x����4p�g�����KE3�1��wt��%t���F��-��޾#��A ʕG	�u��r&����̻z��u�\�|���HxP��3ɵ�~����` ��(vHN��G��O{�~�pWVu�r}H��#�a������zE�����~v,n�Ѿ9ڶ
lN-�g������s�UD��c����cдݍ6\��k���P��3�.^(o�������΀X����Vv*t��Y�A��hu�ٳ'��n��rD�L?�.�N���n)��7���.�b8��7ؔ��73o��"(#=����6��T/x8�Ù9��<�SG�x� )gu֍vV����+H/��H�r��z?q@j�V�fG����ȗ����� Q_�z��Y�-O_ĺZŠ/׎�Y�O��օ.�>֥�N�@
�[۬��S,��W>��p��A֩��)S�]��[�������\��ȍ/�H��Ux�8mp�,��A?��p��,�ёq��A�����9��Pd�+���)���<̓�l�{�1O3��W�i�`�pɜq�e�U��_So	av���q��S&s���FݠO#�S{�n^;_�x�Zz�p@gX�Рj���(�V�,�ke�@��Qw��w?B��e-~h"W��ھ�C�n� @���ٳ�(�4�e��1����:���[�u:-�!}?4��tl����e��i�h��7�Y^�J/�����S&��tH��5���qꔛj`vP���ҲGL��#�pJ^vs���Q#Mz0
N��4�� �;����<0t��	F�H�G��tM�o���������u�];����r�챱��6P��Kk��1�@��.�##Y(c{�tN��r�t6��`@�"��&����A4�C�8s�<Z�R�Au�^�IO�[�o��A�UʐGi����I�gڥ~�*�*����Pi�&�5�w�H�4�ԣl{��@f[�/၅�A�j�2���H�ݰ�{{�!S��k�����*�|��7y��կ����a�\G�]�3 M�L�o�����N�}wjۅ��O!�r���B{%Z�!�E^P��z�.b�SC��{q�\p���L�A>����,����N��L��M��"y��lh���c8 	�N�'�W���Ӟ#�s4��������u�ܤM
�2��Լ���)�o�sr;>��	}����Z�����o����;w����k	�t �SD��0�2�����.(���M��F��ER"��_8��0_��r��\�D��*�~���kQ��� �e�`=�ǎM���/��	B�CbE��k��
?����ӗek}�NkQ��?�6`��5�6��N:�ʋ�\>&;�dNN`_(C���A&׳�Ɲ;��=A�����	���x�P�tܻ^�[zΝ.?~��g?�Q��;;Y�E�k���zKƬZ�ʒ�i��'�� ����]��YwF�^ީ.��S�����}����;8�����iM�EZ?֫Nw����π����i�� ��hgv����s���s?D��k�ݹw�NY\ZȬ���q�j����)7U?�l��Mݫ�0�[`W��No:��2�猼�';�ɍ2ו��l����|֚Ŗ��FG�?ur��o�O�*���ÿ=*�mF!�����~ub�xV�����BG׀��~7qe��A����6�����$<h���]�|�,�ۏ�:�ct����q[c��H^y�!�*Ǧ��ف#Yv��s�Kr���V���ŋ�˔������"�I�ʑ6A�U����:�h�p�C��[�~��H���ꯋ%�BP3AY��c�:��#��"�+����� _V�/��p��8w��;'O��)o�~�ܼ~��>=��O�SN�_%�>�~���)�ʙκeS�����V�0����1x��Eϑ�S��V�+\��dԒ���<�lf��c��H>�7�eЏ����K�{,:��ю>:��i�+.�F��s��-r�Vb笇s��؉�r�����[���i�u�PtX*���A�uvO��={��m}P7B:2N�����ʎ��3��wf�[X��؁�˩ش�z|	�6PfH���5 ���>:���{�_	8@�:ϩ���Y�[�ѳ���V�í~^����Y�;�'�)���	|VLl�|Z;�� ����꠆���ڷWq��1�k��~��%�#�nt�>�?;eٲ�;�+�'�^�Vod�D[�U�T��:�u
{791Z&G�K�A���;]p� ��.Xw�r3���~��{x�H��*��AU��Y���� k#B�_	J92����)aD�2�錘�B[g�V��42C`�SC_ג4=��)��W�aMl=�-3���ϑ%�!]��{�tD�����PN�qj�M��r�]�=�~$X��Q��s�#0mq1e���1�����g!.�����>��]�g��pq����I�kV��RGAT����1�=�Ϟ��9�㎫��x�k�苣%�T� u�q����]���~k�62�fϋS\�ˈ�����\h:�)D.5ؔ�*@���:�o[%�=}:f�Rf��Ƽ�;������-Rw����\�D�&�Ǒ�l��Sq%��!r[=�u�n�Zu����5b� (5����}I��Ϟ=�~_�6l�k����Q��G���at8��Nq���=��A�SF��S�:	&^�#�a �&爻HZea��i{�Mz:"��v+Y��9�y�ګ�9�����}�2��6m����-x�28ݍN��F�T٣�#_�O�C�ʗ�u��Cڶ�L� ��k����P���ke���+����]�G蕧O	p��קO^�j������y�� � B���ى~���q���l9���hd�8��r��:9�ޤ\�VΡ=��r��'�5���*S���i�){�^�8�%Nt����z0��{_ʶ�s/_f:��@��.'��.S�N�ё�E��$���������8(�0�\HO�涛g���Ǒ9��7�pa�F4� �c�^�[B�>-�o���z���k�w�(�0�N=5(�7RD�P�3��4�9�2��K�u�P�Di\u�Պ�B��)�,NA�{,�
�(R��?�,���Ӌt��i'�1X�����T��#��xQ��^�r��F����'ș�t]��'�-N�=���S��*��:�ڦ�,�8��܉����3q>��Q:�	zh�L��m��!��2ܐ��,�f�U��H��:Dѷ޼Y���~�멓Gi�q�t\̫]����Q,�&��x�����|��k�@�;Nm4/M����>z�'q��NB۷�ػ˩:'N2稲:�ɣ�ٖY��*�4�ыt5 R��{!��^q�݅󧲉�����S@���/��2A��8Ϝ=]Β�i���|��
m�Y���8�t�ێg%��@&ww��vF5��8��FK�Wu����=	�^���|�2������Y'��� �>+���&��	�y��ϤV}��̳����ͳ��&�n�LA׹��O���4�m��,��zX=�]K�h���B$�A�O�g�W�ߝL7t3����:��V6��_d����]*����LyW�B�-xkqi)��>�t�ǎ��ב�v0;�k���{�\<�^�C�)�����|���n����˗��K�k��n���/�ӱ�	D���BQn�>�t��V?N��rF.�c{��߸Y.]:��)�-i�����)ܱ�|܂�o2z���u'�Օ���.�:������΋��k�jǠ"�F�7����C;?�{)���t�De�2n��J�K�a���k7���޺I�H��Zg����'��ofܸ���F!���@�r?�`���kW��v�(0*6���7�v�톮������G����3gNd6���<+�J����v�6B~9�ǳZ�r}f�a}�~�A|!�i��(g:�	�חKz�L�s��,�V`��%r�)�����&�h�\[/��1�o�7���їH�;�ޮ��SB�;®���Y�tX�/ub�\N��n�m��wr3}]?�n�&��'���kYs?��5kc˶���
�Z.�ûY�C.K9ul2A��a�C.�������w~��]P��?��+�e�Ez ��U����*n�q����HxO�'#O4L%�ƃ4m�`�H��.I��H&jdjëa��G������(��y�.j�
�⇸"WD�DS���YS�� ������mz$W�&h��@�J�f��d�X��k��om��T��|��&YԩZ Bk�����Ȥ��j�_wǎi����>D9*��(&�����ﴙɑ�������z�� � t�![�Ƴ��۝��r��WK��k��R����]�Z���moV7�
��Aݷ1=|1=�0�ֶ�@�{:�*�1N0B���G����m5�5����8Dm�/u���<�(����w�g�~l��Pv�ٓd;�Tm�6h����Cخb�<o_|� '���r	c���1HFG�A�e7��>
���?v��G��X�DP�p�<2�06���}ee;ӭt=��;w�/0v�WuhYଳk9*����cO��x�@H�A1;�2��*p����_}~�}��W1����1�R8rr<��Ci�֞��X�ܹw/�>x���Ġބ!���������0��6m����\u&ƫeЎm�33�R�"�����˗k��]�GN�6]�S=n���c�d��SQ|��j��� Ϟ20���R�����Q�y��7�ﴯ��&[�I���h;B�[�Aȳ9ֲ��J�}�Q��?o������%F0|:�<21�m;��0x�z����_/ڗ��)8��xt��)�i8������R����)c
�I�M;�nw��U��uV�{��&^�.�����f���WG�t�WuXwp\�1�<�f�HX�'����m�����HG94v��e�-=��s��v�]Є��,S�;�@�|�j|.Q����A�Ҡ΁Q�^�ȓk��A�Ԛ
E�#֮/�s`Z��q������o>������ ��{���\��+������,Ҿ��y���2�`���|?�����:�y��uqC�;M���ΑU.��BY�!���qF�p��Ϸ�>x�}���q$�8j��)E���ണ�?<Lv��K/L����r�����KG��<땺����F�SBG�9���L�n^� 9�c�]^�G��ŋ�
a::<l�o;]N�t$�3ײ�<:l����8�E��)�N#�������~�����pz����C�� }�j���Tlb,����Bkү#��.8"��f=M^����X��H|�A�����5��r��O>i�޼]��W����vgc#;l.ã�����k���$|5]R7�o�v$�c�:�['�u����#Lc\x��S��ϿȮ���y�b?��������Q'g�y��&�x��}}����#������׎./+�Ww��ݶ�b�-=A�A��%O�I�c�I{�����-<�14�j�Ҡ���0I�~A����F�q���:�O�D���/�h;>�rWK��~�ƅ��O����~��ÛU�ٱ�PY�M~�K��
�st�ƽp�r����)��硫�Yg���v�:"ae��:�'�1���=�r�M��b��XO;����[����/�w��'"���<��q|��M�������v���6����7�e�r���#}��{��3.^���}�Qⷛ�|jS�Qr�Y�q�*#��	ڐ:fζ�@�G����h��T��������9e�#\���'�w<�=���}�Y������ވu�������y����ѫ��z�s�P�:[��2�d�4���������4�svz�Mg�r������������ۿ�S����qd^G�����mqn�ͻ���4E���ah���33:��mc{	{s���ؾ���v��\�wMr[����o���ᡇ9?~����.!Ko\��\���a�K�v�N��W.?�Np�N����������d�nS��^��,7���ݼf
�f�rpg�Pc�K��衃&vT*��	�:�ng�V��*���u�Î=g+`s���3�L�;GG}�Û�G�`a��N�3��(�i���ґr0'N:Dg�飦w��S[)���N��9lG�Ι�8�=73G��A��XsƉ��|�i�|E���齞W�t�K��8�:[�ԗ�z�d�֚,�m�1tw�v�d��.�X�F�̫�y����XIǞ��4R��M/�C|��@E���t�NW���#F�
:�W'�9�z�~��M�e���!;	�����c��oC8�E��c�8�|A���Cu$D���5:�(�҅���wnf�~���=Ơס��_������>O/�^�Z��M��JeE�BD�{�ݡ��sp���!/�8���?�v;]w|r�������̃6o���ͩ\�޼�p��Y�۷��6�̝F�h��� 1P�I�4��)��ç9O���'qwW�Q��mn����g,^-�d��Ν�����h�>����661,���a��i�����������ּ�m�O�]�pz����#wa���2���#��#�0������?��1���)��)b{rt m�ۯ���k�=ꦱ'��-���g��K'|n�o:a��	�N��=p�T�7wM�#�NMr�k���� �@�P7{��{G؃�H@�ꁒ+�����򛻩�#���~�όJ��>���{(��rܼ�q�����1����)�,k8���W��ha<�����_�����N�S�i&/��g��߳�^_u�Nq��n�,M;Uѭ�=�	��l�j-��!Λd�u����us���8��_����[�n�E[z����x�/�WK~;
�rG=<�-�ݬ�F,8t
�K|�Ӭ���kϕ�'eT!n�J㘲V����4ݼ{pY=�n2�ܹ��yw����LQ6����i���k�֭��G�q���~Ҿ���9�m����+�Ti5b�C�#.�}����}p��#�y���Z;:n/-�d�������q$\�xX�Ϊ
��]v*�m;��J݊��⼽߾�=w�Bi�ކ��?�ȵ�4
C���;�;�%��g>�;ʹf�݁��N,w�|��5��~{��/�����^�ꍌ)o;���T��C1�1N��n6��+�8�CM��8�߹]G�q���ƨ��u��:Z���5; ]�9�~�������L�
(�e�i0��4i�܃��<}�S�:�����a�4�2�@>TY��ᣇ�6�>���G�*�U6��@��j�^zF�#��<�۵6�����I88�=0nwi��ҺK�ƽ�\h0/]ڻl��F�[s?�f�Ӟ�wg�ƶFdP�SoaV&:Z莡�iS�e>��(#ln�s�?n.���e�j:v��[no�W��.�t�ԣ��?ϝ⽶֜~����[+���uI+���x�&��9���$��z�O�-���^�dzơ�n��INQ���e�y��f�Ws�=���ܱӎa7D����{��࣏��[���#�n:ၵ�����ɍ�C�sksi���t��Ny�J�7;D��s�rzXn[��Ŗ����ǽ�ŗ_�ϐ����m�vX�|w��:U}g{����E�ׯ��8y�-i��<�r
�kjqy��E�g�ex�ы);�q}�_]��bnF�FbnV�9���Δ����]��c>f��#��ʯά��q�F����zn@���o�Cs/��Y�,��uÎl��܄���x/C�[1�ȩM���=t�:<lGÏ���A��qSN�~]����L:pt�m�v���C�Ud�s�Ğ|�ݛ8M3�X�c��e��X�ti�Mt�����q��y��q=�j� ~�o����Q��=~���}��q:�8y���u�H�9�/���OF܁��.�fMΞ?n�e���"]6�@I9=O�]Y���#޵��p�a�� ��_��q�pl��#�`٦��O �L��8`3_���HK�pইC@�_z�)�&6�(�x�F��?1asc�Zu�(�	�-�&�l�e�i���i�C���u�?����q�4�0�d��}%R�ƛ��ho�#Y��\!�bA�����Ѣ٣$�dA:E"�F�t2�W*b \/W9�7��J�E���)�Q��hY�Ya+� �2=����WH�	���(�AE�i�ۆ��<K�mdδuǩ[����0���ܺq������N�=/0<Q�7��,�j�Li̯�XA�x�#������(����Q��8N�s��N�s��5X��`�0��|���\cc�3�Huݕ�5��Uցy�pr�CE�B#H�X'A�������\F�Re��L��.W�6�s�u�<g�10k��y?z�"�8�38�`����F�������}�+�t�ě�u{<:=�n�R��S�]��tG�<������"{j,��r�7��)h�yB:�~�ݩ�:p�v�3��s?Ne�}}[J~�0�\��=��k��U����`>:�/m+�����(M�f��o��{w1�:M�E��#k�ۆ:%봏STV:;
�{wݵG��Q��N�#��m��.��V��r�bׇ��x�pK�~�ӥ����iR��=�N*�Ɲ���ә��;8�ޥ��3�������6�隞��U���TR��������Nb*E�*2{�u�2�g��3�:C/5ؠ�n��)�Ғt�<�N������=��w�N�q׶{w�dT��A�l��/�oo�ӛQ��hc�j�țwp��M�G�k�F�T�{�s�U8�2e���TQR<;]��GN|�wj�6\E�̩8uf�(,G�t�?�����_��}����[�.h�_qw�n�9��j\j8(G�{Sd:�:�
6;r��XW7A��эa0�޺y9���8:�"�.�B���B����ԑ����Zץ���Y�^��n��a��&k������]y7�P�9ʬ"Q�#ڣ/���*;�}95��g\�B9;D^����rZLj8�ӣ'�Q��)�uF�a	�(������e���[8�c<��Վv Z��K��)<��7��7�F:YB�P6��N���t�:��J3N4'{M�r:}�(���g�a���8���z��?(:O�lЮ:-�u��8F��C�}�Nij<�OwG��
���vq��Wu�F�]r��:�َQw}�q�F�� ���M�Pw�̽���>��w$��NK�W]h�ө]s��K�|���G�R���/�l_߾}�����"εK �2x�Do��N��M�Q�O��)�9#�o_�q��{'�iĻ�7;,~��lx077��b��X��<��ez��Ⱥ��8α�Y�Y�MһC��>t���ۅ�b��<������b�R9����sZ���h���Ҫ��ΐ����O|j[im���@�O�� ߿�����}�b)�!�ԋ��.���>v�b������Ѻ@pd#1�����O:���ώ4�uy�����j�i�zص;�J���Koߺ����-rs6�f76�1O���iK�).?��g7�q����q^=T޳�h3�R�w��
��:$\{��L����+ŵF�а;���u����w�_�����?n�x+t	dzxA���8gm�NO�^��C�ݤĥ	�~;k`kk�m ��ۻo�j��v�v�Rs��t`V�:�>Y�]y�����W�� ����5Qx����Y��>v�:��
�>���j����r]#�O9� 9��&��P��n�ȕ��ʶ�qtP�q4�F�,�@����F�� p�]�z'iG�Qw��F�V�n��Ծ>:ɲ�S8�H�|u������)ޙ���d~:���#e�ĭ�*����:�r���~�G8<X�8���2Ik�����8Y8�.Yѹ�vy�]X�k�2]:��f�����
�#Y�һ�
�L�/�/�|Br�ơ�� �{j$l���KE l75p~�C��F�H���1wi�4�&�:a"�Z�T��)|N�PX�]*X��im0��Ƅ�!�|Q��e8�д"А޽� D��|Ś���'����ъrws��u�׆dd��U�����W��N�؆�_�\htzb�C�N#�{�&��'�94N'#�m�:�vE�[^GAG�5��:Z.���@k���2~���8�L�#���~ �Sq�"�i�q�h{G��qdk��M,�م���.::F2���Sʑ ���77viG{��R�3ꥳ$��B=F;0ml�
#L
�,O!��=Q���y�`��w�4:K�c>�s�W�;w�#�`��q���[悧�I�t��_��O���:	:{���z�N�?D઄��#���Pg���<���:�����yV�ܹ{�}���8�Oq�\����a�(C�̤cni�:�B�Y|Hx
�M��p*	55��Q��5�S���w=u^E��=~�������HO�x�_1Xt�t�l˔�6]���Z�^:�ƃCG���FO�wN']:2�v#�:�Ҝ��ʀlr½�Cv��\>ӹҩҸ���(�Px��1mRN�˗:Ie��\�NjK!���hT�-�r�t�����N�ץy����#G�1�\c�r��6�0ng�N'C��A�Z�J����q蚒Mp*�Vd�F�# ��Ő�(P` C���C��P�.��ŵ�W����jμY������?�����n���oi����Vb��Ņl2��S�t&)����)����;C GNP��2���:U����~����,�3C͊lz��y��a���7�w�a�\Az4 �{h�ﴷ0�\ϠA�ȍ��;a�Ƀg�0�!�4���.r\ùF�t�ʘ��5�s?��K�}[������y�#��eNƫ0��u�/����_c¼lCu��*����oqGg���-fiÃdAS9��^B�<D?m�ܻ � ��3&ݍ�5�n�����ڨ3��S~^�9�����8VoaT9eKcM�=�E[�;�Y1��W7�q�ŝ��)�޺����n,�Qp�S#�����<�CV"4�S�?D���YŁ�����^�s��֝t*��Bcg����e)���f�@/ã[;�Ј�[Y�
��(�ڱe甲g9ƿ���?.e�(� �u��X�}FC�Z�� y@�|��w��V��r���8~���I3��c$�ӭ[�qv�cڗ�5���#����ӕ�,��m�G�=��=�[o��F1��sD'�M�� _��J��3�<\�C�:�3a��t��;����Z��A�8f:vJ�������h[;ڵnj�vt�]4��~�M��-���w�t-�t"�*�2�
:̮l;�!c�ӆn���q��w��.�jqz��#����<g���qiW�r}53]�ܹG�/R���Z��ř�����G���������(@��Sy�Μ�)w=^�ґy�/dm��rzG���7A�ƒ�G�a�)���N���{�r�jq�|���ǒ�L�ų��s/e8B��.׳�GC����Ƶ�����o�㮂�lIR8�$��l�ϝ!t�^�u�~�:��;]�ȲD��m���A����\z (=d�|��
�s﨔�j��&��:�������;yD'��ft�|;3�šδ�T�+�Yᮃ��H�s�����|��Z/K�N9�)���w7���Π����Ik��#\:K�pZ����a��:q��K���6�P��8���
��o���r��s��u��Ag+k�h�ӑ��.���9�I�!�	��(فK��\��a=>�уƁ��^ � ���B\R�VU�T2C� Mdi��̪iz�*�l�J�"K�2�,�����V�ˡL�%ӛN�g��~
����9��E�Yp=�0�_��é ۹�.�������p���X{�][~��u�U��C�,a��dz�,Fҋ�U�z{�j#ø2�����,N�y��k��7�8�V�d~.!�_gC�V������9���9�
�l��hcI�z���5Z���@���^�	pF��[��8v���RӵQ����_f�)��]s�O�]��E�:/n�:B��#u����$#y8*��S�_'HG���^npk�g��L+܉@.��~�o*e�;D�4Y:�~��:��uqd���e���Bv�V�H���;�����5b���Ä��qFݹG��5^N�ۤ�1����)�t�\��q��;�M|C���:��(;��5|��s4E(�c�B��k��r��!F�N��Lϗ�#4'�F(�!0�7��P���ݥ��)�8=�Ò��s)�q(~�֝���:���S�4�l��ݩ�.�u
����3�<mO�2�ˎ����Ѳw��n�S(N�&8�-�&���O�������;ZA>�w��{u�K"��it�^�P���6�A/�� ��
��������N���Tq��p�ѳ�ŗw��;�S�O�����#̝f��q��Q��0e��Ʊ͘=1�'��YIǃ�tR�B%�%t�nk/_��������������^A�	{��ڹ�y��~��d/:]���nK?��y��0�s뭌Z������k�3 ?��{����Ltq�g[)ֳ+A�f'���_9��s
�m��B�:����j��}D�������B���y3����v6X�b�#{�_ٟ���ųe� ߁����1t�"
����!8$3��*�tDj:��	gz��VnP �ȇ�̗�F� ��5�yͷ��ݺÕ6����k�4`������T9m�Fgס��8U����4,ݵ�7p,ߩp:{�?o"�j-��t��U�K�p�Mю�*�_�� :�D�k]�4q��\���k�.]Xl7n\�q~�}�Ïrp�{�Ӯ8�T�V�Sy2�}���8>��"�݇����Ϣ������ĥ8�G�ir*�:��+�{14���)�NG��dzw4F�fo~FE&ƹ�w�liU��ɧ4?-!��v�vʁ�.��Z�ߺd�1?a��K7E���<�o
>�9��*@;�7�az�]���W��7�H����(��zݥύr���<H{�����)�NS�!��D���3t�=G�����`gl#M.ζ��U�:��ZF_f�kk�I�af�����<v�$�U)��C�e�;�v��[�G'�<����p��=�U�Y�~ �����TT>�US�D\����[�3G�4N�S��:��xu��i��R��ͽ�%v�mM;<��y�J���o?����~�Ad�;�:��j��9������͛ql���5w����ȉ	�#W\3�>�w�a�(w�?{��_�`���5<��n�fu���pDG2r�����)����hV�쬆#���o��vʠS0k�/1��]��f�9��w��i�}q��tC�T'���K�8d��)����+��1��緱�ht�k��Qbτ1�L�uM�by�cEt`�?�Љ��T�ɾ'� ���u������H��ҔE�i����6y�uGkd)x#���r,_�Ȳd�e8�!:�}yƍ�G9�A��G�
n�g�����܌����r3:�x��)|�W�Ӵ���*����.���3S<S����R�r�v���C<vG�U�?(��H�I�,H�E^ޅ�z�z��z���:XqPV>�����أ��d�Y��i6b���YҨ�+�r	�^�[�V`��qBt�Pz"\,�������:�(��h�y��S $�AkoօE�]��P��x��{�_%�z��8��aT	Z�x 6:��5E�'H���	�.l̎���T%�ib�4]�6]ʆ8���E�0epklk����4���7�I�9$�(��@��8RI"\=4ϩ�ƵW�t~W��|�FM)%�v�a1N�F�]úO��� �Nن���N���s]�VgY�H@2�����et�9�:X]]�o�Q��r$�e����ߴ��\󖩭��d^�����(
���ar�$īv�����}\�g�a@�~Ϛ<�#O>+�'&꼊r2�I}��,!�,��9t�����t�4�pZyf�=�Fޝm{��t��&󊃅 /�]�ٕ��M\I�N������y�쓎�T�Қ�pQ����#>��]ȑ OAXA�=92�1<�M~t�Y>UتL" �P�䌸!{���[�&mU�Nxa;��>댊3���e���� Ϸ�~�}��١�5D���a��t��_�mw�?��Ѻ�:�RaPk��8�%�\X��.]�sF#��S;=L+?��\�����N�m���۽���\���m�����ޝG�Xt�Žm�L��s����8��rT�*7Z�/gA��wމ���ƭ���[o݈st�w�/S�P��%}�>�ͬ�����e���%��S����E��~�7?h�?n?�ɏ0�ޏ�㎦�L��S����`�s>�4��ЁU7��Јt
uu�]��giMc��/^�`�m~������ȞL�:�����)� ܁6�� h۠|u��W҆�!tҮb]����Z����l׬#�C�H�5�]G�>��85�o\OϺk� =��I����\#�zW��9�v',�P�N��|Ҹ�L���v��۴�#UN�r�g�$y�����\y���i���\�I޵u���h;U����i_��^ oo��^;G��Yo�B�� z��:��.\i�.{8��Ж[�������נչ8b���|���h�M��F������5�\��~��e��!��{��Q;*ÔA%������^�-��֐t��t�o��R��t\Gt��6�����N���A{��?�"������n�3e{9׏�<�Qq=�*tg'����7҇����Ƿ�.B>�u��2��w'�����N�u��Q�f��5����)��p��V.
�Μ�2v@9�t�䢓׶�k�u�]��Lge��#<�5Z��������;�}����ܕҩ�Ҡ#宵u����'������Ip�]�Z���Y�	�GĿ�I�|u�]���.` �/����\<t���v�ͻ;�����{헿�}�կ~����g����`:=݀�%N�S��Q������LW��8֡ȵ��ݼ~��8:�h�+��1�z����_~�~��/گ�U���i:�c�mi�����r��B��m�4���}�%N��VԻ�4�Y�������^�]�ޢ)�\\��B:���';�sy������`�&��B�:F����;8Rq�<�w��W�s�b:���{33�i%R���}��y���2�~6z�"���T��C'˴'����]y����C:YvR��`�d-�+�c�9��dm����;'g�iE�F�B��a����YVX��9�Yr$� Q�!Q|!*��J��J�?��=�e�j��|���jx�� ���b�)!���\>�.�i�f� �t!*3��Ȕ�O&�Q��y���{ �� ��a��Eۋ��	��"Wړ�o�;�m`������$Jr|�Qh0�8�����<8B�}l�m4���;�/���-ou5�s)"�mn�Ǚsq_�ӷw�����p�b c��4;d<!:>Ni�܇���8GY"�qN5�2T����[8
#���(m�r�u�M����ЁĬ�xq�C�4���Q�_.��w����+�ҋ�[a��1�®��Ut��`�v�_�U���ң0�`�\⎒�^itβƵ=�ҙ����2�1�F{�Up���W�4��/ڧ>ĝE�{��;Ey6��<���x�^���ť�iCk�s�%eG�`�����F���|h�s�m�_E��PX�cҎ4�BtDW���me|34����;��s9N�ڮ��|dOUz����QW��n�GNd
�{���s�m��ϖ��1h���/�о��x3r�݅3��I ����mwx�6?Ɵ��k�n������L�s�~D	u��)oeu��{�}����s�(�FwMҩt<S&�B�-���"� �����BGRah�JVg�u'����������W��������L�����)�,�p�@:*H]m	_�=J��2����"��G�H����y���(��K0R��;����Sc�|݆�mms�e��7�������t^G�5h��g�{�}��ۿ���������0�h�ML*o���,��20<^��r�j���#l��98"�Lu�����\�c��#?~Sy)S�稟k4."s���P�R��E�1���lu객�+k��;G�[y��?�)��;J&���8N���Җ�i`#�N��!k��y~�{8Wn���u���{�3ou��J��Ri����)�&�Yf�zuj8}�ݻ��_Hb2`Q�9:p���.���p��v�����yog��`2�
?�c�n����oj�ӽ��4��W?�K9��,������@K8W�^G�q�>�޻ܝ6z�n����_��G��P�z�U?��{:[���t��<�{����ȓ<�I)����Gݝ��`i�P�)3�)�">}6��w#��յ�1;����pF���ߎ�.�θ�TG�����.����yv8�s>��T��w�e��g]�8�ТzRݬ����6��~�  ��IDATY�c��� ��?=�a��r�:rgxuB� �t�Z�x�:rd�b��IӒm�{���֎&iL�uz�����nz�w�n����T]�����Yӎ��D�ϑ,�em1;�u�vw�b�(x�x w�v:��˗�Yí��i�:����mw���<z��N���
�&Q�;:�e϶c��� .@ѿe-88eҊ#�����7�_��7	_|�Md�2��N�̿v=���<�JY2�/�Q;���2]]�eG�6+m��49=M=��.��9�"�������%��|���� _�����i[Y�m�i���&:��@;���~{N�/���~�����>2D[Dg����P��9M��Hm#`��.m���tE�8L�s�'�t���'��\rq3_�e�-w��\to�{�kl��6A��8h�c���,%��|��'啓߂`$˱�NU�m9�M�Q6��9��劜	�`S��v��NO�\��u'k�d���dm����� ��HV�d��P�W�_vvT(S9C��p�Ɣ;�X�1�)�MZ��n��*�z��>�h0"l�ʈpӅw�]��56k���W�{�j�S�6^�)w�I���q�(G�ʃ5������:3��f�u�w������JqB_k�[p�
F��Ta⶧2�F������tFTn���W��.=ެ�q{E�=B-Fgox� �@{\�U�&N���d�[M��s���֖5mb��/�y��/l���v�sA�K =a�g��itfLc�]��G ���X�I�L|�ƈN�iN�tkx���K�c��g޻��	��J��Bu4ϯ��B�g=���\S�>-��҄v�[Fτ�ůu�iԨ�]e�����5�m�(U�8��w�IK�&)V#��^���0FIFr�	�H���/i�iI�h��Wij 8�$�t@��N���6m��*(mG��w���
F��N�8(����Pp���:�h�q`Ҹz�[�!�U9P��'��s?Eu������[7ٙĀ��n޼����5�U�KKkO�W_?jO����20��8%P�����}��R'w~�9����x�(޶���&�5�!�����
�>��7�K�k�T�v�xމ�|4DaԘ�w%��ncX�oLCXZ6����b���AI�gҨ�.�Y���c�A�mm� c��Q��;�g��9���N�����=׾����?�׿k�|�Q�vm�ҙ�.�n �\�^��ʵ&�S����S�W2��ܾs�����Hӱĳ8oҟ�F�(������N��=R΂n������`,�rJ��mG��+�T�4���Y'��#:7?���;k�4(�uA�f�1��О��q��;�`9MN#�雇�ܯ@�txq�Ёɥ�Ѐ�-7�u#ZP���]�˳����JҶf'�ul�uBң#.8�msv�cT�2j��rR��H�����\[F?k��Mֶj|���;��<�n;{;�Q��[2d�o��::i�q�g=l�p ,�e���){z�p\���8j��J�Fk�[~��K�s�«%'�=u/��t�2��g�2}��ֽOGef~����<*?��(q�g�y���*��48���g��5	lV�Y���N:�x��6�ƞ-��юz�K�����:�	!(�K����'N�sz��m4���\��j�)�����gܜ��J�q`ǎ���:_�P-�y�]�*��-B����?�����6Q]��I�ܹ�ܤɣi�͡���g�����\y�^'S�qwEG��/^�����?���V��^Ox���w�����}n�
�_�N/i�v��Uv��NQ�Ŝ9I��cK�A�=��ٲA���U����}������'Y`]�9�t_3�mަ�����T�,������G����sh��i��^H���N�����Hs��o�%�;Y����#��6�4��k�{�d�H�	r�Σ�z�o�Y�N1aV���$d������0���؉]��?��J�\�F{�t���-)qī�7�r��f𪼍[������+�)�ˋ�ƽ�Ų�\��w���;.|����I,?e�֧�#�w��b�C�Ρ�R�\�?��H����l$�su㊻vN�6���o���u��z��t�`���1LKn����dM�������e�8X��DVF�`��(�b��((0|Wx�ANU<�t��8XPL�0*�BT�YiD���FQpN=s�b�?�F�z�X����e���!��,C*��s�ů�h#!{�ϓ��ۓgoPګm� LS�BՅĮ�R8�A�qt�\����q��w8�_�􊐇x�)peC�p�6�?�U�������c�'ړGQy�����:̶�A���,��%�uAp���#~���aó���upn�\�ց�������n9Dr�>�:5aLpdݽ[�y	C�A�l7B��?�G��Q^9Xӡ�?���O�ԇ�i�/1�u �sjA�*�#X̟�,���x�֣�e�]��`��,0d���3k��Q0Mގc�S*h7 v��rz�O[�ls��A�Py��ao�mw
kR�*$G���r�xO�.�Cwn(8=H�@�Q�9���͵:V9H�ߢ©rq�hHqi���7+a�p,%��,=�1��н�>��.B����E��5*E;#��A��D���pf�]�8�]����}�Yj|���ۏ���%|�����wW���Q�Q�e*�up=[F���M��!���������sm�#X���vws�������V�C�4���'�M�bg�施�e�yX�S}ܺ�Q��Bi��n$�u�;(���F����.��J6���������e-�;]�éVʟ��i��A��ڍ��0���t�jL%���z{(�j��u�	Lي�-�-�փ��]�Pz�q�5�M��<�<�:�~:ĥʶ�����NF��ذgRm+�8�n,��ysßM�<��d�g�B�a�����h:Mp�&p��b�Z+&�Ϻe�z1��);*�#;.����~c�������v:�@���2��=Pީ��Mՙ�W2e� �+>Y���
��F�ҞE��O��X#+��ւ:J��ڧ�~��<ȃ��7����Ne{-�e3�=�yU�v��_�ɑz��Cv3�]����ރ�͝TMZ�(���t�P�#X����?t�Jv����WV��:'��w�����{�`��.y0D֪��9V���#���p7]�l;�mP�WJ� �P�v:���|'79q��/���<�õ�u���@��%3 ^��͍�v�SD#�lV��-�;���e\��
9�8v*�6�
���O_����'�U$��ږKpM���6�i~5�⮤:Y�]7-�����QrV��)�c�4�\Yos�k���l�0#뙺:K�ȱ�t�,�Dy
|o���v���v��Ed���g2�ڻ��k��R�PI���/�4s�d����|{����ܿ���3��ݐ�F,O�i*�ѐ5<>��ciE��)��hB�V{���Qd��k�32����*�9��n൷7������}��m����pD����6�΢S|]���?�u����u�կ>�lv���2�!��1��R�����8��J�Uol+�C��Uɐ�\�K��H>�V~1���đغ+z>�Ի��.OJ�w�'�~t����F�s�9��2��\0��,U��\etQ���\�W���.�R���^*�K�7ku��Ϸ�W.d��[�g�������L�v� <�DKP��Wf��c�d�y���h8kPj\�R��$�(s+��4�5Ɯ����J�`�c������[�����WB��[��{	Ab���Օ|I��l��)��C�F����8��0�|{[�%ȃ)�߸�\�����܊�ݑV���VJ6Z�_��u,l����;�.A+��� I�X��x੦g�ϙz��}⠉q�w�j��o�o}u84�M�1b[�a�L�p1]Bz��᩼k�Z�QL���F�:N�p2qU('#=�O��c�~��2�ict�i��hw��������
��wU/;��ډ����:�;p&.��Rh��C�ƔF��{�3NQG_>����w�W��FT*��<h/�]^jN�����9k�U�<B�GhC�:R�+�
K/7�:����(/@a��s�����*O�-OpM���b>�]}̳�W�>�H\� ���N:���*�ՠ�v����E��T���dM���_�׏�Jq��Ag\h��.����A
MJ������C	m/�#~�S�8ZF�(��:�E��;{@����2e$=�N�U&�V���u ��A�XDA�������oV������1_���Js;|w"�����o~�N���1�$j ��H���e `�d��D�h�ު]�wk�/�]'cQlnlęq�hͩZȥ]iH>��Ts1�el�c<�䈊����ڧ����|E]�7�m�P�9w��[o]JG��X�S�\(׹J[��oῙ��N�˚��y�k�֩������
m� M�� T6xO�3)c��Y[�X�3���)�1��ӻ�c�ݡ=_���n�n�E��)���������9;��cG�Q[~��mo�G�)?l��L��cG�����}@��m+;^�^;��i��EN[����/�O�U��T̕Mx�^Y���י�ISQ�v�ȶ��7��/3BL���8Fv����\¦!���qȉ��U�	��6ރ���Kw��n��7� ��qv�t�
۷Fx��5ň4�C	F.�����*x���y��~�j�yn�=�$_כ��v�D	��PX���8Yi��t`uih�������^�u�M��5N�K�;Ȩ�i�E���,pe�ƻ���Dl�g�s�ӫ�7�2�c]�Gpg_۽?�T>|�xN��o�d�Vsd��A�� �Bs�
�:�����;�����Yln\�����v�(F1�*}�ٖۭ{|���OiO���[�L�we�a�7�!_ԗ���o�N7ux���f;!�Sěp�L������I���3�ա�1�.��K֠Aw��gCY#��kk�� ���e�>�&&��7Zq͖#i�k�*�n�ﵭp�����ES^:9v8���_~�M���&���9�!K �f�d;-�q����u�R�
?���ʪg@n���IxK�����3���^"�?}�<nƣv�=�Sd���݃GO���olb*�/���ء��v؁��W��'���_������`�� "�Y��Σ�Lh>�Zjtp^S�pr�qu����%���C�k���e�iW�|W���g���=b���ґ�d&�F>����O2�;�Hg�A��+޴*C��qv�u�w�'y�:�4Bb3�޸�w^U���-|A~��e��ߴ����,���H��N��������
}���̍����$1"p��W*��L�dU�1�a+�eoOz׹k�� YVd�h����]F�Sj��Fd	����&����CM�1H8��#?ன
�N�4�c�ڃ���@D&����/��:
"Q�Ef����~�B��'�~�|�ka���x���^���f���h�E���H�8�D�k5��\!�G��� 8�0a�j|֙)�����z������o/Mg]%��v�KY_qL'��A7r����Zo�%�4��!3b��Q�S׵=�9UgHE�s�5�H#�SCubā�06ߌ�Z�(E	Y���¤P�S�����v�[��z(	�:�@�B��$��%AȨ�{&j{��Y�AQa����ѻ�� q��uΆ�}ViTZ�|�ѧ�nE��con�F��LFS��#h� ���ĩu&��d�� �1m�F�q�����8|�c6���|*��T�k��x���pB����1\;�i��������f*�%
ҷ�K��8�L�c;]��n02p�K'Ɍ7�� �?�N�M/��x��F�=���=q��i�����;pj8*��y�I����K��6���:��{)+�^nǔ;3���]��&gf�!�}���oo����F�J��ɢh���htժ]9=����T���z�zcuE���.c<E��i�GI*K\@���tD���U���=�GQ��2%�v��~�WG�֘�R�c@<{�a�ƅ�Cmsw ���XmO�1�]��f1�;0<��i.�8r�[8#���G����C��1���ܱ�v�6w�������9vG��!���q�T��X��ሠG ,�n:q��?o�ű��_~�C�M{�����3G5&i�!x���9�nj���V&�ɗ��9�8k����$!�߷�ǡ�����JF#���>��S�� ��
��!�k�5G_��t4@Ñw�V&�j=y�_��
�Q�:m;�8�N+�`\�k���f�9~���4���&���x��FeP��~�#�w�縻�=�:~E�NiŠ�m^��&_`$�I�S��2�Q���r�PgO�`d����?�@�/��i��is����d��%h|�f�=�m�{`:0��9�v��88%+֨�;�yΟGA V��699�nim}��eҿ$�%����,���_dm�7���A��?kK���M2�^�u�:j�V��i����GsE�y��ߕqW���=u[�?� �2\;�G�o*�ݳr��S��l����#��CGip26��3p��Q�G��q{��%�6h�����B��@W���!A����Sv�tx���~X�,��1��Zd��ȥr��TF:�O�83P���-��+w��i�Ι�/�	�=�Mtы���������8Z�����Ό�T�i'!ˇT:�};"����6wu�2�<x�����<;�����o�z�׷:?JJO*�&wv<jţX<��s��/�w��`c�mgL�;����n4Ͼ��H��;����8�:��a�����B[X�#G���pD���{�N��B�M�����(��@^P�k�Ch;�t4�_�,MZg��A�9�����:�k3���Ѷ�5��,�.�v�yv彻/ۃ�����K��n��t*��/�_�3"�\��<��A&�`I�;�a�/��l��~�>��;�z�6��LF@�4 pB�����^�[�jl\{�N,�Y8	��c�j�Gm�9]�OFqz��7\!.�������b_�OqL�ߎ��q�X�S=���ҏSٗ�[yֿ��t���i(	<H��Ծ҆��A|�e@;��T���v��e�I?��y]����-r�l���)g��΢�L���#?u��^XlW�A�o��^��j?����?~�i�5J�9�wc� �8Y@��)��tAO��[�1�p_����#{x��&C��Q��)�����\(,i�<_Ear ��\�e޹��Р���!N�U����5�-D������%x}��^%��*ã�$�	�t��HC�n��]���v�4,�϶������/�~��G���K0��yo�_��������@��&
&�*$[���
�j�VChd�@~w�N.�I��G��B�q�-�~7���kS�W�p��gq�2,[Bs��Nf��Ѥ������Uh����e���a�)�lG�}�^��Hk��5@��g�8=<רi(�6{Z�~v*�`{����E|Ȝ���t
PFz���c`��.i|�Fh8%�42d9a֝����TpR����0�SX���M���iI|r�hV�d#��|W�jP �#Q����Gyc]�V�'�)�t��mT*�
g�5������|B���㸙�����n'ktR��ʞ{����Kr-
�k^qڨ�EDd�-x�����%�5`��ҫº[#UEHQV]��iuʢL�"�^��?l�����w׀�j�#��A���!qx�.g+���j�������o����3]�mt��߷���Y/��(7�1_�
�Q�R��[EG�=x�P���ɶx~��q7�������:�R�3��7:k(,��~�����:��"_�!M=<r:"F�=�T�kw8sc��v/�^>;�F8=?���Ͷ�����(�fGL�=��; O�l�� V����H?���n����n�{�m�/abp>%��}�P�@�M��|��_��{���/ܲ�-������Z7�M�>��?0��M�R�1���q��l@����v+�Wod����t _<,�8;B/E����Os���)���fN#��j��d�螛�o���m����i����7v�D��^��|�L����(:]�-�!�6�Q	�����x9�Eg��KϷ�-��Õ����Rg�y���V���Z[IG��ϵ���j��裬C�whO�n�������m?#�F�iU�Z�9B��}��N�D�p~��s�����kW����1�-����M�_��y���;R��cD���@�9p����t��P������)�K��R ��F�˖��ŐW'b�����Z���Y�ǟ�� 7O9�#Є���]�vW&ˋ�{�p Mg�[�O�I��D�N1U��o��MG���ʫW�4��|u4�9e��hۡ�mni���-��0�ܔ�Nj^�q�gm����+�.���=J�3�槧��v�R�U'���q���W:cxp�2�Wg�=�I�Ɏ(�	��gǉUG7���<:>5��6L���k�tP�)��@�G��y� ࡥԩ6�pʠzTG��{�)�g��KN-�C�M5;?Ğ�8g(�<Dxjb��h����_s��<3����LK�v|�-m�g�8�8kn��&'�p{H�����܇q^�G<{��t�j8��[�Yp�n��>j�O��n�ho_���Q4Zۂ�<pۃ�����8�� �F{��:4�n��(����Q�4�������1�;77L���&N�붹��15�m�vNE����8::K��4�]5��yd���NmmG|�7�8ǎ;m"٨��h�j��6�)�e��FYfG��ș����Q_h[ʬ:G���]�.�<�B��K��\���'�K�����Ĵ,�klK�HP���D�@�B��ݼ'���>�h+�;x��3eR9��I�y�s��}t�4�����?|�������w��\mӣ�������'�.N�Z[ߑ�a4�Ue.�a�e�����R��X�(�ݐi��E�E�Ҫ�0F���'��;aEU�u�i��9
4��"�Sq��v�|
x�C�d�F�m�x� WP ��]w�1O3��ߥ��)cz�͢$�mI����U�\��8h�����[7ڿ������?n�{���"p����n�կ�l���������a��88��\9}o�k��{�_���S���C(c�<=.�I<�� O�����5MK��C���i������<�vY��u�d�SK4�L�=�k��t�,ǭl-Ӽj*�v@ث\��)Eg������|,<Į<2��X�)��O�q�~fڝx<�C~��ޫ�_�}6������)<��
�j�"���鑤'i�� ��+��3oFi��r��p����P٢�Tlfc�Nߡ���!�����x����Lቼ���F�cu��;��͒�)lS�y�\�%OG-�)#:&�)0��;\��%/��S���C��O����"���N"ѥI�8S�F\��rȋ5B��LEn�4B�[+=q�����(ġ����x�އ~�L�1�?�}�!"D�d�r�C�7���H�+�>�׌+8��]m7n\k������������McȮ����~��_~�~A�曇�"2{��)mt�̣�:X�/�[f�L�Y��1�F˹��rd{�������d�=���q���U�8���w
.`���_2�hT�f'FɊ���)7g�8w1���Dd�g}�d-c��x��s�w�'�U�Y� :��t+�S���<�������68|���10��t�4+�t�3���4n%�tG4"/���A �0���<!�h){\��C��1q����P�L�3�0�GF�k������c�ea�DWW��B�kѓ��Ff6,�����Èv]�X{>�0r�A:��A6+w��u�bY�2�d��3N'��?G��5��pJNЯ����&}��{5�J/b\��N�n��S�q�3*�0
vqDm�[����'�~����v�\~u�i������?~Ѿ�ηv�	�ՈM�ߡ30�#�,	���ܕK���o��b�n�`�d�����u=Y�nḹcbGp�.mNTg��&;�hku�܄<s�6�(�2!�|K��X�7�˓�[^�w��s�ǟ��=)�giP�Q����;��4x�F��� u�n���iy
���=Ng?�;N�D�ǀ��Q�se�ċ *_2"E�u���d������2���C���ϭ��r��D����{ؽ�W � �sF�=�Vt�4+O��.񥼓��s�85U[l�&t��Qm�~���Je�xToH�Дv�VZ5��ܭ�5�|vq壝��s�Q:̚v�G�NJ�4��Ax�a�(��5v2�C�9b��A�۔���Tܽ�-����s��$+��yĀΛC��Á�d�;+�Y��Ҿ��h�66t��<�s�s7����SV�a��7o��
<��P�ڽ�nfgk�x�A�=�M:������٤>v�Q�r$� ����_G���F�fue"��!hB�!����LU�ZR��;eZ�
i[9��N �X�U_���!�� D�{/��8/�6;�T�U�Y�v��,g�wډS��}Y ��>�v�g=4�7����zC���o����ʺ�x+�Dϡ�h�p��3 �)��>���V��󞥌�i�UG:k��: ��8���J�8Y�o]���'���>��V������5�����?u���<yٞ;dA�Ֆ��IdL��d`�h�iP��4v*�, ��4Lz��Cj*C��:2�U�X�!���*ÿ���a���e�I۳�W�2x8I#�]Ceޕ���$~��� ����!�y4.5$h�bAg�F��Wۏ?�^���wڅ�cmT:G[��.V�.8O����j��8���l�;�=����ƭ�g�
5���8�~j��i����f��'�F�gZ��=�s6q�+��4�#���Θ8���J�D�;����L�Ŀ=:?�4�kә�maZ��$?d�]��^�4Ng�PA�՟�,Z���AF���:1�aB���J�g':d=��<�7���9�q�,	�X�Ο��p[��L ��`�cqM:����kqf�x�O��2�>jzqS�)�f���J;릀�v.c��YE97�s6���`���)��2j*b񁸪���{S��T�����he(F|8���|0���os�)� ���n&!�nn�զR��0p�oR`�����Y���9A^���/�2�:(��nW�:,*��q�������� ���s�v& ��Sׄ.^��Ƅ��:����kW�[���29)#���0��ZGS|�ܳ���+	�5���8�����VЕ�B��ٞ�r��?tj���l�L	��d�r��1�R�)��]��ʒ����44�?7Dp�r��qrQ�Ӓެ�Hm����H���k����2�ѫ��47���i��`��Ħu��߷�u�ݥ.���U{��iv�sڞ�,s�;���w�[��9�$[i6�]��v6�pȷ����y>  |S&�k�ӗ�QGB�6�T*gXf����P~��-�^~Ua����Q`�,�׈0m�l X7�p��&�]�����<�Gz��#f�ҹɃ���v���U�Q��o�@����Fk���:�îy���1r߬���_6װ<�>�9v���[�&��6���(��<�}��v�ڕ�o9<F� ���L_tSG�A�C���q��w�v�����}�����i{��C��e9�f;;re���n���b�J���`���,�:���]-^��w��)]p=$�{�f]�O��q���\�EjkiP�i����𺆦���%�pN�Ӟ�mڜ`�_�z^����+~�������S���B��,'૛rY3��(�����r�c|��Q�x�$M,�/�)ߑ�M�Wg�ye�e(�Jw�4���KG9��/���+#Ч#�q����t�� R?�p���e��S�a����Cu�G&�a�v�(�9N];�x�
_=sS�%�@�����d��4�o�[G��ZS�蝲ȳ�=z����t^��3�ۡ�8�M�!k+��ǰò^�����UR�{*u�3e]9\/�-�>T*�{9���E��\�Fr�0ʯ������g� �%���mG�A;�]������e:����ƶR���G{iw)?��r�z��35�s�((푶/���wj,�C['q���_�Y?��2��o��Q��NW�_:���v��յ���y�.��0�7�a�j_����)m�����'��s�7��A�LS'�8"%lڝ$XN�^-;�:)�o������-�Ż��!�u�A:3U�|�\��l�gq�G���;$����j�?�4�l�,N�&7���d�	*��&�&^�i�W�s^0��j����&�6�[iȴ�_�k�`x���x�1"�+��i�i����Q���wu'=qu%�1��T긌J��|��u���nj��^��UN�F�QAnCV�2�J�.Z��yÈ�1����K&�)�tXW�>�n�2�}����o�h%H~�^1x��+�uN�5m����	�}��!g5U#�����l��¤!d�2���J9*E�ʞe��dn3�97e� Gؓ�d#fZ��1��0��J���1ҩ#p(��T�U��6��+��KϮٳ�
P��#h\S�Ni>k��G�~����H/�F3��2Lgy����rR����ď�U�	��8�[�:g|qX�o�+�ROBS��x+dTE;�Cc���4���s$t~�M�-��O�_l����+�{�����6�p��;�-\��	<OΜo�S	���	�8a���4|v�#FY�)��N��u5��u(�q�¬��h�೻������BС�P����|&�h%	i7���^
���j��w��D���CNPa���w龣A�*Ȅ:�督_#�:�F���G�-��>��B�׵�c0Y>�S�_� �S嬷k'�o��]P���֔m�@�p@�{�U�v�P�N�ECCY�k\�`�׏�㼹��� v�u�Fx7\k�6�v�����ݧ��ۏۃG�K�8�:W*ԅ>:��9t��v%҃�i`�#���:Q�_8�ϭ�5�\�0�r�=��G��y9�4�S��v�,���D�0J����'�EY�T7�p-���(��e��ٻ�A~N?��:�GG�9�`3&����� �!�Evă�������gVy>�|g Gk7xs�Yw�u����>���f1��mE�?�θ;ii\�a�A��{C�8�Q� �K�;���aP�/뷊�⎗Oh�g���{���#ȿ�m���v�����~�>��ߵ��?����v��[��L��-��Q&�T@��-��;����|;B��L�?׉�gK�9�݊��zm��m�>��IBv���v,�5��mGH�+Ym�EhL�_���s���`<�j^��
������0Oy�/���Ԁ��M�3�$�t��iΣv�M��}�E�5����Vh���ݶ�C�����S:�3K���5*P��R�@��_��60�f���2�����KY#N5�_��������W8z�"�3�C����G; °k:��zEO�Tsw;�ey�9���<^S�D!3�߶��w� ��1�l�.h��"?�!|9�-���7i�1H��<+��G�9B�Xd��8h1�!=��Y ����mn�h�d�܋���k;5�'�ϩry��|�A}C�I?9��w�}����S� h�ڭ? >�Y��.ru��v{CY�kn�a�9JY���3����ygt_ݣ�]	�h[;9��uOy��0���Tm7�����e�#��8[��U��ؖڦ8:j��KٜeG���6RxI��y/S�v�Qt�bG	�x�}+]}�4�'�vi�*9�uv�e�<חe�Y�'A�k�ص�3ρ)eHtZ|��a����#��e�V ��V��q�x�e��#�r�ܗY7�T��G��}檌�"ff��D���x�8:D��FW�v��2V$�)��1c�W��g�:*n9 �'�ͻB��.�"��2�E�����p��M���Ǣ����Z���#��iҫv�/;��%-�q�M�= 5����Dւ��+��0Yn��8y���Џ����M�#�R��@�n��D%�p'`&e�
���p�1� �G$S�0!��e�?a)��]� qH��1��4��Q���Gu�T:Fq@�������FR0i,�9��$O��6��c��F�d}t I�1��[�� 3������J�Z3$>qR�{p&�y>���4�y�������61�a��y�92lʌt��v ���}�*&�84<�������l�
�#�-��Vӓ�sm�ܹ6�x��.\j3�}�M��3�_� �ئ.��ūmz�Z����66{��L_l#S�̹k8_7���y�U�]��s�:d7��K7���on�~�na�J����&q��0F{�lp�x��([]�LG�݅͞qx���:_R�M�G�� ^��z�6���8,\}�Ҳ3ss5m�NGH�m��L�1�9C\s�G�m�b�\���
�4G�������,%Y砡���訽ts������1JQNﴧ<t�?d��8W����P��U��q,ʂV���v�������&��{��0��덚����2W�"4��&{`�u9�"J��-[ǔ�H�����3�5�a1�>����wGS1�0t�DC�t��7<e�g���De������̍�n���b��uz%z��r��Ԝ!����[w�ά�ǧS�����@^<+�kC�B���s��#�Q����n<���:P����3���Ja����$t�����%/@S�cd͐��ȝ]hgsZ��k{���ā�'���׶`$ח.^�����ڏ��ۏ��?�������I���������o���o���)���"o�>|��ݿ�(Ӥ쌰D�Ri��\��ȕ�8�Aa��]���H��,Jw��Ʋt�@磓₶/v���}�$�g�{��&J@W�֪}s��������UgC�	���ʕ�yȏ�"�,�z? �8�N�����t�\��@���`�'�@��#�[gL�؟������Pp��,�kk�ci���5���#��i���N��ء]��L���"�[7g�� o[��K�4B>�vL�Ɉ3f|���r���p$�f)���]$��ua煭g;�ME�ǥ)#���(��N f�^ҩC"����/X]�X䣉���qg�7�EysH�op!�0��<�67%Κ-;Iƨ7�~\+(OIC��YqV(۩�vf�*�t���۶�\"��#zV߸���u�3�9W:���������z�:�ݬ���P�v�=��VvӲ��919M����4�L�-�b,�Ɍ%Bě�^�٪uזϨ��~�9a@�LV�0e�i�*?i[ʊ�;�I�#�s׶ɨeF�j��4�A�c�
W:�I+l�Y;��)؄�6�^�Z#�����V�r��M�ѽ��%|�3�tl�6�ā0BY�k���i��|ɿ��w�I}����<��b�[����E�;D��Sc���R�,1��$�ݼDց��*��4]���,�����)y��'Pxʊc�=SJ(ǆ�,�b��������^����dA;p7�[�U�@͏F&?�ɪ(�,*#c��4V*#��� E���h����EBU��7�l�Q�ip���1>}F�'nFU�S�.��K�ғ��
�Q���9 ��)���N���lӖ#n��@����R�u�i�|��@�����M�;�s�� nL[g(Ya6M��=���mo���6���x�-s�OG�r�k��F��(<2�el�T�5�`^�5���G����XE$\nP��� pQ7Ɗf}�8u���"mFulW�'*Ǭ��x�c��:%���j��"߃(5���: ��5�����T��kSs�8B:V���3��ad�|�ZĶ>�Fgx��5y�*�����ؼIs�`p��8�l�z�J�ɚ��f�o��ś���[���wp��m�.��.]����8Yo�x�p�t�fp���qg���TD}�l�r����hP� 4�2� N4��%(��Rp	��a�8�<���j��!��xa��w�n��BY�.��w����:B~���J�8c:��:0:Ђ��&��ك�P���dy��T���5"����r�� @�7Z�|����R*����o��%e��`z�ɏ<�b>�^4�bԌh�+�Ӏ➘r�
|#
��h��)�ʏ����F���+�B��A��R�P�F�#���mgZ������S�-���g��UO����G��@��C���hk��F)%m�G��H�b\ 3���(+�G�l��R	N{��A��iY٭�@��[��ֲT���M{���.5�\����!gm���u�\��:�pv�_uB��`�6�z�Aj���>�c�oa,y ���	����l����퓟������}��?n����v�[��ծ��V;�r���<:�N){��a��/ۧ��?}��c�U�/58tx��_�7��	v4�{�)���6�����Z!��^�q��5�{c�B�ڜ����u�5������Lg%��j%)���`�^5?�p��y���5;7��upy1��w�m�w��vwh3G��߶��qĳSL�>ġ���_�/�����@�y�A��e�G���#�l��D@��u��[�$`ր�uVt�t����yF�p�»�?"��a�joCUg��B��d��*/w��,����6#�<V�	��r�_��m��	�[Z�ybv�!u-Րp9Ep�r����͠lp��]E�ѭ�
ʋ�s:]FҨ���ߔ'9�N����rj��9�� a�}�Վ!�ӺN�u�YW����m/e�uTVQ����]L���M�o�i{���Et�#o���i�֛6K��U߁i����� w|�́?;���c,K�O$m�3�G��9�N�r;S��]����4������Y*�/�9��K@�$KFh7���"ʂ8>$�G�uꘝZG�l0/��i�۹oA��1;n�E<� ��Z�*�}/��N�,���%BY�o�ı��#R)�Rg+�e��)�۞AV��NW�۫�N/�r�(�N�
ZF�eu���������|�wQ����i�p�0�GO���7���9,r�y��	Qd(�q�5�(�#��6B�$)��m�M�#�����.���� ���"���ie-O��9@?J`^��u�JG�!?��3�1Ӄ\0,��L9¥�1
s�\
�u��;�d�q&�cjr#r>k4\�m��^A߹�$��߬��Ɋ�&+c�T�5J$��[p*�����r�w�w����R'sg͓�-��.`Xe�pVg�/���l��0Y/b~�����Ws�j��q<SG�I�����ڷ�a@����"k�uu�`������i0����룂�a�Q�@O�q^pM��vlk-�<vq��R7~P?{j�,w�ѩ�hKӜ0�q��ʉ���4��u��X[�S�qlSaT�R�8ёtdM�0����F22%�&� י�j��H�Q�j2��P�Iӈ����*lYcBn
�M�a
d�SƝ�����wZ�B{�	�{�3C8p��q�.�'�!�h�K#�ݥ�1�@= ���0�Kf���F���4�
N�%�k�j��T��� s����ԋ:p�qנ�nm�L?CYU��7�o�T�	��]e&O;�M,��ޅ�LN�F��95�)��a^.ƞ�k�s���1z�ƕvn^r=�땞��fN�=����E��k'�!�� h�

��;/�慲�{�$��O�l�X_����\��8�x�m�dO0y�SX4�#�z��ϝ
�I񁛹(ls6M)8 �j�����g���-:C��䩜�4���J}8m-�L/|Ҁ����o�Pv��Hr�:V��.:���r:#M֬�J��r�;;�YcYv<y��m��M�8�N���̫�3�35������(�(�#�|�]�=?�W?jZUܙ$�#gq�s��
X�).  �#���`���q*C�� x��w�'?��}�8V�����sȄ�637������L�(��5;�Kv����_�/���ݽ�0���X~�Q,�����u��$�f��Ձ'��+���N�.L=���W�Z�<Wc���/�tnB)6|)�gޚq.������ղҊy���;Rj���"����5���H��Y#͔A�׌"�O�j�:^�Ȼl����eР�;!��ܪ�P��C޵�BS�Y]�#�>�Ъ��/Ӡ��P�����ҟ�2T�$����.�)���I\�γ�!3-�wf-qy6������Ͳa�]�I���L��8-�w�ˎ1+� �������^Bc'�=�V��]x#jk3;>\��� ���XI�ٔW�}:^�R,��:<I��:��W��t��O} �퐵cV�.8#M"�6�#΍z�Ed�(,W�-�ù��w	Ԧ =�R~����+� |:gC��mk�`��Q�lP���������Җ�2}^����W/�u�X3��_pJ}��⌉���o6O: .z�4�xi����z����i9����J:[�鷂�p;�T<�7����eN��r�5^����Bۄ�yUGz�c|m��Ɋ�!N�w���a���ە����:'k�rMV9Yx�F�(s�W2'����*z#�QT*�1�={�(��I)�K��~�i�D)�қG:N/���#7�YT�g���x-o��m���Q�[���zD����;	:e/HYE�4$NV�CpV����	`0��4�5��;7�ϟks�s��1�#O�x��s?>~�sE앳"�4*`��� ���(�w�s���w�{����a�ġ� c�9�Q�S�u���i��h�vL0]	�rh�(�>�~����BG����2�$�8f�U��d(�%H1{�dZ��F�#��e�嘇�����A�q�!f�����̲eh뿻��,�_F��⮧�Tګa�� �Ih&8�e� i\�"DO�f��Y��vaP�P��գ��^(	��Rt��J�N h�%MO�6k���������=�*R�eۓ�.4V�eC��m����|���kcS�9+C�j�`�����\��t*�
�a���t�~{�Ӝt�p=����2��P�I�����1�3B��^�~��'d���+��{�T
Tڬ�q�J���%���Z�L�F	x��%B7��̽�g��Jn����gk8Yoݼ���Ѻq�R�������������=x�Q{�f�쀳�g���pR�u:�j�ʃ���G�5镉*�вpB��W�}G��#I�YY�*�ޛw_z^��pk*l*r�KI���sk�����8�[D���4=��uB���_��1&�>�m�?D�U�l�������=�*e�?4 }��^�(g�%�F��s9B)����#�,�-HP�7i�L%_��E�Җ[X�Go:e9��7\���%ͩ��ku�Q~�Nz�6�� �(��\	#�mB@�?����u�*4��U(;�O��p@�R���y��-h���>�������<2jV�t�e��#��y�ѣG��o�����ѓ�Ẏ�c��R9x� xOu���ӹ�SHz��)*+���+�9%�kZ��ɯ�m��;�({�މ;U�V�ۆК"��,��BO�g����O���{��pL]k:* wY�k1�c�R/�ɗ�N��q��"�6���}(SYh@B��}ۓ���}�	��>(
���f�A����4R��t���ʑ�'�j�A �C(H&W�=_�Kˈ���	�ꔩ�;ya�޵����XF�%�V~���-�1%�WB.	:T
e t#?_v"D��`y�]F����%��}@uu���R���Ѝ�����V�6V��Q�Z{��z�@��^�*��F��n��b��[�#O�dE�w�����qm�4���zXߌv�~�{���w��ۮvlG�i-�$Oa����Ē�j� �� �-��4I��T�Z�MI�L-GC�o?��L�-TXH�H���*k[:��L'Aj��X��m@��c��%�魣�lߢW;���R��L���g���m�w��ؤ:��B9������fa#��ph��o�;p�������w3�ql��s3�ʥ�l|qaa��,G�>]j/���F�`V�����i�#�u<2G]�5�P,�A����9t�Y�Z��Ґt~�Ʈ�Ɉ�(D$CZX.e��.¬�#"N����_pmCo9�K��/��,�Z�JPD�q�`��=�q*�G��4�O@�R���&fF�9{�J3���֖�7�`=y���j4΁��2r9M��x.Rp��jK�Ρ2�+����	�!l������*���嗣q�"�Q�`�&N���]#���K��c�oӈ/Gk�B%q�bOO[�>L�{
�]ě�o|�mm����r��\*m�hQ�Ndl�C�YWf�1��Q�]��^���.�5�2(�i�ǈ'��)�tŤ2�4V��6N��N�G�'tCYE�Tec ��IkO��f`a�N@��_(��]UrU�����%dN�>xЉә5MM1PP��.�O�����\`q��؄S�\���A-ӳviNwRr��T�/���􃚦�P���oP��PT�Z@�o<�S�@E�w�����x�5,Q����S�kpX���t�і�"�[��j�w>�\����_�{�Cy\:�@Uf��;8p4��t7ΫW.��޺ڮ]����I}��U��ot��?�.a�4Oۢ��0	�e�/@� �!����ށ>�C��d�|�@�E`=�7�䝪S��A�g���"�X*o	 �h^����~,mC0�8|�Yp9V�M��S�)�^��'WJ#�u���]>C��>���xȸ�2-�ąu�9�bd3�0`�K�� ;z݃3=֔?����v�3����M3���t�����A�N�i)ڪ)T���Ѭ�A]rN��z�_)f�DŠ&�t&v�Q؏�#��7pXe��z�LCm?7夗�#a$T�euʵ��(��K�Ϸw߻��}�]�K�!p(h�<8��(S�n�����_�_�����W���'/���Vx�vń��x�ړ*vV�'����U'�#g�z� 8 Y�qʐ+^(C���B�=��B���߉O�$��J�p�]���Ⱎs���[~�1����X�M��OO�:R������K0�!�Z#�p�FI�+��|�7��7⵫\�邼+�����x�Dީ��-Oޥ�^OX6_�%�M��x��2)-�t�{��e����?�����Q�7^ֺ�-��I�|�y�n�h��^�3��,i���ᨩgU*?s�x�L�O:O��a��1UKuz[#z����; ��d%����b^=�h����I�_�tik���t�R��O�`�����¢��韻��(e��Yq7�C+/m#Q ���u�M�,�[�u�P�������Uy7d�(2�Amۧ��0 |B舌��w�p��i��'ӑ,R��]�Pu�u/�L<Xk��JGU9�I�X�X	���4%��Ɨ�+�r��ڬ����s��E�S��2�8r�w��oӞu��N�
�y���|�5u �8��e����uq�]���������O�����|�=z���X~��Z�'��T$w+v��q#��OO��Rk`����e�6-��(���U
�Y�AE6 r����)��s�B���9�;{��p�������Ձ�a� �h�I2c��vN�-N9��ޢ؎P$�0bN|�^{(�����F�7���o��W�TG��qz���L�ə�,�}�z��|�Җ_��WK�mӃ9-G�B�D��0�!�.�*" �j�3���H�@#n��=���z���2Ycs���YC��IһH�d�����߭Q{F˔0���v����g[)@B���Wz9���K�%J��͑%���^a��qT`��JB��1A9��Z����n�'�e0�|T��G���/E�	�a����3Y"D�'�q;RJK$��7����$9,��v~�rF9��h�
��|�����x�TNb����-e��*X<�8ܲ5�d���(ut��6�|�&q'2��%t���t�#2u��*��>4�q\�9r+tYa��Cyq�d�̩G0�WX��[���l4`;��u��12���"޲IzH��`z!���עk�G�����%�0���0�!�\�_h��2��T�Q��=�!0�ٛ��+�mqA�s���҆�)���� D�M�� ��i�+:Y7���W/��i���8v۫W��ɓ�����m}]���D�7�8�6��۰�M�a��u�n���?�ո/C�銶~�YwݠSO�g�V��9wm�BuC9�^<�.�G�T�ʊ'� L�*�V�7q,�!�#���_�:�&_�W�t���*�;q0�󍴤w���%�N�,��kh�X5�T��"$�8Kx������ΐ����Gk)l�4.���ʋ�*O�V' ��(Yd�2�gg��`T�l�)Z���Q�!��5�tZȽ~�T1��'m�_�����Y�%���SiY$ B߉A;:*l��}D69��&+~��qڜ@�����\�ts�A��|p�z�sz�Ƈ�jU	�:hk��ٓ����ڗ_�m�?ooޠ��g���/a��c#�4�җ#����GܑU���ŭ�' ���vR.R25T��G�Ʃ�G�m�,�,KZ��8�&a�@	���� NB��UI��W��6����ܤ;�	n�,o��A�و	���J���>J^#ǎ�����^�@y:�J��[�9�C��C��Jw���8,�%��Q��
?�	���;����˼�x"ҞwjCZ��Zg����P��1�q<$+�T��i��r��J\?j1�&I���T�*�G��bѨ�v�lǦ�����,#���Bo�q�cQ mP��.`���H����$J�>��.���&#ś���N�]����H}��:����LW�j�x�4kx{~���r���qv� ?�����dpʉl�M�c�v��L?%#��U��V���m��go���k*fk��G���
��,6e)��i�C��/���Y$��C�C�z��G��{�M?ĵ6��vT0���%-�� �HGY�����6�eh�ٱg���ƳV�X��2��f��TD�$����G���A�M2S�V](K�Yv-����6;}u̴=���K-ĳ��s�o����V-Lc�K�_=�hY�hw���d���lW�ϵ��ܬ�M�l�����d���r��K+9�-~�,s�c"뚬�.�| �hL�RH�᭕i��u=q�H��*�R(\�bЙ�WFbh��H�w��R��*�h|�]���RJ@�M>`q���=��-òd,Uc�<�Rb9亅��:��s�m��B[X<�ff'��������ޖp�޼�h[0�þي#<�8�Sg@�*�S�A�g��K ���Qp���_ن��֥�1dX��@fc��
��ե�<�������<�0����#&��bM�6_F߫��Q�/��N�s��+�H*���ey�;�E�Ʊ���G������C�]?HE����f���a�Ѕ��mm�|�*��4�2��j�B�0^�.���)��k�,��&��w�g�*��xG2UJړ�0�H�R8N�1�)��<�_�u��%ؠ4�8�Ўla3b�ҁ?�(�߉��,w�+\�����ԣ�����Fީ�}ߏj��Ճ�s�<�K^����E�q*�o�M=d$3<�� &ꬔZ!�������o����{(�7#�A���E#"�}�.]��n^����t�Qp��;9��#�O_��-Q���d��`��ˉ�-�6ڢ����.���|��O_�%�W�xw�s��X���_ '|}��n���i$~�91��U��a�>m
IߩsWƷbR�z�]I�G.
j�N.~w�}��d�E�^�pT/#7�i�	��O�<ŝ<�=����t����S���?�t۲:��2jW�A�pW�H#u��,�h�[C8R{����"x���v������Ӝ��G��:Y��K�D���˼���2<��zNdO�w��{��N]{%���?��^&鯼?�P�LH9��L�1�PW_�i��� ���>/�h��w���Y�'߫��c}"�m|��!F���@l��'�j���M���'�������m���ꥡ��)�I_���9�	_"��Ӵ�޸���V=v&3�B�\ң�b�i��	����J����BQǌx�tz��_:�ŝDX�P�K�}m-���?�KSG��J�L�C#/T ��#]�S��幜�,qLG�UF����?�TW� ��:��B�u�\��7�K-�w]�\�����K��t��zu�}ą�X�=�+ǁzr��e]��D���L�^��V����ԃ�Ʒ؞ST� /�ov�Nm��|:g�q��9mJZ+L�}�)MB6�Ԗ8Ih�h"�I�3��6_��h��g�fdr`5y���ԟW�i]�DWh�����)�d���ۦ�G�&��v���vnn�MO���:'k'k�=x�"�70�0�4�ͥw�D��o����(e�>�'���L+�JwLP�+R�h�ʿ��r$�H����q$P�CD"��!B�SDQƧ�a
A�EH�[h{�G\�ӭ�əB�ar�j����v���v��嶸���������ߖ������ب���9}/�� &��W:\މ N;c�g��L�G?�r ��t�jO��x�֩���Wu7M�PF)	��D"f�g"&��sa��K�Й&^L�3a�����wa(b�9w��.�doc1���Yu�}�����sZ�6�6��ev呱ij
k	���i=�N�,#�#EC�|��/i04D�]Ѐ�v�_�u�1rI���;aߗK}�qz	~�qQ����S@���o�9��p�����y���w�6N�A�	?�+�UPnU|B?�_�+{-���6�?P�H6'wۨ�
���&0�{�_��V��t�v���t���yW�~�QU���~�N���~��^9X ��+o��=o�׻W������l V�'m�|9��Ю_�֮]u�q�{@�.�����ы���R���r�cX��O��ʶ�g�-�M�"nDj[U�����ÙD�:[�our�.��W_�Y��V�ϻ����u!���.�?m�>�����;���w�����*��W啇��-#y�ϥ���o}�/��Iw<GV�L�BfwYH���ʷ�K9Pϼ�x���-;^ik�mc�#8W;�7���v�����W�	w����S�Ud�EW���~�q���uߞ�
�<��@^q�
fy r����}Wg�ϛ.}�Ζʓ�|���;��L���-}�.h�eotϑ%���t]��+��� gz�aj[�GO���z���f�L�\9ɍ���	�(>qx����~���Rl*n*G�)w�F'�ɿBp�Ѣ��] #b�N��x�Ӑ�.ܔ��m-e����*[ӣ����8
�%IF/
F D���2����������*�N: �K��-���*�(o?�>/�dT� @}g��J�0��j:��� l��W�B����~��/4a�<GO��c�v�W�.6OmV���1�rz]o��F��Ĉ��CtrpM����I�6t2Z�3廿�}`���]9�G����'��6��M~��ە�x�F�=�/v%߬���C�=��6Y�G}�?G��\�t��#l�%6��2;\��]2�Q��{�e &��G��n]mɓ�'j�>�z�����&��ՉP������RO�9�sr]�'��b��)������������?���~w�=G� RrNV�Bk'�r�>�)"��l�X<���*oV�-��a�"���I��T�+�;���� hH�7�Pm͟�h�P��b�:�J��s�,7����ps_}�J�y���{(���&W��t�ݮ�����ƍ��mn��8Fdk++{���f{��S�w�cn��V�u��(2~� �8ʀ�-~�B��Ν犹���)Rv�z9ZNG	���O	y�Gv�t|%�"B�`��ѱ!3���}�Gzl��7���x�'ܶ��k�]F�lS�� ��*������o�a��Mh"mL���~��� ��t4�4�eH[+��S'��t�:�ҍ�Ꝭԥ�<ҟt��8Fķ��A���C��m��G�|�J�mval��@a0[�rSt�;z:�n�Nn0Iw�;��`�V�Q	;�/�aϟ�6m���D� �#D�=�4@#��^S�l{�N'.Txĕm��LH/+���^���e�����C����8Z�:`Y��Gע;�M�Qb� ����Ѥ�j�(@�X��B��gw����V������pi�ePTXX����ڮ]���
N���ڳ��C��'�[Y�&�!�q��"G�/5�l��mű��KOjx����/��ҿ�:��)Z��N~wW��+��q���������������.�����:}��U�z>=���]�x4�z���U׾g���ܥ�٫w�J��,	|.���]�.M>v���%W�H�;3t�6��q�<r`+<�F->i�o�m_|�M���w��O_���u��F]��*ݬ��:y0����K8*�)l�I_|P��&���$$?����/���{�8z�ջ�2aW��)���x�Z���μ��(�V>�o=�6S£KK>'�~ۿ�,R�I��G�g�O\JRw�F��0~sD���]`�\��Rv��;�R��v$�-H�˹t�)� �瑹'�IMZG|�6�C�cur��)]�W��o�	:X:"�玶�EО�"��Bi#D��V燏�]�E��"�������r�d�\K�R�>�9iX�����1�:��|��,~��l&��wFX�z^�L}���	�R�k?�ۅ��X����"��j�i��G^#�Cؑ�J�_�"|�o�Y͆ɴ8p�=�S�Fi�\�8��ZRO+���B��Ց��q��S8V��ζ���������aum��c��QN�e[Nl+�m8��Z�!|q��"��^l��A������y����K�f½
(G�%8o�{�ލ��]��w�:�qS0�m�]!P�0�5��i�R�����{�z�&���y���k����^�i/2K}�}D�t�fە����m~�F��d����O�q��<[�)�'_H]�޳��j��+A���fǢQ$������<F�����C5Lo�����2�^�=-06��"s�`���B [u��r$wb����6��ɩ�6>9���>5=�fg����|���o��smr�mm=;Ag�M"�%�ܹ����ﶷn��.\��&�f��ӈ�q�v��7;mu���a6��g �9@�8����rG6(*Ϧq>���8q��?�]�+m����ޅlr��LIԈ�'��6��������n���s'�u:�Jd��TQ�.n��O)�d��swa�(8�~,;	��&op�ru�e��u�|�	���	���VA�T�,�B�m�n �a[��O�q����5;P�tb�:J��Y���r���3'>�EA0���ӑ3N-�Eh
k��t�T�(��/.e�r�,#�"p�H]��ɩ�6��}ҝ��׎�ɇ<�$u�ų�KAP��I�
w�V|���0�?�����ͨ(�]A���}�F�Yq��s�JX�7���"|,<�`C&A`��u4:P�O
�w3��� ��!-��߶��J��U�v��"��!_�s�,SL,�5�Bp�?ST�`��;���g�=�Ib��;l�ss��˄Km~v.�\_�k/^�i���O�.�0�E��"x���(	��P�	PG�a�Y�I�P�"���e�?��L��.u�����
�3i�H���ȳ��/~'Z�4ٟ�������������!pte�U���_��(
�V�dy����!9y��}�#�����w�O,uX( 2�7��&�Q�"��w���c^.ү���?����N��M���<n��=l�p��?_jo^�9��̕[�}=���^�%?���ӫ�����J���ь�����;B����V����e��\ͷ�H���������,�b��#���9�+����ްw���;j�A�_���Q�J����`�������]c�������!B��uԔs{�k]�pd�K��৪���㷢OY���d��0��=��,4h�g�QBm
��e6�Y3\���'ـ��Cm6iZX�.Q��D���Nxć��(u�Qp���sǎP�z|Ϩ3{��Z��aj��>�Q �م���'N`�Ʈ�S��������?�{u��I� ܨk��W�A��z��,���Ԧ�^�o���1��̹�
��`��`M�fj
�;֍r�_�7�s���:HD�I�6�e�w������� ��Ӯ�G��o����)���������2���u&��	�>N��n��~'d�k�8���D�w �x0�M�m2���n�q&&=pz;e?m�>��R�����u8�q`���=�SXB�!<q�N���L�s�嘹y��t�{�>/Z\&��#vl�p�=�4��%�Ha������x;��u��Nօv'kj?�F�������q�&�-�=_��,������F���d�JD��Gz�2-�ŋ,�M�9�(�	��$N����<�RJAI^J 	���������j�� 2��Sf��F��(�ff��9�N-.���N���m�in~�͟[h���:Sh��-�=�gxl
�E(��0��L[�x��s�v���63�������8���okk(�㶋�:8�)�	�c�d5Q������N��OM϶��9�IZ������b���}NZvt��8�:.�	B!���݃�L��������8]�Ӗ���3�ޔ���f(�CJ�Ɋ�D��A��Gl�=q]�!oG꺀(L�{��IK��n"B݆5�en�O$(޻B�f8�(�FC�Y�sd&�&wS/�8I]�CbcD���;�R��)mH���`�vq4O�%3�{�Ό�N��p+ǁ\`@�QC6CPЦ��:�<T9�>�s5�}zh�|�T0�Gz`Ҷ���r���NO�DH�!�8om"l�~�a	=���sv����l�l�#~R���*��BJ���m^��J�PF����ֆ/�GR�ِ^P1S� J�~�ptH�(�J���9�ӓ���]4��Y���H��+��i���S�V�X��烂2�Y��0�ӻ����u�M�;G���w�s���W����͛5��U\�(ʂ�:8|���W�޺Ĉc��D˷������S���_��c[;��D]�Y2v[>��������֖Q�	���]�|��z�?����-���s!���	-��7�u��O��W�ϻ�P����YGs�7+y��S�&}��r��њt�;?�F~V��"��ҳ�`�~������ S�9��N1����H���A6�}�;�Ca�o��W ���|�07��s�t��������������N���/�����Ս-���ޕ�pY���=��m$��i��3�.I�}��4�Ī��2�}��ʰ�^b�L�z��*v+�|����5����弐�2��$�p)��Q�4e6�Uv�k|{/�ɀ!L^nFq��k�,F?�L'�	ɧ�)���s�W���'v`-��C�d�x�@ָ~
̑9�8�L�����a�o�tAR����!it|t���x��޳1���}��R�:����E a�Mc���u�
҈a_G�F�C\{l��p5~đ�S���q�ϲ	t|ߩ�@�Nց��ɰ��Kg���v~贏iwi/�7w3Ύ�2 8�ѹ9l8�z�[�k��1� ~hP�xl:�#\S:-�v%�eX?G�t�БV��#7Ea�}�ٖ�#���:����=�N�H{���g� x0���t%l:f�G[�";�'�Mz���Y˙��ah|�y�M�*l�3أ�"|�?�!6�B��Yu�x���Yl}�*yU>��!�LF={��4S9�<�d�������-��W���ɱ����5�un�'��d��O׿�d��k�j�Z1�A�O�`�٣��hq���p��#!��R(�J�d=�<L��ƌ@P��F�'��թ����,Mc�� ���n򽌽�?�IF���L;~G�r�~�j�z�z�x�b;�B[<��[8�����/t���"�4L6>�����fg���9�^n��\�"Ԩ:�1�k?�����֖#=����\�\��Ն�]�t�����
�868Z���Ӕ�TB,G�H���5��g.��YZ8�����0O�W��M��#hNM��Ӧ�B�h39�<�t��}�s��4Gh�9��N�́s�ع�I�11?`�����.����>'��"�8NZN8�<�]�K���z*pu�,o��wʡ�ƺt�����Oş|:05t\�t�2�ceZ&ww��=���9p��HVũ�D~S��o�n�
�$eFA�@���WH� �'�a�8:��/@��.�E�:��8Q:��|�O��t�63G<�Q����8�(�,Nw�=��J�'�Ipk��q�-I�1�TٽN���N�aʬ��tDYg�'��FE2���|T,1<�e斆��Cd��3Z�y&�Y,��ƌ���{z��s���,�~�T%:�&��!�B�>��;�~0�q�4+kՕ�%B�6��]m������a[]�hKK�s�4��Z��yT�^��o�ו�����_��/��G�����ϔq���w�����ͤ$o�����������*p}�ݷ�����A����j{�G�Կ�:��F����������2�����s����5��ݑ<k]��5N�\���T�͈AC"�ķ�t�W0x�,��(��B���9$��r�W=��W�e��	<u���9��e]g����[�6M��c�&�`)'%�gI���[~{9�S6/R�	���v!�pB���<2��R�Iq�4�p��i�Cӻ8����h�lF�A�y�zi7	�i����iҙ/y҆17Up��7���alGwf$i��?�3��+w�Ʃ�|�8���%}�:�����':2:8\�*m-��� w/��\ƣױ%�&v1��1_m��~�w��IW���W��H��v�irL��cU�&��Rt�~&��Ym�����H�b������6�Mg�B�qrtb&p2l7�r*���2
B<�G}�O~�@�8��o'���x�p��a�L��i��3�S�l���2�E:AV�F)���2�e
\���!��sj�N!����l�$>p�J�������L�$�f<��v�l'��T#YP0��tb�w���g ��td���/t4E���q6���gI_�hZT�Tj�؞�4Z;��u�2.iͶ�C�K���oM!�^���~����8��t�-?�wNXd���{�;)켈�5?�.]<׮^֧�j��N�#Y;�&��R{�9Y��fH ��E��NH�2�0���E�|c+l"sX㓴
'�ʤ�ƲN���=iz���Ù]B����~��b��:̊����67V�h	.75�9��/\8߮^��n�\ݼy�]�~�]��*k�F��/.����T�I�:6G����( ;J�x�5^1���75��F���l��4��7;��ti7��T�f��X�5�a�A���:+::[Н�S���q��稏=��n���::I���Lc�]��<<iGD�_G��q�t�D��)�:K}�ɛδI��ټ\��G�k��,�� smv�\�����`%=�4�YG��8X8K�:?8�2�qu�FeB� �(it�t�t�gg�QN���R�� ^�̓���B<���9�(@pr�(jP8����йM�u�N����yʛ�����
���(幻fbZ�S's�43N=�l�#���2�Ϧӑҁ;��ӯ�EX�y�rsP5�ר�Oĥi�;�A�f1�����x*N �Qx�AF�'�:��#m�{k�˗�^�,�p�Q��^3���ִ9n:Kq,��9��V�N��H8�d@�a�ę
/W��Q5������R��N!CQ���4�R�
K�y
���4������Wd�7� �u�m���{�r�T�s��9h�)���t�6�+8Y/��۫W��I�.UZ�����ga��+X�΄�W��.�Uu���\���:y:S�Y����[��E��O�5��W�3��-�}G�5�y��O^���2��<�����ŋ���c~v������ ��L��M�6�G���E7I��e?��[���<,Z��>����Z��s�x�pU��di��O�d ��̻�%��3������^�,w��O�L����+-��q�K��
���?���:I���%��BU)�vF��eL��di�	O���g9�U�gZ쑠,�K4;��|���ܽ�>���w��+�md�=�� 1@ο+'��ձ�n������X_�.4�����A5�����h^	�K�
���%1���kMV9Yq&��F�:f"QcVz��F�#;�J%��p2m����q��+��5�k'`g<�r;F-C��ߖȔ7J�3@|�HۘƵSq
���N�l<�	�gd#�&�������5�����3t*���n��Pi����x�#i�gT�:�9g[�����ҩtdJ/�[8,����8�|j�(Ԏ�!pTJ�ߑ27��=��҂�Mk��'����#z�I�q�n}����x�#p��M�
:�>;��i��=�h��r�t����"a��WGة���J���	g� ���W#c�z���s
޸[�1hA�����*���c�x�l���,K��mt�ě�M�M�^�H,�9I��,��_KGPj�,ˑ��Pqt̼�_^i[���R�����.x�¹v%[���:Y?-'�s���l/_�����;G+�Z����d��5�V,���1W/Y��!2�]�ʈ�#�湳��8���)�+������$� ��08Xk�:��+d(�٩��/_�ɺڮ]������<�&^����TE�N;�8��u��%P��]CPG���@� 1b5��]X|{muu��Vp�����F���&�N�Ɏn����ye��9:S�1�{�݅�w9\q�t�X52�񎣠�ᠾ� ǘǮ��4�n�+�t,���6�9�����ұ?��M�{=�_��C�T��]9%��o���EȤ�8Y�Ε��L�&#�c�<�'
���:F�)���,�F�g:d��ϨO��rz�F�K��dbFx
��|�t�tVm��B�������o�(��e�a��
�n���5��cFY:F��
�6�R�K4܉?n1a�L�xNspz9X�O� �?�`��ř�����)�<R�9���f5�g�k���{�)]�Su�`e��3/�=B���	0��C�(3�Su�����h��=j��S�#Φ�1����,��c���Ĺ0:cʊ2U21 x�Q�;ڥQ� f�3�)C��5�ӌ�=��W>���@ ֹz����t:a.\��.�OC�m{g��^Yi/^.�e�,�����W8�YX@���$��5N���N�=y���m&��R�]��X׷�Q���ǃr�G�ay��B��V���	��Gߟ��s�b������� ��/���믆�۷ޝ^��l����h��V�.�s}I2�$���W]��:@C|�����aӎ�G��)߼L�����Li<A]�x!l3M��;����Eɱ�W��&W��r ��,�S� ~�{ϷI�%�Z� 0��Kַh�X�o>'p1�y&V�"�*���|�����Թ��/5�Xρ�#��)w$�fZ:Y~�{_�I�yC����e�5��K���3���$/��W�!�ȣֱ�.�§c@�;S������E��^�Hd�r�:r���cෳlGJN�&��>u�hT�h��q �~�B��z<�!!F��6Hl-G��D�VXm.G�zGA'I[ ���rYXsV���|�O���`��/;as(1N���8QF.��n��N�˒t5�c�:�QgN'�Fv<#�o�;����f׀�����Љ�:��gm�NڲG��r0z�����[�����w.������Y[[{Y�)�I-l�ܠ3e����)��gշ��)��)��Ӵ��A��	��5x���l [������Lp�f]c���N��n}���j��e�D阙Fg�N�����p���l���֤9���;�0��_�"t��[���;��ͭM�'���M|K�:X��y�/�f�*e,cǩ�З����V�M��m?9>�uX�.̷˗����ck�=��Z���0b;@r�,2�h㟽z���K�n S�[TO&�֡H �"+Ï����v���[ u�<J��01�9���,ojr��������yh$����N�ŋj*�B/�+�K���9c��1��8{�0�1F�>�m��e�P�Q����ﶷv!��&��]ls�t�A�C�nt��@ڬK�,�`�x������U�Ҙª�����tq�$��/%�;\~�G��0�3����N�7M�}��8�t��L+S��>�'�C�eg��nH��{a�iU���Y�q �'��	�.��M�G|����#�ԍޕ�1l:ʎ����DZ��	с('�~[#{3�7q/&��8A�Y
��ʠ�I��l���m*GI����Wkq�S��:4Ҷ�'�t����%��uY����1+��7����̳y(����M\;�΅ө���k�qLqfu4ŝ#���-g^Z�P6�b|�uT�0 u.�@�ԡ�q{����X!~5ȷ���Y)���!U���O
C��&B�����#��z��M�T"��{a 	y��ژ�!ς._�Cc=��P�1"X����=�5G����D�\���W��I�o���W���8Y�Ȃ�٪p�?a�N�Gx��zv��2����?��_uY�z�N��>�d������"��~�������?N.3������XI{p����\n}�u��v6�*���U���N���6��A@sb'jů�+A��>�EĞG��*�c9^]F4�t[y@v�0��g���/Q�FڞǢ�����y}�Ѱ�L�U(?�OzI}�F��?�����w�6���)����Gq����o�&b�gRԽ��#>N�A|�=��<w�E�ir���"�	֯�'���lxD�|E�L��ߏ�x�u�V�ӦA��DV�(�i�_�J�<�M�����'��'~zcR^6��׎n���HݕR�Ǔ�?�6v�%�#�רU�g�����˔Hℎ A�t�r,�O���lg�D�[G�%�v��l���M�c2n�Z�`b?�����9?�`�1�SP�m$҉S��ֳ�S]�y�;�[ ;2�]��Ѡ�8s�*�u04�]�-f��^�i[�#:\�<�d� boRVL~�S��3��\#:�B�����-�@���\�F�82\:=����08-N|Z��`�/N�|�]�E���Np��8:L�"����8{%pW�ĩ�>�n���i����>��ě��fN9�������ea�g��:Zw�e�k���;uvc3�,�UmAy�Í/�[�qř�Y뺍�S�V�y���Jl��K�����-N��޶�8���"�������K,����+�$�:���ebl�-�M���e�yG���V���-�����������������Ͷ�EV�N��0%r�,�;or~c�L��v���&����Y��I�V����vr齃!6*���!F�E�kkk.<��� �� ���Fn�8����wb(ö�0r�������	m����W��[o���z�F�Ο��x�0���;�� �	"���P{�B�o6ګ�[���N[��qrX_b#]�"D$���W]�r�b��+Xb��p�D,Y"�OG�V��䡄R1�'����%���\�7�RA����	'ϊ�b��<h�o��	z�6.�%f�G �ޔ�ۗW��c�TH�����u4T
�r�<�m+�w�	h�����]�h��F@��o�������-�3"}أ1
�;��t�;[a|�I|���m
{�2wH;��UJ)HI�0�� �-V�������p��T��]�Au8(pܙ������(�l�����o�QBT%�������@bv�1����e*�]y��w�΄ݝ����¥��a�Ys@��?x�Kԗ���)�_��ml��>������TVO�㝽Z���߱�T��v�ه����R��E��l������`t��U� +vv��8���nZ)6
�Z��� *ߤ52 �iOy�ɢ�ܺ�~�Ïڏ~�q{����8�=}�>�����_��}��ȍ�Ȯ�N�{�˶�y����u��9��;�������(9qN�뻿����r]��V��3�UNKQn�0W}�.�fj�I��W����'���$�?��zW��/_=k������������)0!��7�|��H�>E�W������s/_rK�£�~�v���i�>���1���i���%��T���t�'��̂uW�����e����ֻ:!N�����r���<N�<���w�z����4]:��W�b���^�(��H]���9�� �V��.z@==��p}� N�@ɦ�öEf��K����U��.`��^����NO*�sF�i f���s�,�v���o�xe�F�~�\ڲ��,\��9r9 d����r�4^��x���9
]�zZ��;�AG������t���v�V���ף:c	:��/` �ΓӳFF�����iW�q�i��[R��:Ru��EM@���ȋ6G��d�{�􎛼�~#(�Iꪾ��v�,H"3Rt,�p97����8��v-���;��"�[�ko�A���~�o��I��3G�m�
�h�_b_Qo���d��?Gu��?�h�#��;ڰ:��:Y�I�c?y�^BzQ����Z7Y�m������K:��2//�`6/Gvt�8���|3�H�X�� "
>��X��'�'���)u,m7F�oq�Cf|���#ެ�N��$&��i��,,hR��N=�c�8�Ni�DH���e�8s����ڃ�$��"��O��H�Nq܂N��N~![�r��>�|���l�������+���~���ݷ/������Wvq��q�~�e������{8Y[m�u��8#��
���t�F��{'k+���aͽ�������"�W�D�{±!���c��N�J�a�.����֎Χ��wp�<�cg{#�j�,�rKH����;q�t�\��n���Ef��9��W�Ǵ?�a{�1�ެl�`m�e��zu��m:K�TG��UU�Bˤ'�y��3�oa��8Y%�R2Os��B >9/��D5v^{_�`�F������Asr����|��I����T�H�/	R&�	SB� e`ۭ7z�d
�y�(�;�i��.��h�h=�q�¸��v�N��޻����`PП::��q�p�)=��TxQ
���&m�X򔎃N��}�I��3��Э�{��[�W��X�r���I�!�B�afi�:X�Lo ��*sp��ҸҼϲI�
H=�9�02�p����7��)���C�t�0�����";T>�[�" _\�JxU:��'��o�uI����9��2��}HQ,���W,𿇓e=�$-'��Eh��
v�^?=0�4�n����Sai���"�<�6U��'���t�~z�ɿ�o�tc ء% ��c��i��~��8X���λ�BOۻ����������i��r�Mzy �څT�RҖ��g}��suxP)u ��+�\E�ً���r�v���R�~��r+`���ʖ�[���s�M���og��5�_'����wu�޿.�.�30��[?���/]�D�땺�_W����9?��`\KNGh�ה���^��u�J|��4OZÿ���c�Mˀ'rƺ̷�B�Ǔv"B�U�rR�3W�^�ힺ�?L�����l�+�Y|�-���E�[0J�,�)���ϼҠ3R�(W�� {��"8�=8D�j_�8�ɦq@�Ț8(�+�Xl#�m~;VH���NeW�^�K�"����wn��ov `���k��xgtŶV�9�K���o�U�k�츣0p�ѯ��4I38�~�uKDJ�q Ե����>i�Iwzvs$��]t��ͽFGgѽ��q�� �z���	�_�S�G��:�B}gEu �F W�Ӯ�u��`u�Z:h;m�thp�n����4��k;ќ�&.��):lꦚ�_�둸���:
83jE~h#LQp.�X��DI�s�caY��.v���$2J}�~Aeő��u��� �C�=]�Z4��x//zI/:Mq�K�!�M�ҷ��mUv�q����O|/� I�r*~����!��K. �0�bW�p��:��~���?������lR��g��O�[W���t#�*x��.�ԑ��i���6���c���U4kR1XS�O|�e�2��"��r�Ӿ��Z#���]:hy��� �g~z���c����z��+��|�d�#Y��������,R��K� D��v�˹i��(V�p���[5�EL��1�jF:�1`jƔ1bt�`�+����Kd�dI02��j��E�-�nﶍ�M`�Ah@h��嚫�7n`��n�}�]��ZX8b0�a�0$U�9�I�@3;��[�d�ƹZ��z�F'k/#Y�q�hd��,"�KiejK�鈊�z�hm<�2M�6���t:�?��_!�3!�W�,<�����q��E�>�c�K�|.�5�)gyfkܔ��� 5)�Τ�ʨAPB��:��A�4��P^~?	�q���z�΋�<��pJ� �+�PF�k���թ����^U}l#q[�>���ZCH>0\�Ҩ�����N��6�H`C0�>�f���!�]=��e*@�3��x6��U���ૄf�����ҥq�Vx�:R�)n���2�^:_�BQ�m���N(�Xg�G��=����|T���m�d~�\��)�2��AY�R 3���&��N��I!Vgs�'>�?�.�����NX��_܀۠��l	LɎX o��c��u�?w�Ukmm�u���h���ضf(��ly�6y���Z�������?��ߴ����{}�nܘU,!�s��/�����'N֗QȖ�;YE��TT���(�hԒ���>�OE������:�O_5���]�\'����*�<z��5�/#F���{E��<�>������ī�/W�_ʨ7���,�Ig��]x2O��S�N 9�Yw
�+2$;�L���>��w'��"K�zJ7⦧52�{��^yWɨ��L:g �h�|W���������c��H>�\U��\�O��E��=��w��qY0'�3W����������}ܓ��+xȿ?��}���(�34�A����8z �=95Ҧ��TSΖn9�A=�Gwa�{�'"��8⎰�����n�9�k}}����D:�T2Ü�p$@(��D׳����nkm3�L�"���e�ĳC��l_�@eM:����ma�lm����ѯ�2*���7<�A� O�>����y5B������ �?�͌&��i�`���i'���:t7���M�ӄ�އ�:���MQ� ���:�:Y�������i��i�����1�����ͪ��x����X:?vV��o$���9��U^�_�:뙤g`�|$Й5M*b�|�*��c�ɻ�&���(����d�6nl��唳�ly���~��v�m�D,�x�Ë��8�Q�V�cg��b'*.�[I����1��8=����G�<F �څ�YٓW��Ӝ��(����iGi{;�Ň����6O��)�1�.�������⏴�C`�q�l���|�e}���&�q�s�So���8<�ɒ�h���vnf��wv$�+���p�.'�����j�Y�d�����E�5�j$K�%��ɉ6;5��a�]���uG�`���.H���VE�,��C^�#d��E*刂A�3�`�V�Ew�Zi�B֡�+a66���se/�B��\���~��L�t�r��s���0D$18�$�y�f�dml��k�&���s�����ES��%�{��!�E"<҃*���5B)XeŐ�v�BBq0���g�0C��==#f�u7a�}+�@�Q�����E`0�uH�;��%1�0���7���)�%yJ�����J�m�6�2���wE����5�D���
g~�8^�s�ƴfYeh�������߫�M�H�7a���-G�]w��� ;�Lk�fY˴�RJ_�TZ:Y�!2�c�R���1��������YN��-�dn�&�{`$U,�t��[	1�4�3�&�g��F|�Xt@m�G�
7�92I:*�[ȴ߃7���6k�� � .q.N�i#�5�8�N��S�㻽l
oG2k$KX?���v��!+��AF���W����Wq�<������6�S)q��8
w�H�]�-x?|������_�'������v��80�d�o���~������?k�}��ԓ�����u�hq�BۍRux�H�i�ψ�eu?��K���K|$�p�2����ۙ�s����^ف�L��o{8�.�VC'y-M��o��? ��}�G�M����~��_�����(ͥs|��o�r�}��nE���w�����?�
V�v�U�W��M֐��h_�"������;'��* ,�T>�3��� #�qq�J>\)���UWj���|L��g}�<���+zDx���l\�}6m_�����;����s_�,eq���8J�@���Ni�s��s���s<� �jV�S�6����㔲�	�ӌ�!��v:��l������勶���l��a�J����I78B�Ձ�c��T�_/�i/�-��W��_v
���y��\��C'n����V��L�E��"ln��m7`���qR7��1�	��C`ݩMzSv�d�%������M';��l�����z!nY>M����	+�˥L&��_Tc�;�H{�F�p����d!��d�`g��#2��RQg���H&[��Oh�:+�]���@�9S�k�v��cV2����{���
�������p�#�YnxEg��g�7�e �� x���;�ގ�9d�e�(K>	�l����_K�}�W%�Y��a�ݫB�����ʔ��}�;C�����Ȝ����|uz9ܵq�m��/�'i�*0���r�Rwx�2t�b�P~��f�n�*�N�m��N��&�����E\����������U����c�Ni��x�H�G�$!����Cg���I�ɺ�'G�u�F�é�8Y�H֏~�n���w�{�\m�q���h��g8Y������9Y8�d�@���r4�邳�18�^�5"������w�;�� ��?[���P$XIrt�M�F'(�3��7<�AiCQ��8X~r��D;��&��FS�Ϸ˗/# /�������Nu��I�@]��ߛGmy}�-�`--o��7��N���A�Ƹ�,�^��"��D�NUO�>۸q���t�-����5�֟����6��+���g/��?F�Y�w.�K\&�3��q&#I���-�����S>�*��;�Jf�>�W_�N����T�ˬ!��̷C�*1'#F
"i��n��4�MP*h���{mSe���QʳV���l�e=%.���3�el��Fxq�CԽ3O�O8�F�}\�^����VZ1�W���'K{X\%��Jk��k$�Z�@�rtW!V�OXvZ.x���P~%+D�C!�I����������Q�
Sh����FgH�A})G�Lg�IK�d�&Ȼ�De�;q	�i�/q�p���N��*����/�E�d	_z�'�K�@���/`��h�+oڶ#Z�#_{:\�'���!�(�L��A� 88Ba�M�ζ}��/��O�?��ݸy�-.N4wu��;�ﴟ��_������}��ϐS��])e�QAm]�(LA��"��[�u�w�R��������#�r�J�.��s���(���k|���t���OS��q��W���O[�����5͒�<���*3#�(]]պ! v9�743�p��▸���<�!Dhݥ�RgD��b������]ݍ����������ݏ�7��;q�_=��2���~3���Q_�WW�sq�]�Qu���2pO���wB����l���YP��~�󫺦��)��	7�!cq;�,�/���E�`�������o����eL�w�Q�7�������p½����2�Zi	#J�3��&}6܉߹��%'�񳶼<��޻��{�A{���q_����w|�|k��ze����xO2|�7�̐{O�>o�~���^Bۓ�㊗���]2{>3��b}�����=z��=��I[�
�v������א[W0�<����U����W�FQT�ƈq��z���'�vbpi 9޺J�����	�� �|We�����<��|��+߫�c�7���׀W�V��	�K RR�Q�j�-���<���M�kR�]���='U���Ġ�c���r��Um�m|LG�zt>&ǒ��E�Bf-��c�!O��Ex'�yI�K��I����\4b��U�*�j�<��ɢI���1�j~Y�q�L���IZ@��b�b]/�ъ�IP:��O�Ў�ѧ̜K��i|��<|NX~�E~������.����l����d|1�Ĵ�
 ��1�p����5�\�����_Wm+'VkK+Q � �O�P�F�yZ�}E����W�	d�K� o�o��F��Ը�9���H<ʓ�ʟ�I\�<����+Yn��w��/F����W��Y?�%F��^�ه��ȂK4�v����s/���X�=�����Iˤbede��������MmO���uu���)�5?;߮�\m7��hw�ʡ~��͞/P����2��4� _����^�<���=mkY�1����
��{YY�"����m�F*�0od/�G:��q������o�@������x�yh�2�������m�������_�^�y��ɧGL�v0fR�V���TLÓO��J�!;o-�����Q�߾Hڦ����Ψ
�l'���|p?i�� �W33�8��0B�i��5��p�t��_ջS��l�ȇvx/�}������]�G���*��-��O�T�`^���<�ĩ�4 ��6�_j��r?9���tO�a�������"@sQ2t˖Hh���Y��*P���t�j膠�Y&i����rIZuI\���c:!UO#vSo�2��@�A}�W�W}�.���e<��і����[X�G{mwo���x�^bd�z��v�721s���:AF��PT7v�<D́�m�Dj�ȓ|�������}���i��V����@�I����O?o����M����_�����%� ��V)����d�N�!K����]�Ԙ��pn<�[�o=˟���<��0���}q�)����<���L��eMUά.��UA����4D�����{�L3r��tU��wE�x��n/՝ڕ^>���6��=��%����Ҽ^�LHt��y�P�2��G��{9��x9�?ʟ�);�T��H�*�*K���!}�wb����el|�U�����te,�����(���K{�����e>��C�M��Axۗ������>|���[�O��������;��G.��M��ɬbmmm�+!�)�t�K�3W�rH��2N����	�mc�1�o!����3g�3"sl=�#������'km�٫��s ����L�%_�˚|�$|#_D�;9��R�[/��dgok71������ϡC��ܼ'	��\��<0ƈ�.$���t��%W����O�����������W/S��d F��t;d�����Jh�C(�����9��$b�V'��UTcL�8&�~�S/:���z&���@޾�%+�!ŭxƷ<�gW��WJ�	�85�M�g(#r��sx"[SPȚ�q��<ˣNRq�2�Y�\��mbd�F�H�L?m����N��u"��Z�վl(x�\~"+~�Z�bS��WҪ�7h�_}���k&�4�B��W�q�����7���5�������'�y��ƥ?Y�/�I,g���F����c�4p�z�:����4��u�I�gW|	�W�I|-%x �Mhf-�Rm��C�P%���f����� �4��-�]Е�;YɊ��ޝ��/�N�=�h�忕��J�+9;f�Uﲠ*�&ۂ�{݋Le�}��v0Y�YT��t�#�\�uP�H�c`QI���QqU�ܮ#��qu�j�vu)3G��tr��=��s��km���v��ͬb�]��t${B!����T�Y�����/e�}�v����;i�[�ڳ���ًm�������w�v����	&�@��D�Q7Kl蒙8�g�=�ap�����X�G�J��a�T�I�}�!��e�49�L<\�5�q�G��tD�'�ߐ^��+�"C�W�_��WUx�g�g|��%�����UI-��"�åN%t��4��$�#��*�@�̐�#��6�ǆ����"�.�s:
EtH;�u�MYtr�d�#�Z��TFVfv𹠁�x����|�x����T�c��_5�Y}	�Ĭ��NW�jP��b}bѧ��ԥ�u���s�bh﬑4I��+�%�hϡ�Y�8Jx�.�O�5�����)!Fz�b|��?�]�+ڍ��g�&�9�v�ӂQA�ns���5u���E���Wk�۫�(-�2�񵿿#�-���Cg?��U�z�5ѽ��9K����{�?��?j�G?l�A�}�Z;:8�b�٧�����m�W�~���@O���ț�<2��%�X/˰M�X�4�7^N�A�/q�tpv| �����ѳ�Eɯ{p�wQ��T���1��]鬻Wڳy�W����|*�t����ﻜ���^�3?�+��C�q��}C�M߈�;������5�+%��,��Ļ)�|T��91T���|�t�(C�a�"U��+^�4�e��K.���0�K�s���e��^^%T2�m���
�"��G�7�֪�W�7�B��������Wշ��i��t�/��V�$J"��˙�g��m��_������?o޾���G4�Q'��&��A[�J�'tS��,�0���t��;��nW�
rќ9!���	�r�mc��!O���1�N}�B�z���gyW�h���4=�A6�a�!�kմ�Ólt�t�����⣱55]u�.�]���a�wv���Y�9�#������?��k?��_���M't��e�^@#tB�;��'����0�Ȥ%u�Y0�bʬ�Y����ģ}ڎ1\�����sd�1���c�u��<�B����mg�i{̑F�-�E��D��1F+Y��
� �5���}U�5�5Vcl@�q�iȝ�k�8:)����Ǿf�$X�Rz|mu�P��
>蹎+�?'ҁ_�*m;�wëҁ�8�[�>A��j����i.��s��<{_sa����m���� Y�!���ꤣqjh2��.$ue҉W��I�,��9V�G�R�k1���IO�j;Ki]��R��-~v^��:�����v���{��q.�K����/��?��N9�g��[��#2�|�
/����w�j%+F�����<��������/�v��'/�W��ahl��*i�Ӑ��0Y@b�R�8	���o��C�{P7�	qU����Yџ9)d|�ʏ�����q?��S��wn���[�{���}��;�[��>�ֻ��w�g���w�;wn��ׯ���n/PeLa�����QBI�4��+�!�u�z�����x����=%�zg5�+u�6C�ӽ�4�����!� �PA�*�;)}�:�R����MX)��Cx��W���0����ØF�/_X&��K��ƫ߃-�G� �����Q%K�r��Pa�g!_������t��O��G3�yU�����k�'�8U�*_?�^��K'��;�*�Q�Mk����~�u�ί \aSP�ֱ!G��o�|D�%F��e�[ ̈��M[s��&nܥEh?�'��*�V>	�Mv�E�:n](�Ⱥ)�|J0)8�牓YR]�\m=9&y%�x�S�:�9@��\�J�@�W`��6�3D��̇U0�Eޅ@��c�5��a���ll�y!�0'h�ҿ߿�[G���TNܾs��j�q�z[YZ� �`���z{������㶾��2 �T[yeV�cX�Y8a�Ryr��G�QJI�|�����$�����m��<�x��@�O���>V^�Nɗ�K��3N��x�/!	�_Ҙ_�S����?�D�?8F��@\_{��a(�/�����Q�����M�_��G�Pϩ?��_yg�z(���r�2y�'��y���.uHxh�m�<��q�'��x����D9#^�}��Y�w�_��͐�(<y����a�^���ĭߘ��Fq��O�$��DL俔E6��֭���w>l������-O�#�Ep!��+G�LN���.��u�ᬻ2M�m~��(�*�u�v��L=�&e�V��e�!߸�#��ojYvy�v��(]ď�����x E�� �4㔒i;�r���l̻�N����t:'�<\*���v
�k=g�.�;[3�_�c�5:=�	<ɩѰ���M�³����
��^�j-��1�`,�wcmww$�c4��.W4�\yY�:JC�\'��F�8�vI�]'��Fo�m��R|�������U;߻�qEN�;\�� ����b�\-y�5u
9(��w�݂�F�9ilL��r�q�rL㊘bx������w����N9`���r$�4�rʤeQ7��ԍ�u�s��w�m?���Ic}lGZzH�����n}�.�C�7m݊/ms�F�����¤�8��pX�|��8և2|�p�:���j�ir�>yI�zo[���4�ݙfۺ�b�UW����u�Q/�~���O9�/��S����V�kEY=*:4�r�Lg<�DO�'OV�!:�J	Tu<i����kK���;Yׯ-�w�`�Y�;����<F�^�,�H�'V�����A��bd�����*������!,g۝�UxH0�$`�����;k�WW�?l��~��oc�o�jo�u�ݺ��nbX]��Hz=�'r��f��1,/%H�9f�P�h�(r���ֶ1����.�L��PA�VA�Q8�`�4��|2���qEٖI9u/FM�){�G]7@���Z����3H̢�x�>�{y�Q�0�)�擠�]<�4���/eT�p����{'��-O���7�R�)I���\v��E����xh�{u ��Uq.⍞�/�!]� ��V|�:��Z	��Vz�j���GA��i�ǐw�?FV�5,��x�"l	��Sr��a��eX��2��)��%+G�uN�B�q��S�J{~Z��@�Ocbdh�W�y���3�
@cgH#���G����������)#aeP�R�G��4qu��5�����B��v�uw��	����NV��Cl�SG��r�.����|>��ʗ��3���nR�`��
��V�s�v�ze�h^���ٓ�1��^�#^������e+��{�A��;��/�=Wn���-��rN����} #�#w�%r�g������� x��K y�M��H��*M�SqM#tŸ+ǉ�!� W��F���E����ט�ϖ]Ͽ����~%ɐ��i�J�CP��&\�F�^�N�T=q�W݄y'Q�׻�|y�sO'�p7,���'ωT8X^��iY�1�Wȏ��E�4sx�
1�*G�<e�=����2R����	Ý���e����ʏ�'%*��4���z�W�A�	��ſ�j8��5�WWW��o�oo�{?�)�y"_&��~����̓���V{�t��x����ll����w����g�t&��Fv�����\[��?�!\kk;�9�_��cg])M ��cgg�|�{�^���W�ڦ��ٍ,+9�e�rW�a�!�	�Th��X)Gwv�I�A���C^��E��n^9<:�<��TY����J�OT�X��%jm�4x�-����z��^�$�yxV�:"��Aޮ<� GIVao��ʘR�s�w\P�D�D)�1��2��-���>K���}�?��2O�/��iʆ�k/�Q�˹�C�0�� XY^�k\�4~4V4Ǝ=�4(��o��9��y��v��0�@����t� �[��Q��1��Ӟ�8���z����R��c&�֝_WV�c�O7��K�p�s'�)�����[��>t��S��U�Q�d&F��j`yҸ�jd?�@�NY��{)ǌ=Heiy�͓Σ��)am���Hd�I>�Nɳc����^� ڐ�F���Gy����1=�_^X��Ww�D�0ˊ��!\���5����b�N�������#{C�,�������έ�v��*�b	=�]|�mV�v����ۗ����/7�|(���ƃ$�d����;Y�q�Q�Z6T�@$9��K�Uf[Y^�����a�{wo�?���ۏ��X��g����a���9�0pF�.3TT�:{0aZ��$N;�q׀Ou�C!j]���ZV�4�d1���!�w��\�'/�[q��)O�[g;��[CTG�G� �c�S����5��4�?�[|-'� �w��cz�p'�[���w�/e� @��C@���L4v�ÿ�O)U>8���9��OA�mD@�sDL>����+ƏqC�x�jL# y��(Ӫ��2d*�ʭ:�~��^�*V�)�� ���v����g^��t�U�{��V
��۸���Àl��U�dCe�V�e\�������KnP��M&U��#ys7�ܝ����؍�ػ���XlWfu׀\���0�R����[["���G~W��Ú�(c���=�>E+��3*?��|A9�9�Y���hh�W1��T)x�v��8�&ʁ�*BٙC�P��B#k������嬧��`�En��-b�������v���(W�'�P`^<ў<~���Pc�R�}�Y5�͔[�;_֝,Ӓ���]l�ۗ�^Mϕa�{�<WX��{¸���=��6�����E��Jݽ�W�
�mC�9J7*�4�?� 
��q�,�2�[U���<��� ������M��;A�x��R�����8���d��5���1<��.��m�
�՝�o��/m�_������FhH��ͤ�p�r;�9�
Y�?q*�?�X��i#��!�j
��޾<��r� 9ee��;��A�[��G�k<�މgy)S�!N���R�6�Ĩ�j�=��Qi�$l�:�8~�f����7r��2�����X��`���9jO1�>��Q��/>k�}�u{�����������z�ϭo�hk�^�g�^���z�>����'�}�����ڗ_>���=z�<�fkSCk����_���Ϟ�'O������ٳ���^��͍Md�ʭ�7#�5����^W=�S��앁����Ã������2����^alitml���W�\�iܒ��Q ff]ٺM�[ՙ�s��c��׏�K�����h!r]���f��M]��"d8��6��_����W�4�����U7Oi����%��� �%y�/�x���?�vn�s�)�/lv�Uy7i��	�9ܫC�RW�����plr�Q��S%o��k��Htߜg�7f5��3?��ު�o��=\�:i�Ջ�����K��!�i,[��0�GF�_����d�~}D9��L�Y�2�܂��I\��]�>�r�6u|���B߷�r�$z�Ɩ�R��Ls��d���e��V#˴���;~J����;�:��H�y��P�_�����X.]��Nℶ��-�'Q��9��pW�����.��Hy�t�Ke�}Ŷ��%��@}�2��C+�Ϲ����*���F�;�dad}�x��E{�����0�FV���Y�Y�ϋ�:�Q��	�v�|[`��q���uP�.O�����$�X�[��l���n������߽�F�֔����4G����B`=Ɍ���
�G�.��]M:� �8:;�i2�>*Rc��]�+'�9<Byڛ@x"<������3�
O�U���h������\섴+"��|�P8�[���!D�F�s�g(i�n�KƦ%��������@�m��n懟��I��:��)��8� �RV��2�7�G�o��s�Mɯ=�����zr�퐞܋~p�
��*��ա��l��~�yY��2�3��b�_�����A2����M_t�'~����i:�����0��8h�ҁ�@|ɜ2��v&E���C���^�vk������;�T��j�p��q��o������xN��*�a(_!�wB�҆`�\]i��Y��Z�<C� �	������e(i�YF�ǵ7nH��gW��<k�1��]�2[OA-n�(�[�m{s�B�߁�8�[�<�\��p�M����%W��#�SI/1�j@��m����-28n7Vo�w���y�~�qc%�:]q�7��W������mo;�mꄉ���~4j��*u��C��+��G{���	q�?(�m '��#%�T0,԰�w��0�Df��KG0��q���t�%oq�t�^@��Y\�ɟ�oz�q� �{X�TDŉ8��2�*�2��o�$Rӊ[�ax��e��a@?�+�8�����x�X�� {q���쯾�} 	�䥟���7��(����[���r�x��땺�ֻ�j�z&�$�� �����&����ÓvH�	��<[�	��ݽ-K��]�w�Է�\P�(_Ȟ0����L�p/^*<;��
��o�В�Q6q�'������ ?U�֚<3�<�6ܸ҆�[���y��y;�:yZ۱�s\��;�n��&ڭ�7�[<UP%
=�����Ρ.�a�_�������_���������@O^<m�~�E{��	�ǋ���ω��}�ۧ���}�����o���y��ן������ˇ�ۓ�/0�0|��1��Dz��F�����_���Fq^�od�� e53�����Q��m���v�.ak{#����g���%�"�^>k�k�1�^��Wo[�o������Ӷ�j�mo�@C/W[.g����Xo�x�/��\�#�5&��Epal�I.]�F��n����#ߙ���g}o��;5.#�F��Of_p���!��8Ȗ/�荦Q�ʇ~`���xy�H�A�b-o�9��qbrj6cEm�7�f<�q��g�5�y߇r�f�be��c:[!=��������;k�:F���=u0���"�y��d�M_ ��ʻ4�d!��A���"3E9���K�"�8i�GOH�������ƾY�kh��i���.��9��D���`�NM��h�juzzc�'e���L�,�D�pU㏱�~�~m��]$�g9~��#���M0�u��E㹍�S2�YYŢw�7��U�T����x�LVM��y�':��OŜ�<�G�]/w�V鬾����A`��e��F-��0i�_c���&��ą�f5���^�]p��S����z�լ��(0|� ��2S3C�Q�˚�R�L�AB�2�� �0g�@J�zqB�VhŚ����O�z����b{�wۏ�����E�Y%�_q.P���2Au%k�C�Ջ~���.�E�l�PW�e\�!~�!#U�����y����������?ka�~�n�"�ÅqSg<��w ��P���.�]���']�XאW��p^�,;�J&#�=��U��m���:���k�=~U���߈��7������<�s��(i�k��VC-�~�J܆���W��zy����x*&��!J]<�?�rY�W+�(w��a����4����p���#�;�\Ϻ`�[eq�����
�V����ҿ�t��le�_�B(ˌ�mT����#�_7���{ō���s�ʙnzt�?��й��{'t����p'z����,��ve%q�#�q�x���wv�/�oݼ���{�<h75�fQ�^���i��8�#�*�dhC�L<�>�L���>�q�.��^ 'F�`P�r�N<ʡ9���f�d ̶n��m^�����7�4�n�X���q{xǳ�S�/��G�
S��N钏�1^p�����ݯᕰ���\�)<�{�������W��� e�0�wAϫ��3��;�/��,��_�k��'�rz`����|��q��ɟz���'�������c�r���P�2�܊�t�mT������/'���Ey���K;���ɷ�b���O�3�U�{H��w��d�}�	��4��n�.���e���z�/��0�q�����K㨨)�I��*���󽶰4��y�A���[�(~w*}�ͪ��W헿�U����I��O�>��a[��A�66���/���u�jO�b� ϟ�
���v����@����L*�"�+�\ǐz���=��y�V�<����۵ʴ��+�v�'F��`�a�=�]k/��	�1����m0��Cd+B���vѹ^���g/���O�w=z��ƻ�zi�C��ho�������ÇϠ����!Q���r,mj���*�U�5z1|T�1J4Z��euVX����
��!w=�)?�����ۃ�O<+�p��<Tȳ�C�9V��k��?0Xܕ ~⤲�������5WK@NB���a�sJ�c�u��X��c��{��;{���1J�	�m��C���Խ5�\��s��t�}M��t�.�'���1>��	@�ں������p+�+j⢿�R�]⧟��F�!<!���7�̓z��:~E7hM��Z$^83��F�}�6Հ�6�l��,d�֒�ݥ�ON���T��4\���~�_�;��lW䬏C���ǻ�'�Vh'^�e:�Ґ-�`��'�c�eD^�PLf���+YV�.��57��~�Ȣ�w#+BV��c��4��PX�,�)B0�xPxb�F��M��]u�'��Rܻ�����������Ƈ&T4���E�������]� �xUP`���v�o'��e��`��?�r�U���Ӷ�O���YnA:�C��y��g�_`'W�*��Y��Ζb޺A�V�p�������0P�7?��3�c�q�������e�{�q\z>E��a�|]������� >��oo�%�Pf�����,y�����~���%W2��_�7���C�^˪��c�/�ƞ�0)�W�u~C�߄�~T����U�� �Ѣp�/Hw�e���'?;Jy��+���-}8w�
:�nK����G�U\rRV�xuw�Hz&n���l��@;�O�֭%Nf�P��	B"�H�6�ƛ��3���n���;�!
�̔QO��e{�3V\�]�,�o��^[�������<~T�(5�&#
!*���}��;G3�����2K�(����^�E�3w�VuA?�/局��7@�'>�4w�E9�_��Ʊ\��&2�*�v�o�n�^
u7	{3��sl����	�?
���S�~Q�]5�_�3| �(�H�^�7@��%8����įǫ�V��_�c3��{/����ߟ{Z��5�</𫴖��z=Ӯ$�tI8c5~�'�DNH+�Qp׎�e��H�B�灦�ᬽ��0lh;��Jq�Y�,'�Z�8���o�W�%�钦ʬršʼL���ʸ�K��w�cy��mB>1,�2Ї����o�]v;���m͊�~\��9�)�ݼq�}�����nݼ�|�Gy�;�ʄO?�������Oۧ�~��^퐟z
2Ɗ��'o�N���~{���6^iTyJ�
�J�I��:<tU����࿋��m�� 2��&Ot#'��6%�y
l�xn)���0��0�4�և큺7���<O>�n��b[{���n��K�:�%�u��t]Y�4�+9 ���hd��`�m�/�zھ~��: ��UK���
�@��3�vX����a�ȡ�w�p����I��~*��t�f[F�;.��vA�!�'N�*ݮ�LQ�<�N��2��u�_>�AnYSQ�ϔ�_���KV[�C5���0��r����y�u7�1�mz-u��WL9e��h�a�c�u��r a�,����p%��oV��S'��.'��k�:�]�8�1����C��I�	�,��ԇ4�"�,xi�DNpI3�d��IC���(@��[��mz8��_Z���P��-~��2OY߬rI7�1Lz�&��`��Q�Y����[��EF5��8-U�� ��QV����w���kW���4�b�N#K��Ε��"V�è.��Ȃ�6���T�8D����e�_>�{YƩ����kO�q�re����{���N������tTm;��=L�������_�Ͽ�����eQg��" |q�.�GŻ���Q�7�~*��e�4&���Sg%k0�|'+F��FV�@>1^dT��[���g������"`��kC�YH���08�������i.�Q��m��Ǖ�����+��p%��w���܉ťc�0\<�C�~>�{՝��+L���P�>��wv��Ex�{x�']ś�`A�a������o��8���	~�ȕ:�\����ׄ[��őQ%�ܑ<�'���j��{�T�(.�
O�Y�
/�N�@�w�o�5�ъT��|�/��9���3(�V Zg�=��=ۡ�81�)���rDAkt�����B����+T�6�z����}�=�˃;�S}s�z�w�n�{�v�z�
CM�lm����/>�?y���*�Q4�a���X�7aP�����pH��� Π��2�(���g�Ҩ�B9(��∃�.�������y�������86z�,�K~�\�_?�E�&�!ݨܡ�Q���ᩛa�`(��%] >� ��Pw�P�N�*�ұhyq7O�6~ѷB7.
��É��������i��_iG�Է�-Џ��Ƈ�����W�Ye�\����
~����!5���hjˑOI��:���dU^�w���U@��<��{�I�P�n�<��b[�_�f�m"���e��<z>�7��`d�s�e�㩃i���E�j�*�"�*���}�N\�?�B��>ϳ�<�C/���o��}�c��Q����Q�;���``��O�o~�yV��Bxyڏ�N#;&��B5����^F����������n��xn����Csu�w�]��*�,d�S��  }�6��H�=�Vc�լ��Wygk{g;+]~˕5���=�X��ܵ��OFt#o?�瑇�����U��kW�#�U��Y_=|���c8"Y��2���z:Ѯw��w]�B|1A�U,��hx
��-���!-IA��{C��Z����my�~p�r\qq�)��$�7�-�Yī�~p�=\�/�V抏�K[W�40<�]y���o����(�wls{�+Y"�QF��%^)P���w�,�G��GM�bB�p�qa}�C��] n���i4� ����3q�
�|d��&�6yĐ�,��?i`�5�{QÇ��.1`�o��j9��V�\���د�mW�n�3~V���5�(M�K~,�1^#�:�s.��L#�6�*��i^V�1�B&}l+�P;-�	_��+Yn�s�Z�ze!�}�#���:U �H����ٺ�5�|NI�ό��� ��UR�CX�Ȣ��\/8B���˷�{J�[���}�-��М,s��gL�<y�>�����������j_~�={6��`|��of6I �.I�u��(���!���튌J9edM�]�,��U��<*V��<Y֊�C9�f���l���	�7t��ϝ�I���d�5�Ѝ��~)9~>����i�M<�zY������W�	�+&L������rW�8����7����"��+gw{�v,$�ѿ���[��ׁ��Ɋ�w=�!H^Ic{z�=@�7��> �7m�����n��{p���#���ɃW�
v��w����߅qGn0���1�ː�LK�Qe%�(��T��q^Ja�[�������C��_|*�X���
uߑȬ�
��I�ap�'�2g9�-d{�q|w�`�Y`����jd��������3�W�,�[�o7�
n���͏?m�~�E���/�IYGp� �2�A��y7@�&xf�Ϫ�u@Q�hȠ�2XAd�B�FAT%�Jn,(}��G�cǔS
/����x�����q�6◟Je.H�QX�JBV���8��Z���U��)o(;�*_�J�F�CX�Yˢ�=?�#�p��A�u(EY%�L���@��E�ɣ�'��nƏq�<.�U����-�H�!��+~#@hu��r`ަM����T�����*�^|%�<@z��#_V�eԐ��	3��Kꐲ��h���6�-��<E��K!�5��7+�i߁W�r8�Ⱥ�;�-_��]A�ū?��/�pk8Y�E��[����x�_�q�FZ��]�tT�T��(e�/�߾y�}�ч�?�^���![0�!uw����O��ۿm���g�%k(çmfvd�,�R%�3�����
�m%�*��*���s�#\-�Y~��G���RWkiU �l�4��y���۾��!�42�p#?կ4�\�:al��)g�c�/Ç���Sg��uYX\��\�!+�A��!�d��y�߭��ny�qa_�#���
�J���+���^��mg�*� ������E�y �D��nd�(��k"���mz�I_|�ĸ.�b]q��B�K���O˸zC�|���|�9�i����g��S��~��.�e���V]�ϲL㮱'�q���A0~�s�5]�K�֮捶Ʃw]\��A;ܦ��Y)��YX��o9����(S��F��|�ye���\}Lz�,��9�t�-��?�[��v���á����)<3�3а��r4̲:���Up4��G�?Wm}�V�NҞ^)����Z>���,�������oyN_:!O��O2��-ٛq�==q���TBCɗ+=e����PD �"�����E��G5�q�ۃ��ڃ��촳6T>�G~�j�}����g?�e���)֯1��α�.m���ʾg��+1�ff���r:���B�"2hp;x���z����0�0�v}ޓwN۞K�'�d9# D|`z�n=i,�))�l���6I��0�q�oCat���v'k�_��.7���&�4����&	��Ly$l�cZ�
�q�sq���~�<~
W�kx.����Υ_)��U?܀����N� �d\�<*�� ��-�o𫛼0�
��k��9��b�s,`��G����̊~���n�xW��x"���$M�����CY�l����E����W�ɆX>�8:p���q����3�_��j���9~�+rGc��,�4!�|��Y*�#s�	u�^�_t7�39q��򿳁n=1�����Ӊ�Y�o�l����J֍�"��V��o>m?���2����v�:?<g�/���=
�����N
v�V
M�K�Xo�U�R�c���`B�˙\pH�K���T&u���l�wӊ�F�yY,�?����qp�K>q�3�@W`G8�O)�*#<�?���!�a*�t�@X��C���T��I�O��p�B����˲̻�bl�t	�%�T*EE� R�tSO�φ�Yz��P�A��k��|(�r_��07^����5wT� -��`��#��k4�;��JQ=~�3��/���^>�<��XA�DW��v	N���E��]�(a��|�E�WҐOڝK^ ��{��o�%�����w������Q��3~R�O0��a�:���G��J�����o}о��o�w߽Ѱ�"��y���~��_������W_>Ɏ����D��o��{p.)�n_���q����.��t����Q�Oe'�aVӕ�Cr5@�?#%3c�+y�]�L9��r5rܱd�Z1Y�_,9�P�dRn���l���)Ʀ�%�����T��R�FX�T�K�G�M=�>�C!F���J�RF��o��|j����ab�
e4��0�DI�>�5(��b*�i�h�3e�ꓭ����.�i�T��W!/C�~��`@�c�P��BD��Șa��+}��S!���ķ<��	"�������7�D��`��j�ᶉ��A?R78�zd�g(G��)b�;wSe<��4����<��. �<R2xR�:ɸ�ƴ����ʗ��R�j�����W��4�w]1�R����{�W��J�;�y�H���73�Qg��Uh�B����]0�b`ݺy��,ϵ٩3h��O������D/�WB@��1i��Q�XC���s)nw{�my���N��T�q���@`�h�Z�n�}������}������?�i�����j��}@�ö���m��t��勡�f9�a���ȗ��j��y6��d'���
.`���'#��z�=b4���gv�ߢ�`\���B3'��+ �_��!�x>���ciF��ag<����8���ÿ�_� ��?�_�/�{*����4��µ������ mHO|�}���bL���������i��:��.�@���nٯ�@���"��߼���CM�����Kj$�o�_���`*И)�w��|:�C�����6a5�E8�n�g� ��qR��סfX����)[����c'W�ұp*AY3r�IX����<5щ��L)���2���	&���V{��)�ã������Eɟj��2��/�W��A����V0�!��^������ώ^��<I�g�"W��Q��K�瑿nú���y��cy&�P���@�$��
�����E��_���g�P��l+�����RO�X!O�j��S*G����4`����[���(���m���ӛWI�� �7�B˶�b��A��_�����m�1vB�p'q�c�)w�*�O9;��;`��Hu(0��eK���-��?zp�XG<�+^��y��!�
҉m7������v#$�l��*s�#�JW�b�Oެg���V�8��{_�e�8��3iN�QJ=�9U�_N�b�xr`d)��I��(�,�[��������mw�@�Q࡭x׬����{�i� ������B�ʊ��A|���0>�\:S6)��gG<��Qj�[ .nR�[�u��枣�a�	y����E��������=������}�>�*k�0p� ˱��e�c�;�fف�!eNl)����U+ܾ�S�'���~��rRI��LyD<��4�V@V�i;����򳽤w���-�z�>n_3��b��QV)e�i�A�k���H*�U~�f�:��g�K\�e�m�EM�`t�o���y�L�o�kHfB�62]݃_��ɸ2V�刟�%�����ʘ+dY��iX����4�����mF��m����iqL��h|�"�����9)�8	i+�$�}۶2Mm���q��7��6��¶�q(]�3�{=gLI]�@��da�w������
T��0i����`���#�ȯ�Kq���wU.��Yϰ_UpP(��A�����x�w��n�[,�Y���{;��)�ӯ~������c���ݾ~�4��x\t-i�>	��y�݆�Q2C�F��A
�k�����0����Hdp���\}#G��@Q"���tw n5v~�uóa����|�=�S�r�uO8=����@�����C���=y��(���,+����:�J���Ɵ�ŏ[������~c��+���p�#~ԯ?C���!q�6l�����#� ����_���,���h�:i�D!��U���';�eɣ�V��hb�G�o��p�C/�S���T�QH^8����xϝ��F�v �I�a��a�f�����W�g:*���D�H^*$�6C�TF�[�K᪼�*���(��I��vP8˻\~fo���Tx�U4'��wU�mБ;�=#��r�O��EV	N�u�mׅ�̬w��� �<����Peih���)o)�|W�2@�v��(�#�{�C��o��`�8�k۷+�~���@ߛ����tG�#M�)��G>�f��2x�|h�N?�3��I�#�R��wx��j��^XAȁ9�!�������s�CT�R܀𷼯�2 �>�{��������wC���ʫ�g�٧]?��ת\�~�o���	��t7�x��Fd1��w�ű�E��6��!?�W�H=č2�.ı�ܺWw�xHÿ���M�W�$u�H����x =��P�N��YC�{�t���i]u1�ф�p��>(|V�ڙџq�&*���=^\cj7����Ϥ���~�U��}�����r(�ȓ�rj۠@��%�`��FV�m�����㝏�N!���.�.�\y緔��jkWFU¤�z���_����(�$��6�Ru�Ih@\g��H�F�J�h%I�J�j�?�)n�Rxx�ޞn��0�|�k{3�ª�+3�E�`��G:��Jo//�/����]Y��Y����Fc�g�O�_e�-c�о*������v"�+=� �c�X��O�˪�f%��J�+��I��r��
��<k]��u�t�����o=,�r����oVץ�-��	��#�+�랺�e��x�Ox��M1�e��s$�3j���X��}�2���zeR�8j��Dg��t^�g������(��>ۅ��xNyC��D�N(#+�Q���i��d�bp	>��|*b�)��ʒ~�i��'���J_����������<�W����8���^b�*I�^�ђ*��� ��А6�BR$D�I_�-�g����A̗�]�����>�"'
*�jﶧ�x���u�C�i�`����	Yf:Wfe��ް4N^`������"|�
�gx�H�"2�<�a�� v{�(ށX�/��Q���]<_�>�<��]�_�=n`yVa7I�!����$nq�9q������9~�`�o�K�y�U�Hx=�7�P^��6^=��}���p{�C��ۡ�/�^�o��¸; *i���q��5J�L����q��n���	�\e*<�s/|�e�0^�$�5�Eac����Q�5��u������2�+�ߊsQ�G]Q;C�L]�P���v?C+�Y?_7r-�xT�Ό?�j������@����^ځ�2έ#n�3�
�_���uU~?�t�^(��*��B���/��� ���Dd~�E1�n���o���t=��G�,���\��A<�K^@�w%5�s�p ���1|��x6����X���FH����uL���մ����R����i���3weF=�q�?x��U_W.�6��a�J�-��lx�Ӈ�W^�/H|��0����Xw��yh�B���q�(Р�m��_��t(�����������P~/x(�<ݘ��Exg<.�q�|Q\C�4/���~2�7A� �ne<���3�f�U�ݽ_�6�̀��^�q('�&��9E����ƨ]4�t�������]�B�K��?{�<Eج�;naM�/�"�T?2Y� ����U�Uy�.��)ĐRUw��ĝSɀ�Kb�p�1f\0�=����3��Eee\]�AzYG�Jd��<��σ}Fz�?�F>�E�����+�K�K��ի�����T��e�U��D�����(yW��mUvb�H
���V-�^#A�{��H`v ���$t%
�1Q���m�0~�������b1��*׭�4�@�1�G��Jj|����Ęv��G����,hbz�.+d�iP�t�M��2�ġ�UV7�>�w��F��S�[F��i,�����2���.k,Q���8�����э�B�Ѝ���WtAq^3��7�)n�gT�^�N ��!��lהC@�0Jk��o�R���]P�7��2^�t�؍���W�:X��i�ϴD7�42��S<�g��~�G�=6���kpz�s�(s�ҧG��"NU8�2?��*���C��r�Z[�~�ݸy�]�v5�VN���2����]mdFļG[x�<٤��<�&�A�X��/�{�8ذ�9R��;VH-"P$�̦��a=��^���� ���2Q��EX���~�<����zť�Q��*�夬<w �C�
��zU�TH�8�c<م�
_�� #�a���A0�����=.=m���Q���o�L�m��p�����5^���ʤDi��q�z�g�P��'�<��8�00�Nr�e��G�[q��C`࿦ �>@o���ِ!��+�S6�զ)�3�#���V��|�t��-̿�����X���W��c oC��]ś(:u���x2�)�ܦ���?4�uw�:F��f_�}� �<�����Lz/�Q��;3N�$�lPb�3�b��Eq�����u��E�q?�%�}I��Q�K}㐦�2�
P-��*+���Q�4��*�B@}ˈ��ď����ţ�<������;��2��_�DT91�'q%�t�=i�Ώ�˷dH$�E�ŏ�����Cq�%�F�&�0��Jy���^�>@x0|H�Ľh�қ0�M��s�L��8\� t1�<n�w)�ک�VmCS>�m/-*��'M�w�Lc��z���5!q����Ǡ%M_5Ը��SVOH_q*^K_�^p��UWjT�zY�NC'�Y��.�b�Q~�x�k��ݱQKy���=<C��L��7ş�	�d蠡�q����ж�OIS�1d�6��߇r��ߣt�|S���!��\J�� m�	��!�}~N���٩����*����&�&i?���ET�]��͏�:�$T�,#�&:l�n��,�҇��h~���1��������4���Q_��������lW�x����R���=� ��������5�T�A����5�Hk�glP�#�K<b\�ۡ�ƨ1Ь�@\��s�H�ܶ�Jr)���n��6��?���# ^�U�l�L������"����Yp��R�锃�=��`}���c,��x�U�`�7H,◡P�b�F�1����PN�W���û�5:�{����T�keZc��g9���9p,��[�@�"�[[w��}�~b\�L&t����>��rBۨ/����kJoi,ӗ D�Q���4��>�wE�vH=��1�Q��Wٖc|Ւ������~�W�̈́��i� ��C����������~��ѓ���#�ȋ��t֎N����PVve��d���MA|���A�1���Hr@��:+�=�����J�}�n{�w�;�ծߺ��Bt H���c�m��{����t��ӣ�{��&1�.�P�)�&�����|e�]Y��VW��+W���)�����D2�1xP�v�� w'�����m�v��;�$'�B�y�eV@�L\
��mَmd: X7�#Xy�˪��̳���4�� T��8��
�Э��d�L!)���ٗD��y)�a����h�'��;-F��#l�nP�0�����:v���Τ�7����� q�o��T��C�'�2�)�I*2~�Kc$�}�y;�'EB�N��ɒ,�����y\�:�$�2 '��� �նUN�H[q�uȻE2�S揿n���[�¼�g�j�/���<�'�'@�.< �p���9 -�S)H�Q��[����+��C��i�p�\��~��1��w�Y��œ���� �{	�!�D�e��Q�p�o��D	�{����G��z��$]��-2�ͤ���(&�(&�';�s�0��f۵UO�Z�w[��=8��4��pg��+F�g�;[mo{��o���?mW�.��߽��z�v�s�f��*��N�Z�����x����zF>� "c2H�B�&4�%�����.C?g�'��ʢ��[��'
��2?��3f<dn�/����P{ګ4�M���+���r:m��S92�u)E����ͣҩ,Ap��3��RD]�n��������Q��;�+w� �A�<�.FiL��l?�N�1��W��-<;�X��Pn�^�
����D%��_�g��%��k�0@����}Α[ʟ׀��2��]�J��8�Ed�b��%k�r����� i(���>eW�QAR�H]�w�`��t$�fs�mqa� P8���N�����e%t��(�i��^e�E���6�K�x�����4Wnꚝ�ns�m~v�r���x��/y��Ƭ��>#�i�� �YѴ�{�I���7�
?P����G]/--��Y��&t�->�僸K[��[�oӤ9@�2Q�T2�ce:E�T�La��:�$}@am���(/A�/ˋ�ݷ�{��bd�@{Ǉャ������'���M�C��T)�{�����K���N;;���P ��?�;�f��@n]B�]B�O�.�����h�sڏ~fw�����`<�̤�1=0h�t�(��ϕ��vtL|�=���k~,8ߌ��|��P�2�>�,r{���B�y{�]�q�-�O��Z�maa��ܦg<r����\oݞ<}�]H~#�x{���w\&���[����������i��dڍ��.�'�=��iWy�ռ�=���\����~nz]�\���<�/#CgO�O��(�����We1�Cߓ�=9��ʻ��?�#�q�H�϶K������N|æ�unf�-b�Ϡ���3  ��IDAT�q_e�%��2h�B�����R9n�:�a}��m��hЩ+�'���9<N��k��y��P[QG����<wK+���;Y1EO��6�ƙy�.��'��x��	�n|��������-�ϕ��`7��Ҡ}�G�z�2���B�Gn����ē|53?�x>f������4���KK�q�Y�2��^ʗ�O��s����?/DH��r�]�ɪ��0ҁy�k�՜'+7����.F����[���H�yc�ݻs���um	??(��]���`m�0G�4PV��Sa���ݪ�3g+9����� @࿕�+Ynv5�pr�;�ę���v�ޝ��G������{�sP��0�LN��������_�Y����q��w>̑���N�bZ0�,�8jCY�<�?ò�|�B^�-���w��"MO_�yP�qM�s|+,�Hx]\���v��\��ϲ@��`�YN����cll?;!m���Y��,�
4��S����(
��&���ێ�@���@P�趣��K���7
�]��?4E���(�����ch�=�i��x��q]\>w?��7/��q� G]C<��<���]"7\�ak]�/�t�ڤFo��ē�1��s�����x�ܯݩ�^�s�u#�5�7�xiU/��l�xV^@�R���ތ���sA�#r� Y�7p�g��� �1��*�g�^�q��q�F�!��k>��gF�4?�Ю\q��J�I��h.�E3ڒV��V8���a�!��G���V����x���4y_b�H�2n<��R�̬"KM��"������@p�n������ZÊ�Ư��#pI�ƽ����Z�\��iK�D�(G�K�~!@�)��p&����Y%t�a��K�yQ_�� e ���8��0�@�O�~���3-!B!|��a�=��̆w�N%�� ����g/q(w ^u&6�@�f� ����δjX�0���Vwx\�v��Ӛ�,�h�KN�GET����
m��V��0b��X���ʞ0�"B\�2��#I@i�F}��t3u��[�\�PY�Y'��*��])1��㼻T�;m:�N��Mu�8 ?�D�, ����*pƯq��Ē��D���T��Oդ����@�B���Y� L�P�h|^A���z=Fh␏�2P~!Z �'u�p:ø9<��b�ܺu���ރ��o���Bi�Җ���,J.����L��2XYĸ1e��S���|[]]jׯ/��W���Ut-�U̝Du�j2�5h�s�K�K��>'p0z�Wf�Ln����u)�*;UfC��P�w\�R?����k�eg��%<%�U�K��.*�2a%�Tn���8�n����,�'��*�~�#c��q�Ƀ1��i2	CE�m���?|�����	����1��
Z?���v�X�Fr�$����pf��(�.��~��n����9����˖'m2�(OS���ƔA�� n���N��QF�-�QN@�>�]�����ʑ����ʁ�����}SU�����l�20J��������?o?�Ƴ>�U�+�m�7�6~ǣƝ�w��f�P�}O�[�+_M��3��P�8Z]���ϧ��;�&=�'��<Ǯ�U�N泸�Ԗ�V�� ���"��d�j"|2)�A��0�4'����a�\�3��p�M�ׯ�o�B�7z.
�p��y:/�u�T�ryy9�b)�L q�F��/c�޽s��M��G�m�����t<;��[~������o�տh��_�O��~�'���FȬ��d�� �T
�ǲx���b���G܉R��^�P�o����hܳ����H^��X�K��{/�ֽ'��F�H��y�2�+ �j�U!�P�:@�q�K��,���R�+N
)A�ي�Ui�nIq;Dm{8wv��̭Κ%���s�D�y�0ˌ���8(L�c̩p����M�A(�<G0F#�x6E5�-5�\���ý�ҍ�8C^���?_\����_�Yh�	�2�`�����npT@90����������=K=�$�
���27��;Fa֣��w����C6����s��e^�G	���0��l���G�8 )k,'�d
���$�&J�w��,,"��=� ��[��(;�U�f���E��k�V�y��Ix���ʼJ�e_*��R�ʫ �z8�T����+�~��41fHW�L1��M�!]藤+�Y�G�Q�\A?�#���ף�\��UA����>`x7��x4{X�sO�(7[U���:$�:8]'a
wN[S�@�+�x��6�c��%��Ih�����5IV�ݯ�ĕ��� �~(�r,v�5�D�+W��+�� ���G��֠*?G*q$�<�{h�K�n/�
� .�����<6CK��І΄[���脷��<RR��|����W�k�N��*j�;����2��v������b��NӠ:|�������p�J�R1�w���xE�:�8�gZeEt��.�(K��B�:�]45����-K���4���<��T�gQ�<�.��@���k�`�����ۜvF������:��t�Z��q⊟�PY��W�O��#�b;?����kW�ۇ>@��~������?l�������SS�s�c��.ϴW��u���T�2�][���ޝ����7��n�w޺��t�=�w��X]lKeSS����:a̢|��4���﮸ц��=ӓ$
���<��;'��K��mV*���})�N���Т-�E�3Q�i3'�mw{A�'e3�s�i&����wm5����9d�m�
��`!��Qf�6>��2�)���+\��O��y<M�����g��θA��-g���W��"�S�ކw8?��eW}�퇔I��4t Wc'/a>;��?��C���Ly
�1a�H?񊜥�.��6U�|��il�-橡�$@�|��g�A�7�>(o��gC�)��2?r>�W�C�h���t"�ch��ꎎ��+��e���E}�H�z��_s%���I�r���|�Xo��g�O��W�Uh$^�u�2�2@�)g���?��y�i~v��LAVe�c�^�l'�J� �	��܈l5B^�"��9����:�y�����~V�a5J��hx�O�Qp�̔���̥v��|{��n������o?h�n]G���ׯ���{!����~��ٟ������q�������x�2���Uȴ�u*O�)�V�7��89]�{�ɴ"�R��F��<*^�ѯ�j�����4�uq���W)��,��+H	/�G�d
Kh���
	:"���5��U�;C~��/�ǸV�
�
 G'.W�M�!*p$l�� ~ĩ�� �G���G���@�2��5�� ;�JiDk �z��6*�L�-s b1d�N����A�
�C�j㸌���� ���ϳ���ʻ�t{K;��^M:zLGN�����rTy�6���c�iӁ�^�Q��[����܍k^�E}�>��	7�e�{��`�8�@�+:}���P�[���1���2=�k�������}(�]P+'|&P�N�g_X&}��V&�22W��$2�M7H�u֡,�J��J��?u�jĉ, ��3d��(�n�c,�i���g{(ل�5�8Hdp�,�o��r�/>B����b�Lv�VE��B{q1Oh��N�wܦP\|�5ʵBg<τ�4�w+��T^}��2���4m0�}���@��L�hL2@f��AU�и� P�U����\��F�J7�s (�c(����-z�>�Og�ὸ���c��o�q�f�7����Δ�����z�$2�7CSH��ݍ�����j�����m�-�~�r����4�iLґ�x�A)�����Af�i[�I.mzBe�6ƨ(��<�C(�*����MS��u?��9�����bEE�=cm�.!�p��q{��{�`K��`p�P)El����������}?h�;F�����"�Q��k��ǚ���
�&��0�b=�r���N;E��@יk�}���>n�����/�ş������V��e���󶂑u}e��^�ow����.p��b{p{����z��������wn%��V�u��EvW�ܺ��sk�'��yt&?�<���J�
�
z�˥�2ձBw�ڟ�j��}_�]ey�$���R��0H�b{���񥁜v�Y�I�����,�m[)k��A�Эy�l�01=�{yډ�Y�TZ#�$�B����z���(�� � �\�/�d���{�0h�6�PVM�sngw��F����[e�@���2�}2�ֺ�8)�kB�~���I �/+����@�V1P��q&�tꅴ�y��r��k�Q֗�4Q�Kk�<�N;n���d)��K���/y 5T}��R�@�H�(�XZ��A���#��rK?�-��<ƗG�#�xKG��+���w��������1 yByPc�<H^~���Se� 'cl.��|Vڒ�2��)A6:W�60I�`PW�JPVXœ�
٪d�S�T$B��!�����L�?����M�"Y[Z�jw��i�������?j?�������q��ݷ۽۷6W[�ڲ,~#�ڕ,v��1���.��A���@]3���U�Ġ�d]�Wx�_�j$�V<~T�n��-:���WKHØO��p����%R�;w�ª���3E�!fB�_p�h�&����&ԧ�R&�B#ʽ�G�E�ޅ������f;َ�7�W�h�U;|6�!a��WH��Ml*���!VF[\Y˳+a��W��4�bf�+=�C�D�γF�q;ȷE����UO��&}@w�ϴ���6��?F������ߘ�6�e���%
z< U��x������Fm<@@��RA�Q�e����Qޥ'�<ﵢI>��":��o�&^���0��4�6���ob�2��U����ꊼ�Ц�g��kW�P�ꄣ2���;��g��
A��<;;{m������>��3�gݢ0�n�Bž_Je+�R��� ����n���h���@	��(y:(9���u0�p[G7�X�$�Deo^5�]����@&��J���/�}5k4������@ݍo~��`�Ui�c���э�
�b@�VH|��sfZ�٦u;ω�`9rf������e��U���tšVu+{YU��>�� ��%�!�?��0n��(�A@�W�kd�F�7�
����Z�x7�
u�4�)r/:W�8̓m��y(�~����|�{�r���V��|y��?0U��%�gNW�־B>H"�)�L|�Jk:?�@7���i_��m	_M���誼(Wr��+�j'Q��р���ދ.�t��!�Ц:*�Qc`Y.������|C�K9*]�}о�X�>m�m�7��}�:�R��-�h흽����β��t�4�i���꜆����^�u�E����q��	���4��ɶ@-�������Go���w����������^k7�εWg���s��������ݕ���k����=X�J�+���+�[�
���T����S��)F�9�tqg���Smee�]Yqk�ʤ�
���m�KҴg&�ԛW�J�ڷTHm�(���[�W��? �mઇ+����k�%�Vq�p�E��郂<7�!�(W���2J�B&mD�j��#g���5L��ޫ?� ��f[wq� PM��/�:��|'�#���ԁ����&3�!��i��
t[�����1G�Ɖ�� o�}���{���(�3�͈���v\"\�P߱"��_�o�1m�ŹƲr�8�C��٧�� ��Y�ƭ���y��X~�V��:�б>d�;��ڄ�����`_�֕�	����C����C�B5y�M�l
y����US�c=�h��_�AP[����3������È��v,��5N��K�ۿ�?�r{��=z��>~�^�m����cZ4�jp	�r�/��3 ���𤳩�Ұ&	3H�!+�{2D�$�LS�xvܖ��ڽ{�ۃ���X�2뗞a�2�3.Smyi�ݻ{�=x��v��Ͷ��k<� �zp_��x
@A�C� )�\���O�&1��Ɩ�shmck�m��P�A�˄�m|��/3�4�n���ī;�$�cW�����y$�б:�0�d�;�LL��)�J=#������҇.@�i5@}�*/_�ve�ʐξ ���7��7����N1�N�I�bt�.8>tU��_@N�:&��<�|�%����1W��ϗ����+��0�;WIG*��"���҉<����ݒg��b��t���Q�L�pۨ�� �Nd���^C.y(w\���W����������e�Viu��Bܽo���g�9L�P�o�a�C�`��!����p�:�U��[N�����QwT���=j�?p)<-;���L��
��WJ�l�AQp{��THDOH�(����L�����`�3��N��p���\��nܸ�����*t52<!��/?~Ҟ>}��g���Yf�{�ʋ���d���ٶ�@Օ�}Wܞ�TG҂/��]�~�)'�p�PC�Aa���I��<�����(t;�Ut<m�Z�s �w���G1��R�X����;J�^�$큟�t�t��z۾dx�]��6�t��֖�r�x��B�"
���*9*e�5�:���=*�����q�w2���O��RDj�� ��àH��kye�5�����K�!>�;]"�����O�H����m�{m������8�)���~&�]����[5~-��p5�`?26��2SM�����S�3�]'9b:iJ�$m��������6�@��
{̶�p�ñU>�,q�w�kW4��7��W�)8|rB��.����Lx��R���sǃ�K#3����Gf��ku�ʙ�[�=-���q'X"��c��0����{M�o^owo��p�_ԟ���ŋ���Ͽl_?z�^�mP׃�!��F嶲ZR�`�`T-�]B^y��,F�|�ze	��\YY����[���[\�nK��K�C�8��L��'����Ƈm{k���|�vw^��1x��([~���n�,,R.�W�+mC�J�	e��-,̵���lt��zYt@'�l���������񃺮����漢=�-�?�>i�Bw��K��L�z-�G�����yd�ۀm*oۧ��2g�����1���@>M����U��P�+K�kҹ�&��6e�G�Ss� 3����Sn�ݙ �;��$�<l���LuQy�t�Iy���
��ݝ衙|#�<�1)����U�26�����-q�#Ǔ�&;*ne��4����u�Ú�(+㇄�~O��xnP�c���?��9n�x5� {���LL�HY27�|��-��1`Y]��_ʌ� ]�~j�;���1�-�|������t�l���� n��Ǿ�7+3��yY'��Σ>�K|m�u|�.�4��t�F���%����e�[���~ _�wY�||���*�ɝ�v��5��}�8##�F֓��K�,02�D��N�'Ȁ�ʎ����Ȣ�Tr�w5 ���p���b-��)|�l�*���F֝��[��¬J�
��׎D��~���hW�^C�]	c8����5_O(�qN%�%F�C����΀#� cq�mn�m����#�0|�F���"�$���LDGɏ{)�@Fq��
�<���;c-����F��F��q�Q4���/�ع2K'�9S��jx�m;}PLkŭ��1�b@Z?gl5|4X5z4�4��1�0���]:�|���A5�u�K�j�8��3:dm7��:)*�*�/�ЭYd����satI�ڦf=l{�g'����uVŏ�����JMy蟎��0�D�<������~r����⪰�ϼ�Or���|F�"|�0��8[�<[�ʡ�W��^���8�q�����C���a�G�����7EVo����!W��鑡U����������I_���@����6w�Ei���J�<,:+�3Bsai�]�ve�*��B�p�S�}���=zҞ=�{���N�Ё�!��^PQJ��yp^��gKx��AdDd�"R�A�t^[��n>�6��ug�@�0d��29�Eg�,�A�8�R��42T�Ke ���r�c�90�0q�R	�^	$ˎ�L�,��;3}ĥ*���A?��?3��[VY�@�P	�Ǔ��Kx�v5�
����O���(�Ӿ�C�w�� r�� c��a�*r�d��S�1��L܀m��q �~%�*�Ȫ��V5w9E^��Ա䠆	r>}��(2�v���� ѐ����x\�F�)�I�m=�'���M9�PJ�mO�b@~��Xc�J��ƨ�V	q�W��<��<��x������.��A�.a(�6���7=�V&W8�h_�j_Ǹ(U�Q%�pr��\��l�������f�j2T�:&�o�;u��9O�=A8�vG��H��$��g�j�{����W���[�&�!�rE���g�ۧ�}޾��a[[[����W���4�y��%�XjW�ϹՌ�|O�C^©�^>���v6����H[�����@���#�b�i��x��9y�1�8c�����6�����s��������UM����3��6�.�^��ж�4<�bei���*i�~ڧ�]@�����.��}�ѩ�<���y�d��[0����ۈ�Sx��	'e��T2�m�f'�qr��~��|#o����_������K��q��q�R#K��<xg��NNB����G�Ƌ)e\yq���]��t�U��P�F���Dq�d�tUOU6z��<�	��}S������ɑ��Sh��Ĝ�Ǿ b�G�����=�����d���&)�ԗ��z5���A�Q����Ǿl��n���3��:dK����1�����/cΚ��t����@c�P?_�в�	�s��Yzd�	eX��xkdv�1�m�B2�9n)�B7��uޡTf�(�c���l>����>ȇ�~�ұ�F)�Q7�[X�|d�����&O�}�*6��~V�__Y����s"�N,Y�����
�*&ΜefցC�'Pĵilx�Lh�)M��"��X����ݿ�ܿ� ��� ���R1���y"Tb��נ��J		�¬�c@�/<��I���4
����5'1���.�󶏑yr�����_�pt@f�C~Cg���z��������2uhz�c\\C��=Й�Ԋ���4�o��=@�����'��p��FF�ͅ�3q>G�{���aUR5�4�#��Z�"M����:��ed�7e*��e�j֠�l�R���� )\ʝ%��+�j%��u �`\�1gS��eV(b�K��q��������h�J�x#�W�����(<V_Կ��2��V�ĳ<y�?t0L?�^��>'�(����^��vqU�����xT/��|�o ���"r��s�r�_,g�u��YaJ!��?�P�r3��Ҳ{�<X��b��Uۿ�.ΔϢH,�\�g |q��R`sk�=y�$3�*S�� b��~�@ڈީ5m�8���dE*鐥�D��W���]���B��T�Vu��M~4i-0}+��������?�����m�ব�`Eʱ\i� UuH1�'xQ����HY�ATH����^��C|��6F(pI�[~�����N�<8�f�7�+3�l��@Ի�%g�XC����#��-�)e���J�Ȑ`0�]�G㍀���x�M~�9��p�1
�N�r�������Oê���F��8���w��2A�F��L�wk`�k�dּ�Ld�0�?�x8F�X�w�;#OɡQ�����QO���������cª�:�����
�}E�T��r��D�IY1n���|G���	��6`,� .u�����$m^`���z�X�{�MB��9d�ؕ�{�o���}�����v}�J[^�ԲI���%��/~��Y��7�W�\�>4#�������{��u��?�����JR�ǄKh���g?���Ǔ/��qs��|{��.���v��d�p�Zeq�mmmf�I�e��W�kw�>hwn��X�F�K���5��Q��������A������b��A�I7H=�g���M�$��W_kd�@a�t#K��2�oJu���K�)��6���n'��<�w�جr�m��PYV��� y�s�Q�����H���Q��<������f� i�)�u��o���)m)����X��� ���ȃ��>T��Q�Ϥ��_�)�e�~*Ic���%/ٯ}'0�>������kߓ/DS?�|s�2�ׁ�SpO�^56@s���e	��@Qd&@5�����QV��B���$�_ŧ��7/��cI��1g��d\��1ѱGy�X&^14���m;��yJ;e�qS^�is�@�C�O�)S��ɁK������#���R��r���Z�j���ua�v#K��km��b���r*뛍,���T�]L<�[);RN�!�3�~� ִ���� Ⳉ�<$�Jρ߾B����k�Xw�}��y�����X��*)0m���L&
�):�9��b����\�  ��x��,��o-q�>�b���1i5�v�Q�����q�;��E���n�������1�m����R��I��p��ֆ�#���e� X���
��(��Z���}{ C]ɗ�m�1P�z���U���aE��8�VP��Ej`�UQR��'h\�������"#�ΥT�K�+��qEx��Y�Zөį�Xn'�v�
+Ғ/u�Z���w�k�H�m���i�s̋ �n�9�N���d�����O��"Ou�/�jϊM;fV��zx]:g��W�ÿ�0��t�O���+@����4���P�>��|.��o<r3M��T`��{��ǟq+d�G���W�|���)���/��B�ih��H�0?�������X�K���O"��I�A�\�Ү_�������g(_~�U{����"��c�
�X���� ��6e�O�.��h��
�H:���}=�ǐ�e9p8�Pc�ۤ-��t�Kx_��L3up�_�+�z��r[�J�����������d@�u7\������als�����'�E[�� �J�/}�� ��;!�?e L�E]ޘ��OAɨ�!%stT�ρޡ���%e��1'wq��t��Myy�3��g�>kA�i����H$�'V<~�I�ϝ/l7P���d;^�L��B_'H׍X/����������O��Q�D�W:��(���o�5n��Aisp�)c�,�芞��M���v++R����	�u�Ji�D�:	��W�\�p�º��(Ϛ� K��E�`9U�Aϰ� m��@W�UWX��ރ{��ￃ����^] иkȁ���'�������#����v����͜�^^Z�*�������~����377ޕ��țY�k�x���{]Y^�a��d~[ȃ����[�ٌ�ȳC��],��Q��WU��]��F��g�i7�;�O}>j�n�#��}9tp��X��vt*�[�U�Y���@Y�����H�g��z�ս����˵�`��= 䨓��u�U~��$�}��J�jb�ЎG�in��d�G��diV����D�lSE��h�dB�q��S�����x�D��WV8���S<!���(f{��$L����,_K>T���r�	�������pV�;'YD�0i`���oY��93�x�b4���ykwFe�1Z��՗�ku,�.�p3~в�X N�E�+Y@>��?ZO�T&ێ��|��m�hPE��.1z���J�e���,����?~���*'@{D'��a�6Gތ��/�,�s+,���2e�)#�,74�_�+$�.�!�r�������3�G��w����n����6��;��ͬd�q�1�<� !��h*�<���$�{Y'P�ƢBVֆ����V���^�w��߻�f!�8v��Ν�%ꬊʏ�)s�1�~K�l"o� ��Wɧ齙�	b��*7$R�g뜲��F��c�u�pq%+F�LV�&a�� 1��`���*O1��a�yy��j�6d")�#n�q�1N��DJf�3��QT(3���j�"3�s�����T4�Tn���U#c�)o�}+�,��=����!�P�ՠ:"/�J�[�8�G���U�Z��x�P����KAS��LZ���}��
�l3HgA�IʐY���sz��*
���Qkȧ���
���C|�URü�ߐb���\��{i|���s݇�
#����^�����A4ٕw��#E͐T���櫔��+i�5�s����5��#Z=�]?݉Uφw���yF�O����r�~����O�RV�s@%s����d�ھ �/��H���?h~���v��-��T���j_}��}���ɓ'mwg'ʰ�z�zq�/9��?�:�����6�u.�6�o��<+m噴�S��:گSH�9�GA����=�S�ǀO_��l��AV�m��}ξ)��7�_y�����_��o����r2������*H�u🠍�_���pט��(�8@����G>$_yF��D���,w�/���.<�2����xt�$��~��L��/e ��Z�7�Xv��=2��$)y.^�I}(/i(�1l�˥d����<HS
�tw��_��^�`��Hq�B����W���=������D �U|���eͳ��2ȃ�U�j�K}2 5F�� r\vr��t"w�F�@��L]d���ގ�V�B����A��|�#i�|���t�)hxif�� c�+�d���z���1��c�LC𸭭��_��7�����Wm���++����++�{�����������C��v�w����Yׯ����z���v���r��?w��+�Ȥk�O;ދ��턾D���L�W���%'�����u�=2rv&�W��n�����ow���u9�����`yO��l/�Ȼ8��լpYY���e��I��-T�G���ўB��O������r��'W���}�ns�T����逰��D�j<�V�Qv��ĝ�&������Ǩ��!���I{�+��79U����+}��E�W��Rח��w��<פA�S��'��?��3�c?M��Q�?����˕/�r�$9�GVj�������]�*"w�Ӆ\O��Y��1�� (,�H�������㬬����a���Ե��i�C����1r�1���,/�Gxԅ�&���xJ�2n��Q��{h*���X1�] ��1�CW�p[���H>���ץmv�>`�v�^c�#�.G%��t�Ed�;:hjss�J{���|�N�k�;��.�������흣��Y?�b�	f>uFAև�e�W	q���8�����S�$+rVJ�������U�6n��I�^Y^����K���X�~�ܙ9����tas \�P>��xw�S
�60�b�-.��g��o\�����ɴH�(� L"'1��0���Ξ{1ݓ)1�lx�B%,u�ì�W�$����;{bW��;�$6|r[�0�ĭ�cv�3���D���l�N7	}S�e(zH���2Gڑp1�pj;��0��`�sW���� ��s�����D�����6]oǇ��`��r?9�"�2ܣ���К���fݺ	21f:�Y��H3�`q��v���v4iU�=���P�Xy9p�By@}����0y���+�~��;�_�q���ߏ�$�^_��S�C��(��:��:���S��]�pq��*��m~O�Jq�h.s���M�ׯ^n~�y��C�@Ņ���>��B,��mMX	�j�\����D�:���'��.����tHY���N������s�7~V�r����q�뾩��ɻ���{yJ��6�"m �a��ig��y8��*V}��}�r�	��c���F�1
Z��4t&8J�F�uō�(;��w�y;@������}������?k/�>i'�#��\�w�K��w�S�H
l*.���'<����ʺ3�Y�.
���Жp�*2���`�ʥq��>�J���Τ���/��"����~�ɒl&NʊQ���ݙ���i|e`&W��8RN�)/;���7�(E�Mo�X��9mJJ�i��Ų��h0.�?!Ql�@�U���m=�n�h+)����Iޝ�������&-��se��*0�rB�X���qf����	?mS�%��EB��	�@^�&�K��v��&��]�1�	��&���jY71q@z�3V�n�5�jZ�L�t@�(G��9%�2���ϑʓ�� ����t�Ę~��~z}������a��,+%T �;;�!���2m��|�!t�B�C;�۲�]
���6>��G�w�$a���U�I��+٢_�3�CK�'��=	�J�>=T��Gx)��Gmk�,߳v,�dx��m//_�(n�S��~d|��7����1��$�v��J{��{��w9��D{�lm�/>������h/_<C��n�G�3�c�+Y��o����kmg�e{�������oR�y>r�6��>lw��k�</�η���ve�*p�]_���v�i�-���r�B�@����y�9)�ι��Jzj�,z��͑�����FO���v�3夓S6F��b����t�곴�����w�˱@�y@�lmﵗ/�����=tJx5}Y��`�'�������muD�	�S�R�G�TP#����g��6�mow���xZ�6a�{�No��'��+������=Y�rc�-a�������㘾�d�[���4��lm�c��*��M���d?������~����5���x�:�?mc#K�R�+2j�>��z'e�Kv ���)�A��N�r�r�{��VLpCW;B�;��-�Ii�i������`����T����7���ދ\T�?��B��_yFD���j�FϬ�F��}ж#N�R7#~OG�����x��������u�[����!��(�G���Y<p��p`�g���zM��6���n���
&�	8��y�߉����F/p�vnY�6��3E�L�k��t��<��޸�ܹ�n]�B3Ӗ�+�ۿ���s�=yY+Yk�d9��Q5�Ҽ4�ʼ3�S �� ��@�m$�����WihEH��0V%�R�L>%�`* �\�
�q�z�(�?������]�r���΀�(�����0_TS�z'���5;Ge���U!��3xN�����#��/���X�����rx ��^���a��+�↑�+w�:ϦOb�윹�g>����Md����<�}��1�5O������})�v��ȭ~�����Sʈ���w�J���� ���4��TrUvK��%�ڮ��� �"!��&�C�U�;d��a��5�	�ze�*i͓6��sEKR���u��?Ǐ��"NJ!�jkT�@P½R���]�9i@���>"d��>J�^Bŏ�(�O��-��Fg��/m*��j�ޔ��z&�W92+��0��_��NY1�盗~񽈖k<��tu�W��SK�Tl�j���=V���\���qh�oi`;+?4l�OO��̗���wY�K匲!���s�l��G:��,���|IWYt���v���v��md�t�Dz��i{��q{��y��ޡ��(��a`���P�Pge�u�Q>βe��2Df�ٗ,HXJ!~��ۙӒ�%oS�y#Q�yGxU��?�B��Q���c0� ���t�g�k�G~-C������W�%�*����z��˼/ʕ�KzT��׻�G����ZyƂ�����= İ�F�e#ws$1���5S/rB�H|R�>Tֹs��C��X����m����V��356̻Oƈq�"�e_Z:Ԫ����c����Zk$R>yQ��l�l��JK��7�l��BZ���O1`�9�t��ɿL?�*'5���l����A�z��1���{)�LxQdm�q��$�q�/K�&����=����K񘔫��qB�0}N��n����#]m7���r���\x��;o�ko?���{;�>��~�����o>k��k���ξ��6�j�[�<�b�is}�=y�E{���F���)�7o�h�z� s�\��,�U�zg&�E</,, ����C�|gT~Ӹ�0���Qd�fE���=͋o��]B�?m[[���ګ����~*�0������ƶN������g�[ ��й���d��*��������0<�JwGM�}+�^켪mm7'��d��;�Fs|�5,T�/]''�1�N�<m�8�k"��q��B|W��by��R�}c�ݹ��n�o^[Y�X��44&,����q#�6�w���vsu9��\�T�+n�D���҇Pm���O���zʺ}��95r�ts�P�IW����{����VW���zͶ�K�zi<�s�|�i��dg9�n]kwnS�������,Xxn��!bg��w�g���2��b���L��>���.��~W��-����.g{k�i[�Z�'��SA�.�([+���%�'�}ܩ��ǘ�>i�x^�˾,�^w?���D�Βn��̖ٴ12��!�_��_9c��S�cc,�f���U'0���0ˁXޕ��a� @⿣xi��!�{�iwϐ0��՘N��O�������^,O�𵽣�n���w�l��o~�~������q�9�#xRK)��a5	Cζ���62{�t"�8lGζ�4�U2�f�N�b8a$!P��3Oɋ� �i72�����ŏ�;w��J���@C9�Agui���V��f�G�K�{�gc�p�����S?\|����Q8�0/P�0a��{Wۻ����x~���������n�g����.�ב/^��<��Pp) �*���)�S�_p�9�(?b�0���˩I@�w��}�)�卌m@�ʘ���p����A�	&A`�1� ���������=�O�*3�t��H�<��x�E�*����?�Cc^�N�ė��\Oj���K�fhrg&�Ze�Q���Au��W���+���2J]'"ט�]�ȳyF�` � �t��n@�(ovv��\�I�0���O!߅Q��e��y{�NXݡN\�'@$8ú����K2D��Wв�B�:����[u���[~�`*e��q�uh��i��"ޕ�<�S<x��cI����&��.q}�R�κ�2,q
��x#Q'Ő.y���D-Ή	g��Q���z�l��,--��W�(!^��g�<]�
���3��r>�*�G��::���|���w������}����{9��˯�h�𓟴����~��Wk�m�Ke=uW�������O��c»m'y�z)��a�*��i3ג_��/T&q�pE)�^�7}�2TD/�����C~�c��y��!#�-\C�r���6���NWWHc���U��0�U8�qٟ�
.��FEZh�� L�c���yJM?�p�WYԽ�.�U%'r~�]P�+�W�'}������?�l*�-ct �?�P7j_҂0���>I �D݄�"̅�����ҝ�����#_��M������9���։[JMpJ�
�:Dzy�J��O;�S�`Q~T��H��d��n�u�)���e���*(O��ݬc���r���u%`�1���z�� �L��/�4V��eDW:�ob���.�K����l2�ɷw��As	�F���a9�pW���:B�G���\��Z9����jN��:��h^�@�n?�އ������������3���o��h�����k��?���~�����I[x���c���P�W�[����n�8�̓N�1D�a�����G�|��9p�my94���n�V�b(=4J�۫W�׿�E��O��}��ox~E��P�K�eKgA��|�'�Y��I�D9��'��ݶ�j+c���9������֦F
2�Ѹs���{�m�WSm�6X^Yls3���U�w�mcX=~���g�l��ͧ�%��B��s�s��@�e�>����t�V��<=�b�^�}��Tp�+O�{��tѳ�"��,G7NN�s�����X� �z�j��],�x�pw�a$�o�����Z���\Z���ܺ�j�1x5h�S��1�y������ï��W���1�w��\���s��z[���(���|Wn�����g��㇤[G�_h�Vo�[��}�|�8�W�w����������	_;F-��..b,��{�����ʮ��/_���=��~2/L/�?���$:�n����wy3�����,�Q����B�ԥl�>�ޟc�1³ˁL��Tn�(b>�W��#���}�����N
Զ��]�����<�����z�I&kh���vD�K2	^�ϻ��x�����]���gg'��l��K�W�%ON��	�&0��u��c����PN@l��7^��y�޺w�}�[�������w����|�����F�I�=�s"�{���-�XK6*�r@�o`��#�NbGp�(/�wv�׽��!Dt	Ud]�{���v�}����O�G��ܿ��9׎`d���6~�fC˙�w�y�ݽw�N=�U���-�Ţ�k�2�3��5;E�1P�q���"�����s��I�JC���/Oۗ���|��!_0�`���(+g��2�kFV����I/*zb���'�`d���0��1�p�)s�p&�x�
]�>��`nU�~� ��")�80�=+�S�2��d�����pf��q�e�"��>[m`�K��Ga��)�r4<*�D�)�/O͓W�,���I�ԋ�"-ӗbp�F�s��(hd��P�QE� .�M|�P�?J ��1�>
?�Ihc��Y���2��\�ns�'�$�r#뺛kfo����I�R��Uq����Md��e����>�h��s����~I�U"E� 4��5���H&ÿvUz�C��k�o�ׯ�n��m���e����8͘��z�2^n��m_�>��x�0N.À�j�_��к_��ꇨ]y=8�C�n=�B#���o�x\�3Z������O����28�_�쐾�>z���s�V���ؾ��o}��u/B���G(2����o�������|�]Bo����]EF��lr�q{����"���(Eg��o��gi�;*S���\(j����]�
-UʕWǙQ����g]i��$�h0�v'���2���}��I0}�0�y��`�/w�@���B����Њ�83�?���SoO��W�c�HC�n����}��g�L�����U�!<�xňJ]5n��4F��3���E<��|3��D�����T�7#�g������W�pA#�D����h䚸Ǜ�*.�<�F^J~�W�h��]:#~d�Dr\� ����b�S�x��iX1�����/�C4T�A�Π�y�"��Ye�����*� 3u@�A7����{n�Zێ�#�Z�s+�����G�g�Q�(����*�"�,��_K�4c��
s}'kn%��=�0��9��H�O kO���J�D�.������?�����uw�-�"ѥ���Y�����_������?˄pY���w�\ź��\�@F-���Ab����~V��y������}�ݶ��~s�OC8~y�HR��5����v��'�l��������?o/^>O��n��&-�s*���U�X�.c������~NV���{yp�����v{��J�6t�X\Xj׮^k7o��!e7n���y�sug�����P���k�?�U��O��=}��|��1�C��# m=����C�2>k�--]��}O�~qJ[xꤻo��:���$F�B{�>8ݽ�睊gh���~�{	�������?�������O�Ͼ�
��m�t_��5o���k����<mA�~���tY�|��}��g�������y�����[o���n����C�T��?�����z{������b�=�oWڝ�o��߾O���[i�X�d�[aw���ƴ�(��]�p5QC��{��Ή��`�s����|O���pW)7w���拶����#�0����>JS�_�;x��B�B�h��-u���.s,E?$���ㄆ���|]��W��.V��e��߶'�����D���Š"/��s�����nI�����d�O���S�]�t}�7ߨ�V髯�K�=xh$�O}�һ_�a�]��q���
h{�qB�h,z8ߎ��ol�͵W�����Wۃ�7����ut��K_�ӗ{��_=Zo��'�j�������i q�lYub��ΥX������a0�{jO0��m0�O4�4���X��?�ײ�e��0
��۫�~�����o޾���!�˗/��~�֩�F�����>����[��R)'������+&_Rm���Ѱ�3�Ч�e rb�U��Ȃo۳g�1���Z#k3+Y��1Ď4��F�и���4������-���?g��(�m}�kF�a��4H�y�n�dj(�˙�ʬ8�P`MMNWz˷N]R���Vg�]�ʉ}�g�Q����x�`��(�T�TRTO��SHp��r%���,Ѫ�b�8�7��oe�CK��.���C�*����T�|�*�5s ��j���8T�T��T�qi�m$��@	�̮�g5�ecv%����7.1�L:�39K�
�%���DIh��W�R����G�hx�Ս,�1.�%&����Zm���+��� -�$��Ȫgi@�
��Y�w��������!���z%�"���s��Gy.q��$���7v�<+>Ѭ����r��� �d�A;��f������+��D{����:W���Ŷ�&�
���V{��������Gs�2���1Ԝ1�F����;���O�����(�c,k���׿j��w?i���?i�~�Pw��Y*�ֹ !a�ϙs%�<;������I��g�\�J"�;(9�p�ď��*mk�4=A��G\�s��E��.�e�QV�� ;C\[c�e�4.�Բ/�$�ߛ)��O�G=]y�OG�V��ϣ;�p/۷�<wF�>j:��x�Sbq]�E�w���w������|[�(w�C��>�s��@�R�����E�����
�WX�މ$d�3�a} ������W�����>�I6� ?e�:�ZMZQ/iAX� ��`���G��S��n'�������.y�α�$��ip-��k��I+���|q\��<�!d�������񎣴�]wa���j���;,�jÉ'9�wp���4
�+*t�~F���n/���E9���Di��KK+(�K�J*o����%����WQM��n�0�2
����%k�#�A��-�O�z��i�����``�������p�-�3B����FF�/~񫶉���*�
~>x��vuy��A��������2?H�rM%�%�N��[����]�q��,�'
m��^ڷ�^��=��W����߶_���Q>�#�B�o���.��Yhhi�^�(��^l��W;����9I;N�|�g%k}m��܆��퉷0��adݺy�͓�"y]��C귪�5�;b�Q��cd����������'�����a��C�^�4�vw�0&��hs��r{ە���y��Pgmw���b{��Co����n�����w�ի��e~3n_��Vi�{`˄i`9Gs��4_�>;>k_?����=O��zm����N��-ͪ�P�ۧj$}��Ü���h�jd=x�v�y�
���6G|5�CXvcs�=z�t_�k/h��hd=h�n_W�1i���eY�-u�m�j7���mK���Ճ���X�j�ƃ���o�m�d�� ��W;��K�f��C��o����:�rӇݪZ;�G\ Ah��;�Q���w����xG�k�{J�+o�.��o��ڂ��9��Q�WV��CY�l�ߕ:�7L<4��1X��x��l��|�zm`[c94�n�v˹�,sL���J{��媔[\�h�	��Ex:k���\��9>hd敁���Y+��53�3��f&�����������ͭ������գ������j΢��\5h�d�}R)O	�|g�ܦ��*����D�IQ�����*��!�Bbc���g��[7ڇｓ��Qb~򓟴���7�k:��b/'�p��C�G�?��O��˨
2�vc�X�-e(L�0{�j�"�0��t ��c��}�YJ���E)MRj^51����U�3x�WOH
<�Ѕ!<��(�i�!~�wض��o��޺m1�U�Qꮺ�<�#�������tV�1�|Y����3E\S*�մ�^F�]�虚�|�p�U�qa�9�fip�֠c�7�;���hkD�335�/� "t�RR	��V��[/��/�a:��❲�6�@o�F?����8-�v�%^��ܒ��J�*���w���-��,�f�u�Ío�J�=JӀ�k��x�$�>�b�/nuY|��_��Xu���+���C�Q>w?A�����G��:�rFa��/���:^����g��V�1@�9f��3H2_8���Ŷ�6�W�X����E�8K]���#��ð���#����{��m�'xݽ{9t�-38Lc�� �]�W�󽋵�н=�gh�d�΃�U^: 8C��y�|�h���\$�ٲa�Ⱦz���d���\i8�XNf�8U`���/�uĻ�4��߬q�5���b�18H�dI&1�(��*���A���a�$q�P9jj��K�"]���N��q@�eJ��z7�ܙ�&1�&Q� #�RV9\@uƋ)�ʝz�w�J�=��2�����=��*���Ϟ��;�S��sB��2�>��׻��Sdi@eϲU���� -� ;�z��
9�,��-�����ĵ�)'����MA녆N
�E_��,����RB�	�9V�%�����L��}4e��?��Ƽ5f|a��%��h_\\��=(҃��:}B%��ݪ�6*�bģd����i��/-��!ur}����h�>u����)�N��W>S���a�����;��o��O�.�	�.�+��
F�����;o��D�8I~_u�O~�i�����,�O�X����Z��N{���o㥢��^u#g��!V1f�h.C�� �}l 9�$?y�=��a{��N�(yw��K��N+n�x$�
���J�	2m���c�m!�WM1�)�C�[%We܉r���G^ZX��i�ˮ�ۥ�I�v.Wz�5Bf1�r�>��]7s����h@�n���1����p�M���}� >;9���F_|�~���i�۷?z��M��N��kW7V��^�񵲌މ�8#/A�,�VN���$OK�u�zމ{�-�����߇���a-P_y��n	�֙�߹}�=�w�ݿw�ݾu��)Wh[)�D����zOIC��j��i��.YzW�4S�[�g�Q����֣��a9�����N]��Q���fi��/e���"<�@�\����Iׯ���n�{�&��j�ﺧ�6�&4�	���U�*1�(oc�ާ�܁��{��	��ܺ���]�~�4sY]5��E����*������3NI/�=��j���HcN���y�nÕ�+9���w��ɟ�b����;�(�F�U�o����uL��)34��zs��u〣[`oQ����z��ѵ���)����bV5�=��[�R�����HN -���_0���_nl����X�X���H���R�ڙ��Qt��k�,��_����BJ�F��3L!������s����86�G}ؾ����8?{����7��4*4Z�n�qV8��
�a��ܻ=����=\R�^U2�{�P�d��>�������ɂ�X��F��W�u&R�C���_�J��N����
�"�x�1���܃)�р���`桷w/�*DUa�[FDuª�4.DW,)*�+? �Q%���;W�_�`�&�/�������
C�V�H$3zD�4
�̌_}���X
[?N84����D J�TE|ů�;A��{*v*�*lj����.T.F�P{b�]����@�҉� �D����>���H�e�)P�<����3��1�
�z�\�a���P���k�Y(>�^��s�өH��T��wEC��_����5��M�ףp]����<$�y^+��������x=:]F�n���JB)��ʣqo;5W]�H8Q1@�%��W�n�,���
��mhd��ao�~��^)P�ߗg|_#�e�U���;1��0P��)8����E`���l�qu>�4 m)�=��"�b��#�s��U4�i.�B����2|Th4h�M�D�j��N�d�g����3ۨ���M��k�LYNu��?�\��V�9]k*%g�U�T�j7�L��mh{IW�YN�
]4��K�[�a�Eۮi��7y����u��"�TN��<�{�N��b��wܗ.`�`i�` i]�`L@In�3<�@��G���5�3䛧�M0p3��O�8:�^j������r��!���xZ�y �'�(��P1/c��b�i����	�M4i#_��=����g�Ѩ���\��U�
8���$�G�h/�Sމʏ+�f\��������m*��+���|�o�q�O��"a�%qF��1@y��Ã�F1�ڜ+L�nY#dPy�/X?W&�B�$�����z����X�y'c8x:y�V����ƂJ��,�:�Sm1�?Puw%XC�J��fz�Y�%d�"�p��!u�����S�t�c��(�|qu���o�ə���_����mw� �Ⱦ�jˤ)4R&�D���D��?Wٔ)���P&?$68۔ѩ�,}H��W����g�ۋ�O�2a\��u'b���R6��O��mW6������;T~[*�Aw���C�3J;����
��=���+es�mCH#kEx	%ܼ�9��=z��}��a��������'�OP��o~4����������4FpV6�My�?�u�WP�?x����}��}�+�u��u�C��� E�)<t�	y'9$�݉�Unppk�"u���E�:�_�Nœ�3�S�$�ʡqv��h��U���Ne�LR����[/P�}G�:��5$��SN���M�^#��fJ7ˡ�MU��rt@'s�n����\u��2ل�����JeĨǑ�}�NG{{<�:`9�x~&�����bj��6FP9�H�����ZH�x���H9n�w�^��Чy'���� fh��9�>��/[����j�U�+ԅ�Z�Lk��]��Y�f{ ^O�g�&�|�����4K�l�<HFC�+Q��˹��y���]5��������2����c�DN2N`��0n�A�ҝ�������^3gC��̥P(���@�����5#*�Ȥ����w�i��裼�����t�X�X�2�BԴ*9O�=��>
<�mo#��$9���h$9{�d������z�:���H�Q�� �������U�(��W�}d��[�0���}�S�������=�cf����,s��K�����*��[����"xz��_៽�+0+����v�Ɲ��8(�"D�]�0;�3
�`��kyi�N�G�a�E�nے�� t;��ˬ�Θ2�qG�F��GO��/����#f�0'b�%�ih��Q�>����ݴ�q��[�=�ӭb4�F���*�]q��b(�|!u5"κ�s��r�. ��?I������2v�R�U�8x��E~��!���)����$�.�~���c<������>�C�r�]����w��Ah2J+?���"!�R�Q����W�� ���� ���,���(�B��2�+�88f��lf�+ӡb�ÿ����8���U�v�ȁ������r����g��n��+O�u��s�_��^Ż��U�l��3�'�:\v[R&@��]a�I�T_��ۖ?n\��'-TB�p���u�Jc���q�JHe��;U��p�'��<�c�QRC�m[ӗO	SaNx�����0}���~��3���m�����O�Q[�9nW�����v��t�wc�ݿ��޺��޺�Zh�o̵���ڽ�(�7�r�]�i��N��W.��gmyE\�=f�=B�R�40un��{Ļ��|y��#�|��p��e���A�Y肛����	�4�!��er�DW���	MOh��q����o
i��z[m�!��َ%�3�`����Ћک�@�;�a٠�GK���R��*������$J����-�*��c����t�ʱ��p�
��ODY��cF����[�"B�����sp���3�3�rYl�X�FdaNr�q~'jv]GF�oX�+-�*k�q�b[8Tt�Y=``��Z{��q%�X���2�讉aqd`&yS�����+�|?���EN�������F�Ky�l���ہ�u��>n'�"C�+���;i�t���y7�|"k"�
���;9�ε��lgۓ�5���%4��	�d�\R��}�Y�]%uӉxZc]��_�4=��:rJ~ ��;��
@��l珲����g>����l��
�W��=|7NCPz�dEhC�����h'M��;刋|�����2��Ut�Ep7Q�3<��[_q<� �]��lS��c���·	օ$��̓�\@8#�i�s{�c��PA9|������E��Ɍ��g"��}�67v���v��B��6^V�If��L}~hY{���X�=���W�������e[{�ֶ<(d�c�KT)��Cx>:������u�v7)s��v���������{���[���4�o���ݶ���^��jkO_��g/���+��E���-�j�d�,�@4�CT�ݭֶ7��{��a�w���1F��E�w�W�k���������t��a%�ź+Y
gPG:y2L���8K�-;d�U��ΐ�vQjm+�X*�ƙ#�z8s�����@/s:��2��}�}��0��¨9I�r���t�zt�vw|��V�)/e:{YL�쑕�<�<"�"�	��F�q��:i�����}�ұ������U�u8:P�u�2�l�x�*����+[0�p���^�{����i8��5�f���6�g�^iL �x��
�@����s��5tF_�����*���aY��V村t�[C��/G(�T�j��n��К'^�ώf5t���5��˾ջ����Y2�3�E>"}��QM ����w�a�} �Wv �S���9H�;�ЪN���|�d�䚘����v<��B���!1����Rq%�mZi��#5�A�~u��1��Y�rw\�,ic݇��5����Ah�|캠M�j�a��R�,�_)_�og�+�;��~9J�z�)C�����,��`�+̻�P�t�G2ku����J�x���-�P�$9�[�����r}O�mH�ی�����׮+YҊ�edsc������h�$�22ʕ2Y#��(Y�c\1z#�8�g)���H*�Ut��W&�*���A�ǖ��"zp�Y�ZuO'�n@R>?�i,��f�-X�g�D�(
CUR�J��'���Ze-�+�i���t���yj�8�޺�
����F��6<�b�N�Ӓ�x�OK�aP`�hp�@ �Sih�~ޅƅ�Id�T[Y�ɶ ���d��Vn���"ϩ�6{Y��%����s�GX R�Ϝn��{�ζ:��}��e�)�|�������`�zb����#᪝�B���0[	c0�?sX�ҭ�"���9�������S������ҧʧ��� yɓ�����i�Ħ����$q`�3,s���AL`�dK<Y9�{���}M��n�rwZeyέfN�N���*���c>�/@D�ˋ�(��\H�W_.V}�K?���Pqf�#�5�P��A�@(�NZI3h���N3a��n��~u%����X�W���e���m���9���o��Qf�>����22�-Hd�{�yy_R���73�l��{}�^��4Ex��+zna~��i[[{�R��*��&��XW&bџL똜#�7����F��E.����/&��H��(+P��&F�Y�+��n� Yy\hs��`=<u��/�j���o���O�]�����uD�1���|����h�,e�+OK乘�:��v�خ8�������,z�۝[,n��@&���{,�!ii�p*��	œ4��2��Ho���2�C�TWɥu�yp�3p��?�F^����A�^��c;8� =�o�iyt��&Qg�Wp�ǝt�tAe�8���Ol��ob,�8|�u�����&�lи��m��/h�5t�?q䪤������6Q@�M��ǳ��enml�������^a���I[���{�m#�C9|��������/0��=�O<�]˾���nj{��.����N��:�|��z���%�_j�����{\��{�������?�-���	��������٣�����M��~PF��:�,lG�^俍1�	^kk����|�����N��5�j��A�%cۓ~>��3����o1����Ȫw��<��фVK2�KfW��Ӫ���{mә��PR�@��՜@��jZ
��9������n�m~�����w�f �▟}Qonv!��G=�B������`l���*F*Wv|� =qE�­ Qx��O��O4ߟ�����>m���SvN1��Au(��pOzy@�5`T��/�_���t	m��S���$\^�4q0�E����BE�f�c`Չ�t�"1�0���À�ۺ~��t���Z��Vݪ�z#����:��ⱕ�R���T��P3f�,��cx9��%�Lh$2�Bϯ��M0��E�i�ch�:�i��������W�I��sw�R���e����Bz�(O+p�ɳ*v���{�e`r��+i	�nbF%����p%O��WT�z�ؾy����Uqx&OY��W�*��(R�\�%�<+"��ty�Jv�.�j�������o��敤�ͽ׹L=�ן_��Q�v�jdi`��9��Q����� ^�(Әr+�ߡqk����}�E��U$�=�,g[�e=��n帖�;�x�����=C�o2���N�:ҔaUFV��������Gլj�[�����y1&��^���A�ֽ�,��E����d�+Seh�glhk�J��>�K���~P��<q�����΢(磪�>�{�^N��ȗ��t"G#�m|�R�طb4 ҿ��"�+�鯜�0��RΣ�i`5d�S�NeZ������S6�'�T�s".V���l�u�o����Y����p���l�,�o�yz��Ύ���γ�@y�0wܦ��Pb�a`ah�n*�c��n��]jR�;J�<�wYf�Ϩ���ety�Pm���Uo��B���M� �)��:9�)�4�c��]��P&߯����/�Lĕ�p�AB�ۆŧC[Qvq�V�*w��8�����y��<�Qh�=]03�U`���n$�В�T�K�O2X������I �|�G�C��H�Ь���-K������v�s�iP���g�k������aE��i�o��usU���Ac���@���?��={�"�V�o'7 ��9�{^� WWV��͗�=N>�Y%�5W�^%mߢ����l):HC�sϗ/���bdih;f���'��wJ�Q�t;����@���a�jJ#�sx�ʬF�iL��Zp��<���v��[G�.�V@���駟�_��7��%~�O�H�b��ܚ�G���[�[~0�M�f��Ը�LF��|�{}b���_������}�Iy�(G����:��e��W�@9ЏvS/1�ں�=o_?~Ҿ����6x(gkk�<<���1z�q��"�B^�����n�"�#���P&�Tڃ�;(���X޷0\�ڀ>��1��R�v��7186bhh\��W�K3���Pu��C/0l��ϟ�G_��F��]��C�����}J���	��Bɧ���)4�<]���OF����3�ri�h={������Gy����_��_}վ����g�����'O�`�l�=������_a������/
�&w���6\��8X�F�|��r���g�G��5#㬿�8���|����5yyXF� ��wy܃B��3�)��N��Ǘ�!8>�_;����0��)c0>�I��Y�+8�$���7��?�����E�������<���B=s���h�A�Rx.��,�;u� �{����8u�C��n�ziE�alѹ�s�(����N"_2��w?j��?j����2�� 9�ar��������_}�:'z�x�*?�h���o~�v�{�����;��} �͒&��t �+�� ��_��'ړg���'��d��긽ܤc���Ϝ�(k7/����]��-mx��s�F���T�$���N�=Q���?��D�_��;�U�J���Wp~>^�,�e����*��%����w��ʩ|�N���B`������&ϒ+����.�}��3=3��Z�!��HFpI�}]�B�(�r�K�bf Ƶ7��i}>�soU� ��PP!�V�ﺼ�'O�vbr�]�q��\�����Je�|6I��uJ���g�d�?�u����t�@���#Wi0���&w��=hW�f)�{jA�
D�*SB������S�.r�gZ䈧���YYK<�*�j���Ɇ�|�<��O>}@�8|�q�
�%D��Q�1=
�2�����|��v�M�d�F��r���k"I�i]��<$�T$�S�+e����X���JY�A�ɭ��"8�5���u�==�ɵ����}Zg0�sⱻ�"���������v��q��g��$�U*��G�w"'ƶ-���:��b��$������	�c8G��([�s����|%�Z��nm����P��������>������{���mrv:�F����W�o����o8o)�����b
�-[�-�c1�xR<"�T����aq*�́�����Ct���=�rFO���Q�uN���Q���9���)�'����H�6�����)�'���\4�3��ϖL�P�5ͻ��4>T�� -��c�� �l�-�'�����r��N���p8�4�`�E�Qirh����By�}z:6�S�r���cp~���\�^���e����j !��e�`끳�D(3ĵ��ı�b���Y�p{�lLc'q=��1>2�V�wz�V�qE� ���փգ�u��^�T�V�N�#u�\Q7Rv��ڱ�	��f]����@�i#iB[���6H؋�\�n�Aqﻓ+��,u(rg&���H9����Ę���o����`�_�� o��	;0��ג���?I���C����7�K�Q�fu�b�S�Z`���b�8���h������|���?n?��p}	C��m������������h������:#��q�0qm#�@[X�i���i�s�����/�
M\G�~������,��>V!� o�*��wm����14����W_�&f�I����a�:A�-��[�;�78�_�$`�۰<08ڦg���������V�h�㸁���l�[��8��h�!?')���lz��qB��o1��W���o�6K�;����8�;Ҷ����8F�^�WƤ���;s�ͥ ��]��������6��P���A����?|D�|�>��0�v�i핫&���19�J��c��ݣ�2�!�G��W��^� ��mzf�ݹu�ݻ};iC''�g�4���o.��3��こ����lo���r��[h.8a����������mf�r�b�\p��,�0==�F��&OGA�`�6���9��4�+��@r���ה������Pw���oϩ��F��h#��,-��nv.� :@��]wy�g���_|Sn���s�t�-��ӧ�{�݉.>r�1Ґ���S�p	��9��w����{f��ĮS^���A�7W����l8��޵�"'�ui��~M�<\aX�ߞډI����z�[\Pr�l��q��vl���Mb�V����;�2p�1G=E�b:\�u%�ݽޮ�LC/'�6��c_��¹����_�'�:Y8A'#�K"p%�L��d�*��5He��lg�R��C
{�;YЮ�b��8X�Ͷ���ښf�����;?Ӿ�ѣ�G��O>(��!"U��2��Y�S}�Vϑ:�9�r%̾rm����<����W�M��<����s�*�{����8Y�8Y{틯_��gN�t�\�H�Sq!� @�B0L�ܨ�#���3~=b�`�u�Y8r�#�,��3��ݝ����#���:F`c�4<�S��c-��ށ�	�����3�<#��;5����\Gee2�8������ڍ0޵,!;55'��ƙ���F�n ��,*$[�u���odd�tG`<��b�}m=�����W���0��Q�qa�:Ub��r�� �-����#�W����3'K�P��<��sUF�?c���<�(2�yG�Ǡ��9N�O'kp��#�����,�Eɧ�8[��9�<�[/�C�l�%'K�q#-���|�Y�@Y���}�)�����d�-�NV�{���֕q�!�K������߇yv���o�i�qM��ut�H3\�rs�����=h���uȹ}�������[�N�@�?'b�Jl����cmo����mm����!���$]'��e�jy���A{�����{��Lۛ�q���O����?G٢��w���k4��Ttq�'F�J�guX�1��[�Q>FIt��ޞs�(����^Cl����'&|�þQ�!��b�dP�M/Tp����0����x���8<�c>qH�����i�FeG��2�����{p #X�'�@2�͏vpcqG殮eOш�O``ML8C������pSF�i  M���9x����
���{����5ؠ���]�4 0@Ͽ� ��ת`�]�~.O1�ң��@�����.�|{�ytt�u�uTx���C�R���A�3Rg9��إ�÷~�p���h��E��J��W��(fda�	W�`�h���E|B�:�ټ�{����Y� 'O�{�Q����?ӋQE8Bv��Y�Y#Y��Q�k�DZ�qJ��ot�\@�y{Rt�18�/�GF�b�=��ꘙOR啶���^0�dsh`�J#�q�Ґ�����r����d��vmq����V����q��o<��f�&"�_<������������V��|��ظ� �[��ݡ��w�,�޻��Y�0+{����������O���8.n9��&�Y�Af������m{��k��𜲌*��[��ҧ�1|��w�^�@=���z���
:oj�s������q�B瞒��"w�ݸy��'?���j��2�1�M��o�n�ӿi?������]r����>\�#E=@:���j���M�)�1�w�ٛ���u|������(���`��э�������}��G�����/�ۯ�����'\��>�S��[�� 7����V��✼M��<:3��q�][Zj�q��o<�B�]�����������.%�k�h���PV�������D>n{�����-�._q18���^wO�}�Xϐ<7$��3/]WC��f��|�d�ԫ�ˏq���	W�8W.CF�yV����޿�>��i:3�����4#?t��󟷿�[7��<N���\,��I������K�/��Eg/�:M^�PN�waV��	>B���͢ރYL<\�Eo�?(k`h����\C��um���"N�8s/XuU�z6��P�6�0e�b0�ۭ���~���vB{6���a�O.?�\�\e�=��m���a{���67M���Q��m'���}����w�v�`n�KJ��Q��dM�ɞ9Yٌ�<���-?�X� H8:�^�BQ|*K������?��&v~�~��?������M�]i0�-�
0��s��n<����{=�h��2��Wbv�� �*Xӓ�8�p�����q��;P=Y/�ڗq�^��d�S9(�#e6p(<t �xF�&�}	o~�0d�,��d�3?������t���EN�ȕ��B�&�4��A:�¡�����W���=q���0A,�iA�2 L-����� p:��c�m��r�N�u����G��8m�E������HG'k|
�P���ٯNo�^m�o��9v#ص��-���
��R N�i�U���)|�o�ĳ-s��C<��|��J�Ж�Q��B@P�@�p_���Rm|���i��g���Q��a[8��B��(e
ᜒ��3+��dIU��pVu���H>�tG^���wY͓��7�%J��(���tu�M���&w�+��>�\F�q� �˅Oœ�<̰�z_1������t��\G��|�*x�����⽫�UoF?�
�����:Fж�<���~�=����8Z�he�b��+�j�[f��� �Qr^��w��<j��A�q�&2f4C����p��&N���Ri+ƚ(�� �K���S��?ꑐ%���xѰ8�8����3�֖��c��ڊR�t7�\��g��"n-�3�q�����T*b�����3��Tr��:������G��3�N��{p����(~h�ol@��������V�P8���XMN���)��Jb1�����5�+[�k�ۋ��0{�&���	��S]AMCB}�#'��,5����&��C��b���������p8wr4���2��Ic&oU���8<
����=���{��1��"ZV>��I>:���.��4�*N��NV&�G��0�(���#9� .iV�SQXn��E?Wީ�KF�ݲg���ʽOM�Z;��q����dx$�#�P���CʐS�%����������虗�$M	#e�D|�|Vo��(]8�Jua����*-W��'���������h���az�>���v��|B��춯�~�����?�������/��)V�H�c�ZZ�d٨0ɳ���G��7nf��7���>���?���#3��i�)e6���7_�^<��9/�aX�SY�<�; \%�ذ`W|�j�=��z�֞x�75�@|���3'kkk?���ҵv���v����dde@�c̹Z�Y��D;���g���E��W��z[�^�.�SmB��r�JȐJ�y���E���Ξ,�DC���yl�v������滷�ڿ�矶��~��p�MNPV����F��?�U�������~�� �=��n��%�l���}�R{j��8���t��P�"�(;��}7��M�u$4�	�l�~�@W������*6�x�a�yqS��H:�_��Ŕ&'&#w�}�~:���.~q�W��\���iE�eO���f�pnё�;�c{
uP��t�n޸�c���'���8�Kmj�����`w/=u?���i?���h?�Yv���"�o���jcaec57E�Z.�|Ak�q�a�<�0F���py���N֦Q@��3�<ӝ~C��]���!6��B5��������ɆC�q�6�N���d:�pv��+��Uy�\�F[�EY��Q�,��r�ƅ?x�~������]_�v _����?�?��Z7'�������5'K(aJa�O��B)՘F	ϖ��9~�����t>PV�:v�
��(�.�N���+�!�[=0]	^B�-��3�6?��	��)���"���[�.i�'�/�5:��7�<���"<L��.BǱ�'�&|N�<�Ċ�G��S��%�~�z�1S<�_$ ��)�Ř��}�S��V�^Ǳ���:>�]=o��mp��?�h
�`��E�Q%
^e����,�@q������}�d,B�W�=H<���q���{�;C=)(F���$�$tq6� �e/�ll�Pa6�J�Q�� �~ΰX�*c�F�+*�R�u6nzay�i{ NW_�b<1�ޖ\��~�庫����˓��$_����'N�<�^zVT�"���܁X3��?�U�ϟg���A�_+�����ﻣˣs���J��(��y�Z�����������r�z��
�*��}[�<+Tm�͞:	�� �����Q������/{�lI^XZlˋi9Ԩ^}�=��qƀ�~�*=�\�!֤9�/
���6�|(��˵��˙�r��S�B��"W���t�<�ե�7?L�K<�K�U���Dy�AFQ��إQE�}V����$R���IY\���g�fØ=�e`#��et�s��ɝh+�����B��2��L��+3(��vmi�-�9�92�R�Isx:�`'��}�����;��cmgs�e�h�3Y�xv��Ϲ7�"z�z�u�v���}��v�����oc�j׮�i赶�`#�"2o�MO�e|�	t1��e�������U�:F��X�\�n�TcWy's��0��G�1���	e�s�������J�����qPuDH����;�i���~rx�,���ב��:�:��h�k$0���1���K;�6��m;����|G��?��E�h'��xeE9���t��������=Y?�b�Ƈ@h^���t��\��]D�,Q�B��_^�\�j�h�.��d��{������N>_eH��?��s���2<����:�����
�!M�@���΃����*o�C�����
��h"piNU8����U����k������^�i�+�bئ`�F����:o�7�~��mx����q>�7�u�wW�s��ܜ�b�b#`lj`��p5&����q&\��sg0�&K���6$���k���*W��zL���:1�8������0_"����{8K�N�=:�j}��uO��j�������۾y���v�M��od>՛�7���=�<|ߵ]������gCg��C�^���7o7�Χ=��w���"6����m�f���]��/�5�m�g����^�����8L�V��4������Z���L�dٹZ|������
�{�s���k`� }{�Ź��v���A�Yl<Z\Z�i��f����Ed��O�r�ɗϟ�'�|�^<Ҷ�7�t�U'~ow�l����Q; $�&|� �3��Q"�W�٠��͹����QD���.�N��|M�Q����A'�.��m�J~��a#,!���mW=4_�����߽0�cG;Z��w�qK�r��ؠnt$�#��'�>�eo���R���rh&��y���������x���됄C��=��{����:���~`:Yah�w���_�E�ô5���d!K%�A�d7�_C�,�� �h��u\��2j�~'"��Z��J"Ɍ���OG���F	� nVoA��4�U_lo�`m�d9	� �ٻw'׃�Q(C� ��#��*ϓ�?������ۊ�Pyy��g\��ɟ���"O|����S6�G#��{�(l��}���bo���&EvA�!8�!���@��Y*5c�1��PJ�Ơ��uZ�/�Ղzٯ�����@Vp�%ak���a'xdd,-���H�-B��qH7��&s��8[�TL)�h��21��Q���g�{�r�s�LLq�J�Vl'�,��ƴ�I;x��*�5J`n?�+�)Cン¿�S�q4F�z:�vn���@�t.��������O^^ֻ����S�..��U��l8+÷�:���7�>���� �y\L���{��C������=��Ѝ,�:M\h��}�G��sV#EN�*hu����_��Kep_�ޮ߼�V�]K�-{�;��ɴ���-�'��K�Ka<$?�GbP���Fe���$%V�y�8��}[��U��P+�V�6J�&���~wM�>�wi�z;8Yi54�3���dKrB9Zg����*��y/�H���+K\,��.�����!�i��r/"�C,�{���]������v{y�-�M�鉫m���O�Ƚ�=�8{*�6�!���C����S{;�'m��lc�lm���m๊��Ӷr�ݿ��=|�^{��G�N��Ç8Ww��;����mi�z[\�ޖ8Z++7r����#~�y,s�nT2�z��404$�á���zD�%u8� 4�E�P�����`�H�]Fl�ɾs,\�@�Օq�\��!��tZ��kX�=�����e�h����=V{'ߨ3e��6H��d����+:��I\��w8U����J���\�չ	!��&��4)�h�'����t/�˻1�H/4&?o�h���i������>߄�5��y��v:P[B'�t��S4�v%�y��꽻nںB��Ȯ��p�/������_�M�����Xg::X�|`�����ެ9��,��jn�oC�<��a�6`j��lݯ��7�4�_b�on���=W��Z��tƽ���Pp����k8
�;�g#v��Rx[�w��\��Kt�\hn~�McL�k"=���h��S�c�k8��'r��C౾��e�C�L'��pjo���66�/r�:��G0s��wdO��27Vڇ���8��6nX�=l�W��ص���'ϲ��p�Se����^��u�����X����T�q͑���,�A���mWG�'SG?� ���	B�x6_{��?��q�[���G�R��}��w�����5����lϷ=�5�&24���ƹŠ�LN��_��V�������N��~cw���OC{v��\}�]m�������G�ț�8�Q/�.qޫ���S���xг�6��m5���5R�R>����<O>����P�Wڲ~�q�T�t ًe�-i��@�#0��ё���x8ψ���P��v:8tsd�.]�����n(4�۹���[�ndsf��r{U:'k�=�ɲ7˞�C�}�+'��+�hq�(D�;�����D���`�0�j�TP�2Q�� �~#�x7Es��e���L�Ҍ 2��m�#-$=r���qb�hA�yC�5��y����'
b}�~uA�����*'kG'�͉�G��E�T����ͅGwM�T��e��/A������sQÎ��`�<+�����wz�t�\�"=X�4��b�''���:�t���(�H\!R*Ϝ:�`2.�����4��R�����XN8�����:Cx��B�*\e��ѱ8��5�����^�/�YX����1^��)�%��ɬ�TB/F4���9����cXI,&����r�U94>�@V��:zM>�T2�J)�JB]]t0HSүx�U#y�БXrKK3\R$f��{�ٲ�g�?��^,�	��E��}���g�_� �֥W��k/�t~�x}�Y5g��=ēG��Y��!B���Ht^b�P��4xXO��H�a-"x�/f��˶b�S�(��P�^kP9,�a<�n9��fz���˗/��o�nO?�p��Q����k���=�!�����>���4�J�T,��A�Jwεf�1�}�ݟ�Y<&��!�4�#����K��Js?��s|Ky2|��������A�X�(��z"�Im�3!�y����'�k���|��G��D\m�c������{w�G�n���^k�V����X�vIu�=o6,��Tm���նM�ùrY~[OmhC֨,���v[d]�D�NLN wn��}��Lݽw?�,.�����6=��F'����D������Dg�(�e��qRGR��Ju�M�ε�)[�1�4:��5���ب��0+(Z�'oK���3���1<��+�<9�q�&G��Y�Ź�47���Н�ae����.�x�@&O���i�'�M"��+�9�(o�S�(�#�Yp8�6�\����O%��M�҄v�!�Y��$��/ݐ���y:#��a��˵�+=��ޔ�9�3��4��"�Lױ�a���cהּ`>.x�w���6��ݟp;[�rc�充v�6r#j'7=�Ώ��j�������ز0Mt�zM>�0�0�w����4�B8Y��A.��_X̰A��ɧu�3r�`ғ��=�d��bO֎C�o�_�	�2���z����&�.\��m����c�|%=3��� _.��X�b9T��E�kǟi�����zY�$�:��h٫����"R����Վ̜`�����Α��F3<zpuc�ٵ �o�p͛7�ڏ>��}�ɇ�.���|*�@�K��<����ڋ����؎:&Ҧp[?��"W.�e�ݻ�~	Ms�n�����L/��y�)5�NX$��ï3�2dA�S�"+;�K��!A:)�@Ɠ��l��q���.�SKG�z	�����Ao;U!���8I�Ȗ'l�F�r+���:�nݼ��g���|��b*O��/�y��?kO�ykk�q�|��Ae�|�5v������wy��Ym-�˱�ftA�8T�����u�q+;\D���3�ʓj|��
&��!��L��i��HF~vt\�%�"��2TçrE�+*�#/�G*Bꁐ�R<��ccmaхa����<N�C��#�����h��mS���j�	s"O�)$�ǩ������I\Q�J�T�
�{��G|�O&s_�tT�qU'�9�p!��"Ac]"�	L�5��V].�e�q|�2���l9�����kA��$*,���l�P0N�Ȗ=Y�G��p���wK�*G��b��-�g��J�氼�.'�z����K���g��`m�����{E��]N+��|ch�{��*��u�|~z�p�n��Ǣ�.����!�rH�^��C.�:��m9�w������ü�ji � ��$U7�S�f�	��2D�(�t�m�v���{[ܼ�Ԗ�lͫ�
l��C&��K�X6���3�'��S@��}�c�� #"�c�j�ы��CA��0��WpO��gzI(s�
�R���ą�9U�u�;n��#� �[����㵾U�T�������ۡ`�^�8�%4\we�I�{^�����������U���8�^�Xz+�I8��RW]}Ep*�l�R!;�UC�Q>8<,� �ҀC������[*s�	޾u;��W������LNPw������oå_#�#��U�yX�}�@z �4H]��@�2&�o2OPc�2dO�ʻ�
�>��;���:q�&����*}����1L���I�O뷊)�`�B�!a�P�>����̧"�U����+:;�v�F������� N^�w�ߩv��\�w{�}��N֭v��B��B���e�A��P�l�űZk���o�d��C �|\X$<|Jn���x��:��y�ޣ����>��G��?hר��%�K�a��5��ln��R�qN�΄��(�{�fgk�����8[��1J9�qoG�'�����u�|�R�Y�(�;��5{�t�\�W'kzl�-�L���6�|D�`C��T�U�r�C���w������Lt���?S:RQ���2C	6�b��ꤜ�!��ٚ���\�ȯ���~�K�Z�$��	�G�$PV�>qt�-��ҟ���)������F��-���r�	li_��Up�0��^��5���q���[�H:1B#���-��,.�035�n �-/d�~���t�mo�/�x�!��o7c�
��:.~��z���O�3��37S=YYY�L�wj�~>�_��r��ǯ�q1��M{���(�j<]�SG��O�g�r(�K�;���N��� ���Dh�9C�=r�p"��ǡ���ٌZ�^3�z�6�w�YG̡��P�e�[k���E^l��p~���(��g���o���t4^{{N����Փ<3=��?���޿��l̉:'m��ry�g�^6�ط��ޢ���^��{;��UW��{�ĝ4���>p�%���\eoF�؈�A�����'��8�6T��C�q2�:O/e�y���9[�} �Y'Ȗqd��!�jG�ԩ8$��,?��x'�\��F�?�+�~������zv<mei�ݿ{3K�� �V�p�~��/�g��Y��~���8C�0ih��D%=e,�}l6�_�m���$�~��\}���E։�.|[Κ��������~�_w������x���,s��du�q�&�4��J36��Z7��֔����LVj\Y�o���Ԁs��W�ŷVn������b<����=�.��9�Ȍ�Fq����3�/��b��\V���:4B�����/����������������_k����c��1�	ypwk��WF��+pzm�[����n�;wG������q�E�d]��ٹ֜�g(�"Ub,:����~�`�2���<����©�=��X�M��k4u��N��M��ۏ��1��+W"h8��Y�	d&H�J�N�S�u�"xG��|�^�t�us�ݺ5��5���_j<��>��N{���v㺛 ������Ժ���.FR1r�7ݰ�浆���BP�* �k�%亞Wʭ�Q�a6����q��9�J�,xv���`e_e\���I����2���/��3?y��b¢_���i��	yޅG���烜����G,��9��_�u�^���a菳|��'�/��S�s��I�\
R#�F �iP���w<�*=���d��<㊙�ܬ߻*�K᪔�3%���J��a0� }�|3�8�� ��G������/l�H��T���OZ�Ut�w5T[��<]�)Wʚ��4?��>D�;���
-���!Z��A�А�j
����	��y�'��\%�ߥ�x��t�$�ڥ�-x��-���wf�'�l������O�j=���^h�0����pbW���_�h�8V�[�	{�n)�_¯�n�K�S�vx����v�.�jw���L�u�^{����O1�~��v���m�ڭ6�գ��Tc�T��4D�9�y��r}t	����� ]D8D�h�r>vq��g�3m`|��L�����{m��n�_�զ����<��x���ӉӠ�aS��Ni�J��z \ ����!��(���aG��S�S8�s��E��
��M�E����27�v�M�Y�Q�~.�쁷�s���w����B��pΊ��.���C�:[���p*yCE���K�y��{��cp��2�N�L����a���=�����ư�Qq��<!�J��ҶF�N�˔�]�Ј�`o���o��E8}�/P��p6h�V�Od
�	��憱n�����t�x˻�E=B3�Cna=h�u�:�*�脘n�@�/�+~6�#A܈��n �3��^xX^�O이�:=�Jy����\j�䈰��9:)���q�~_���	 �8َ xw����Fv��2mD�D���`!����@�ƿ�S�.����IZס;Д<���8&��q�������7����`{�z���h�tl�uێu��=W�ù����3�h�R!3�c�u_.m�Ap��v�eh�������]ay�e��>!L�F��xgfp��A��
��Ӯ|���Ny�1�r����i���QH�Y�A|� �#ec 6�{����	�9�`���q_w�?b=h�Q��@W置L���T�Q����ӧ���?o���/��8Z�A�0y7�u踎�� �#���,8F�ؘ�Y���yV�X��	��ɒ8S	�ql����7��4�9PI[}k�4�(M^�m�TDZ�m����?�<��o��%�o�F�f�1{;�����/+Ǌn�����_���ye��}�	G]C+\�=�?�ߎ5�1^����:�O8.�s�vV�xWw�����f �1�hW��ﹾ���e���k���?��������~򓟴���n��^�|�K<5�o)����j=�:��F�x��/AY���r�=�x��w�.ƻ��µ���P9t�P=
�~�C��+C"�,�d5&e���CB'�a蒧�׷ziHI2�!��QQ)�4�l�C�v��
�ڽf��`�c���շJ�k˔{m�!��#mv�ea�������e�5�����8ݖ�p������h�heȢ¯Zi�^.�_�L�7
�<��N8�&|�3��N�u�w���d.��^L8X���װ�����1*�R_�\��ϩ�~�������>vl������
y�?�T���^�'��z������Ͼ�δ�p��O����7�o��S�z�鲗?��Z�I��������ǜ������_�.�!W��$>�^v�#���o��W"|�둖d�٢�+�TW�QNF�;����1��m��W�G�k�0^Z_;T���/��L��ҟ�w�޺��}X2�<Ja�'¹�(�bf�Ζq�H�a}Y�:�Ş�Cx�a��9$p��,��w���n�~r���{wۣ�7��[�my|���f�^{�V��^>�M{�����+�Mx�S�>�����%F c�y ������T���^�������`�{���p�Z� ,${�lt�|�#q��ĵ����N|��ᘸ�Д�
����ӫ���\�Yi3�7����@�[��fV�g��Թ�v;�b���t�V�h�l�`��'�{]�������#W� ��aP��t���m���񦐕�Sc��<N���	��8=��u<_��:mW1qz\'��+�?|7齊é��Js�8[q��&d(Ut�	�+u���C8ݧ��C��;�'N�p��a��θ�H!q�E=���i�}���le���|���Vz,>֊��5"����~%Ct!C�x�c�'�F#�FCyS��0R뀇�ӽ=1ܷ���Ͷ�~�]Ҹ?"�}��ԩ��r@��urD����<�{���~u�4����SAy'[�P��G���O���\�NY�&otVS�����&�اib3�"��MaPFT�:��m/�1��`mC{n�*<6P�0:,�o�E�b#��d�ud���d�"���Fdt�<m)�*8�[P��b�)+6��O���I��o�Z�u{M]������Ջ�m��z;98��5��G����A��82���/��O'/U������h`����@�`��P�c׌����v��J�|���Y�𽇷۽;72�t	g����a9�=��8Y8��Qn1t��_��ҿ�8���W|�?��}}J�.04
�ad�8W���u$��ˎ���rA�o���u��/~�>��g��~�޼|��n�:�h N�+��:u}��A��*��`���8Th����;Ñ��C<��*�����^�E㹟�S���3�� �AF���0� �c{�w�; ?�f��A\��Yއ�-�zS'Q�v��}�fH�r�N6���b��r��Z�C�A�᧰,��D�n����]<3�B����>�ޘN�w�R����ef�����onl�a�K��u�ٵ����N��@ n��pA�F|�5�n����
.��	s`��+�y.x�g�eltϿ{P�z���d]���{���:��G��_�P)se3�J�����(X��(��
:�Koq�$��8O<���Q1�@E��p�_�����~��J���"���zg�b�+�ҥl�^�H�(5�c�������/.��lͷ�7܋Ca4��5���ϮW�gs)�ѮW+�Ӟ����W(�B�"φ8P�j8
5��ǳl
_Yn���U�z��n8����ǸԈ��e$$L�|%��F/�����q��]<�J��.�.!�\ϻ{�OZ�^8]ȟ玟��kB�����}F�y�\��?�����\W�>J�h�T�>�L��W�E`��_[UU�:@�Wc���Tg��y@:d.��~\nĩA��b���әܤr��~�=�V_�O}Q+/�e��a�w�����|������R��\������	|���k���'�;(Wnr�r�g+�Z�i�Ø�UϞ..�8��e�����ɡvmy����F����k?��C��{܍c���2=��5��>�m{[o���m��7m�Փ���%��z;�w��Bp�Q�0H���NQ)G� #��s<;?�n�Ñ������{�k3��o�H�(������p�!��3��ժn@���n���︡�4�����6�C5����Wn��k����;mq�f��m�p���P�f�x�s��g�}��\��o�b(�#/g�e�G�c�`p�@_�Xq�����05�n.͵;�2���R- 2�p䰫`^uT ��=�4�3�,g�z8ԩ���N�O#doGc�:p1�}@v������d�f(�,s��˟�i�.A~� /H��ق���:j8\��q�}�"h0�%��S<sDC|{V0V�0N�P���jq���Ս�����_}��������g?�U��/ݾ��I[_ߊ������C � ���L�zs��z��}�v����/N��#�:��׹t��:[G��*���q��.��I^�m1����@�6���yK4q�]����u�dRn����M��w���D���o̞�Џ��q'&���Ts�{�Ж΁���$��w�Q�$C��o�jV"Hk6�f�ׯ��Ʋ��C�o���s4Nm�B>��	FT�/u�C�m�v��+}.�S���ġ��>��>N������?��'�_��?n���ÿh�ۿ�������O~�~����������xDf�1H��S��ɼ�7�;�Ydj
�2���7%�9�򧒌�\ N�/yH:�}�U��'�㶽��^<{޾�������������g?�|��ϟ�m_D��������.�G��=^{�]���*��d��zt��2dYe�,�E�̗{�ѹ�3���{֤�؟���8Z��r>�!i����f7�ׇ|sH<������JY�w�R��|�J�6`����8��F��aM��FĎ�{�����?w.�K]>quA��@��	�X�R�4H�ʗ�!z[�v�r&����J�z`m���M���F0R&�g"i߮�57]��ti��1`F���o�_���_~�^�������=�n�-�+ח۝{wڽ���4F�-]�� �\ڧv��N��rŃ���Kmc�n���mc��HZ�=��+C(<��Av�V�VX=dfҞM?wF�kٴ���9�u8��k���C�\�"�/k� ��-	�T��R��T�[f�]:�!���˚^����@�1�g'�]��`"g�_i�P�j����8��Xc#��!�>=1�������)� ���-v�CX�
,2�"� ���-�&��c�k��mjjŀq=����N`��=�	c_�GM�t���m����/	T�5� j˯-d�|���6[qm=(��(9L��4cd�4^C ���ܓ@
��7�!0�`�k>T�����m~\�Y���)h��\�`'�F�-M�#<)ۜ��?�r�=p����@Y����;S9
��=	��>|�^ةSpח�wT�3�2~]�a9}0K_�|�0����;L�o���ַ��`�%��i�$���V8��3ot�M���,��p�t���]	Oa��X���.k;�}_�c:���n����M%m˞U�.�X����w�C��p[�y�`�>N[��z�H�|!���_�p�ϱ�D�`>0��3� N��
��u��������Ud�Y���<
ZMu�ex	�}��`��2<�3�>?�X�;�8�
��O|�q۠|k���F��dȯs/��������ۣ�����x���m�jo_=nۯ~�6_}�6�|Ӷ�>���v���?��#��	n#��mX��2���U�7<wby�9�݃d�v�anf�=|�}��?h����j�ݣ��1�������$�8���'�O�ԯ�䝘��'�|��ɋ���6h��X�>�uex��C�na|�r��ƛv��3WJ��Q�8����Rp��pe%<�!���e�T����D$F����la���St�%p8D�c����@�q͌��QTe����8D�Y�~�����3~��ʐj��C]˄�^:Aߧ�� N����*�i��b�<�!F�4(��O��[��EW�O���v!�g�2�4j���r��aO��_j�gu7�Kп��:�n�O	����\�A�@Hy�k#w}'ok� #�q�ca�D�_�����h��<�ۍ������Ͽh?��g���|�V߮Ʃ��Ё\���.sԅ��I�c�Ч۝�������sLnI31�3�[�X�,/�	�t:���u)�u[xx�s�Umt����	��<<p�<W�;l�������|�>ש�S��qN�N�$�CW6�f���0N��!h�$�!���=�3��mzn�:�����/�o���ac��]�m��po7�r����,���hGhkK��;��ҁ��3d)�f���w���ڄ��C����n�%���VۗO��ǯ^�5�����lQ���ҁ�m�O#FF0��(��g�!$)��> 7��48xp�>�{�>v�kK8\��_~�������p����޿��޹ٖ�\Ƕ}�r�mn촫ɸ4M���-s�oh�*ϑ룃��72� }F�eCa�=��h�Xڤ< g�S^�Gg:�Y�w.!S.#+��\9�BC��������W����}������*�[:)�H�qִm8gG��u>�������{���0X��I#�-A笝���<�gJ�����l�x�w檱��6���<��ô�U���D"�lB�'Q���'�m�G�kfXΠ�B��G�m|���,����R���@������ß�m�d��.xD��d�`�2x�I$�p9tʉ��C���FDU+�� !�������a�繶l�1�."ɖ%+n{{�=y����ן���_�t�-�s��q�+���-̷��=h���G(һmM+� 2�^"����3��? f���mmk��O�Vt�v�L�9���ā�VJwT����=.��:ξ�Gb��
�����5�#��UdJ��k�"x�U�!$�<��hlJhԖ�/��=�Y��y�sI��A�
j���K�ڪ��X�*��:F<�d����p��c(ں�`��/ce!X[�4hN�uú���Ult�q�_(��
�9F�d�_������õ�N��T8�ZfU���OL=�H���#F�o��G�4 �����}/@���M1�l�!�h_^���W�0]��H"��#!N�q�Ϫ������ག�;�����8I��8�}�Ξ{���"�q}�������x^���k#��ż�2KȽɝ��Fҩ_&J�q�<:b�C��uZ��9O��[8� ఑ݝm�p9#�hH=�
ij���O*
A���9Y�#1�FfI۶r��� @��Z*7gtH����t��b�:5�� ��l�c�?[�t�z'*��NR��V�T�i�g(��Ƿ������ ��Vy���Y����mq����[�1]y��"1D�K�G��E7t�s�V�	�8/�d�}�f']%p�}��^���w��A��������1���A����,�7�x����`���GǴ��`v<�g+�~; "�f����[w�}����fA
<��}ėqC9+�_���������#v��?�y�!ŇF�J;)�~��zA:�`;��)D����z �y�β���ƃ^)��G�Q/�˱��-��Щ�5o� ]d�M�/ƒ�׵�'؋�q\�'�e���P�'e&��S^�����3Ϥk�[��}���r\�,�'�*�O��JW�����l�"��l&1x��s �#xء~#͹mZ�Mr��]�B��s[�"���(��3-^��ao��B��X�a��\��
	E���ng�t�N��ql�׮6��N&Ω3��k�!Cځš^�7�ڠ9�S�g�zuj8�r��Aʎ,�ŷ�Y'�N��@N�6���@�m!�leW�W���6�omi?)q&��[۵W���&��1�S�8{�����%��� z��Ü"8l\��ͶG�V�PWq���S�/۳/ó��^��llp/)�Cg7�Pv���FV��ƪQ���-xf�����XC��k���r�um�M�K�`d�����I[]�jO�k��|���n���mg���:���pb��X��b�i�B:�ewgx/��ىؚ?���S�v޻Ӗq��y�0�n޼�n\_i��Smzf"�%�`=51�;�R��L�M���^��vx[> H��ӎy���!P��Td	���3�u��V@�Ï�SLW���+��9F��Ӯesz������)4���}���`[B��V���$�%�����in��{�'6"����N��盺���r���8��ɻbՑw�Q�UT��.e�0�<�G�O:.�پ�r��Iʁ�%�g�iOփc��67���m~ngB?^p��7#>Dp���Qh�܄AAak��֡%�
�v��:Q�Z dI u\�-TV�ޤ^(�{��)�C ƈ��i{����o�o���=}�mmnS�&ˤ5gjf�ݽ�}��G�����QE���C�H�>Ғ�X�n$'�'� �v�(�ݙ������N\<�{�1�s����|��AB�Ȫ8~������Q�vM�fȚ��`�*�^:[M��QZn�:
��9W^�祁l*_T�pl�à\QP'+X�/�,1��֕s$d�t	��(x�ɪnS��1�{ibbl"N�c��m��hڥ��٫Ɏn
缳L���2dR�w��d�@��o�5�j����]ŇI���2��x�$�O\q�m&���,5�/<R�O�-t��8k[�9?r���\���ԙ�#���B�1�
�\u���ĵýL��\�?�y���9"L����Ͽ�#e�����o����i<��I���#�,�[�Y����j�J�R��#R�7iL�A��c	��[{k�G�a���fm�ʂ\��B>��@'Ǘ�=m;�g�P6�|�6�ꡱ����-�QX���;i52��Ѐ�ՙ�EP������d�e�W�U���,�q�A\a��4��S��e�_娆��{��g�+�֋���P𲱮�'��+>+�K���
���675��\_j�cx|�ރv����47�Ɔ0~�6�ƛm�����B?�hQ�٪ZN��h'�s��\["��2��Q��PPg��y�Ɠ���L�̶k�o��w�;���eP�A�}a�e�E;�<9s�ȏ$p�γx7��đRNk�/B���ĥH�	% ��Τ��C���:W;���;�w
�9�hvH��B��U��ּ�G��Й�_��c�%F����2�op��!Q��p�+{O��9l4����n1=e�嗾�t"�ĝ|T�(�$�i#��N�Ys���F�O��u-�H����hlg¼xla�����q����5I���m��n�ob�y��I��|�=���g����|��?��e�	 ��6\���*r`-rA��HÔl��Q~�����=�D��$��/���lS��Y��at�wa�
�x�Z�W��@9'�׻��P,���̜,�C����6N�2�!}򖋰��6��jo�.�U�.�(��e�c��1Q.���v7���iV|��i{��	�r��(;���r8��L��e��j/�tu"�'s٨Ӧ#;@ҹ=N6�N���-��ח�H�بii��,a�mn�da�>}�ެn���ضҢN�����_��Y�f����,@O�m������?����~�>��Q[���o�S8U��9�.��xPN�Ώ�>���Ȭ�;�@ڡ���MG��e��޴�3����R%�E��g���x��_3y�U�t���W�#O(�E���-x��kk�s_�����������4K\eqx@:���м3TO{&oM�4N���߻�Է��u���)�+��Y�^���I�;��79*N}w1�dɏD�`
X��+�1W��?_��N�N�X/y nt��j��kg��x�\Y^���ٻ� �����:YT�i	:Q��Cf�pF8)�]࠘TemeS�P'�/DLp7x��W0��c#mY9�'�k�hm���W�Z��y{��e[_�cIt��GMʹ;�G~�����l���G��c�Ax��S�����ow����w	!q�OV9Y�d�ӓ����|UO�G���:K}�{�X�9r�j$+T�1�&}`HW&�!���x<�\;�C����9Y2K�R��/~e�)��R�N����|'ю�߾ե�/G�[�\9Y�:�R&8Rw�o�j}����[珡������h9s's���ug���8�k/4���P�w�eW�; �����OV-�  _1(b��c+�e҈�0$`l���NA6	X���g�J��T�P5�c2���[��dI�(	�v"��Yգ%����)��;y��o����?
�ЇpI�yv��C�]"��}"u�]�n��J����:u�]���G���@;��w����q�Ԡ���W���J�[�՛�w�+�� v�p��j 2�B���Ri8/І �� �<ʭq��W�Ώ�rMDW�L��
�����������8Y�"X�l��1J�,k�����Z�ԡ��[�#�D���Y�M��$J��z&/�Z�9y�N�s��7SO>�ly�ҖW��D�^5(��U
�w���w*h���!{�&�1tf���+�;7�=7�\�o3cC�2J|o�m[{����~�v7V����rB=�.yg(cǓ)�q��(�֕#����,���:._��nܺ����[���$eq���q�a�r��C�\��y�B���g���[d^�X�s���ީ��3	Ĳn�ho��s������u����~�^�GZ.�Y�JC8�8����q�����\��w�RWD~��s���8�ܺ��;�Jǵ�'$ǻ�	�%�"I݈�'�I\YW�0�R,�20_����\�c|�̣j�ɒ7�/�I��W-���OU�	�P��o�&�S�r�0ab�L-�T=�~_�4�-K���K�KcA�pE6��e��j�:�N�{f�����(�1(=;=Y����qكj�����W�g�^*�ʽ�4{��_kb��-?8�g,�<���\�@k��}�2��v`���ޅ\�ݡs��J.N���3'k(��J:y[�M�)�8��>z��"6�]2]������
�P*@��ց�կ��H���ǖ`U���!�9Ls�S�1T�������٫���������S��S{�z��Y�!���2e�	|��3������Ǐڧ8Y|�~[�>�0I�A�	��!xV�N[iO�G�>�̀�8H��g{g�z$G����(�\�륓���?|��
"�]�;�]� �9��:�[�m��'����F2������6��F}y��ᮃ��� ��xm��L{���)���KG�H�)�E���`�J�����o��)G���+D�R�J��R��7
�����c��@�aC���8L����1����l�0ӆ����3\�9Y����SsV���
~�<(:���;u��������`=C4v7kԋu�]ضX8�YS���wp��Cql!�UC����ٹv�:J�ރ��'��=lKK��"ӂ�1�2�0	
�V\�qD2��Y�'K'kO'k紽�8J���6e��B
��UA�DLX)����GOTƖ�e��\Y���̘��}�Ye�3����dG��q6]R<+�y�����Ӑ�.�F���54Ľ��`�9@��z���)qχ)���L6��Fp)����:�?`�Z�P�T-f	�q�#�N#(��~��"�Q'�7!����*	ǋ�xIZ�\�a������jG���4���(O[ �!5�3� ūM6mvH��a��*�ac+�b�Q���	��+�ِzQ�.U6
����N@�������N��K��/G�U�mz�=E��wם�����F��w���w����y�%٥i��z8�gH���壳��G`�Ρ0����q�|�+a9;��U�~.��)_ۓn^i��l� ��
��ނ���Xv��ɿ����� |�+i7N�=�8X���k���z�͛��s��m�Ei��{���
�55�x!����}x�k��2I���z.n����)y�+�
}l��FY�6���P|L�*��B�d<���W40:�\�R�!�O������߿�>~x�ݿ���'Gp0
���������'mc�y;��n�����`�v_'�MK/�'#��l�"�(f�C��Z�NL���%����v��{m���6;�Ԇ&�S��)��%� �x���C�絵H�.�O]u�Px�d�g�+�k���WŃ��Ş�7�U��X׹�r̼����G޹G�c����.�H&z��U������<g*CgdeH�F��,:�<Cϕ���[����p^����(5�\T�.�4�X6�	�UK/y��<�7p����!��C�<����?����R{�|�9���	��� k�1X�ieS�dU�/:���tH'��	��z�����Q�p�:���J)�
��Ti	+��
-�;� �@~J�߫��(e�.�zN:��;�Y8��Q"3Eƙ�!g�j~n>��9T0��u�a�P�u��'(�=W�λ�G�p�d۱5�HY3�̡z�mr�İ�h׾�v��.��� �AtN�+���i�����lcc]O����q�[�mݽ����kcS�k;=(�M�Ʌ^�g�z�t��7��!�%�t��&�6��T�ϼ(=�-9Z�]��G�YW"v���q�\�+؏G���W�����-蓺��bEn���*h%����^�
K��˹K�3��ѣ��?��}���ڃ���������XM!
=Xo�?|;��� -^uf�G�"#�;=Z���)�I�C�CT)u`C��w�E��Xz����[I|�>�8��q �v�����������Q>��S6�#c˱Τɭ�l��lXz��9q�-�=��E��ӊc=v<nZ�P#7J����/�<r�g���3�X	�1%�[w\%���z�+y׳|a}����>���H�����S=�%O+�e�DN���/L��M�'k:��f�?�����NV� �_�4�$#��ӈ�'K��ɒ�ҊdT判�*q5_9I�d��̭�%A['��	O����j�:����V��A߭[����ڝ*�Yx k���n�ի!cW�8/�P+�� ��mk먽�<���]�d�p�3'+�&aS颢#�����NVUv_���X�mE
�%��xY
�՜�^�6�d��û�s̬�9��r7=p����)�A
�"�0��؈���[��(����\M����,@"��� j���0��㪆��G��o�V��-�^}��br��Fa�u-*1ru�0��p�����QǺom������a��8�5d��+	�!/Y��b)��U1J���\�a>��u���V�r�Қ)J����֯� �(x��{$�<!N=ٓ 3�+X=�����B ��B9���&��g��� l��]P`�S�(4gZEk9L�2ɑ�ʄ$�|��T/���Uz=|��?�a���<�|s~�n>�e�S�	�]C�\�L'JA,�����zd� ��{{ke��1�*=�
;ɵ�nu!hY�d����YMDw��gU�C�_�y����8Y�x������N����{��PM9-��J�U��������
��U�w�W�8���Yy1c�)��>��~�=$����2�8S.rqc{ c���mj|�-ͺ��|{x�Z��{�ۣ��۵��6B�w��������%�7m~nG{�u�M��Q�KLK���*X6V�KqalJ���SR��J��`���V�ٹtÝv��Gmn�F�$�Ɣ-Ãq���~���U����OVA���]�������՜���qT�ЩN�s�t�����#�{��*7� ���j�+�Ў���)Ԕ<��L�z�Z�Ѱ~)տ�'�L�I(�&M ���Ll����\��#6H++�އ�6Re}^�2�lyE��6�q�Ͽ ²gg6�H)N������S����̵�3�(|A�/���yX���B���І4_A��G��(/O�'4���I��m�<2mΑA6�w>L�4k|h8��
�m \��
_]n.�]s�]Uo,s?���1�V���Ó�����Fo�.�-��K�߾�b�@-m�X���2ҍ�Z���(�[8$n˹�;{;��wʡ��\�����_�El\tъ�Q�*��]h״<;"%�z�1�E�290�G<�@���>��GvQO����JZ�_p*�hwZ:�<�)p��ep073Җ�����R��=Y/ۓg�귛�
����mb]�>q�	򝶕{]nׯ/������|��u�-,��Gk;��m��M7����ն�����������۶�f��l;�C�����l���rH䈛�S����p@�ۧ3�,E��(d����U�q�T�i����#�=i��u"�p�eW����#'�-!�����r����؇��8r����_]���#
n~ʱ��%NJ��#��ta�{Tٽ7��Cx=wq%����,a�G��O���Cz���������T%����F�#��u-�ц������RwB�ߚ���M{��a<:Y
++8����P���2	�#�Q�� �1#a,|�4(y�X����#Tb�q���isssmfv'k�-,�g����T�{�L���
F�B���� �y��D��sxx�����8�av`���r^V�dY����������a�.��/��0�v�����)���c{��������N�WS-�^���r �Y!� �{���8��G'Ke���j�3�%]Yh7o��'r���x�d�W�a	
Q�^��I�YV'��q�,KZ��Q�\GY4� �;�_�p��q��lmo���:aA�6���6ζ�:��#�Tۚ]KO�|!|-S�N�[�A*���[�y	X��B)-��U�q*d��ʯ�?���I�2�?�^�(�j��y�WZ)�̑��:�"g��"�@��ҽ2�$����\>+�ѿϧI[�+^�����?��*#������;�m��e�r�*�G�B^���[�������Z�ԩ�B�C���QF
�Α&��l����S�Dr�M�WJ�o��y	��B:p?8')۳���9d������<N֛�y�.���s�m5/�OC�;뫧�a�蹖򺣅�O!�]����xX�幯�z��J�*iCZU��J�Q�*09���*C�8YWp�ZV7݇s�צǆ���L{p��ս�!Fǭ���t���6מ��5�M~������0^��Q�x4��!.�ŗ1�,��'��o�;Q��=�)��`���i+�7p�����t�J�F�/3*�����?�@�pޏ(0��-��������a?7������e�E�,J�'kGtow����F���z���2�Sշɀs����C�?s�/�6Fϒ?�
�.2_���Je��q�	#�Pf��	L�G��Gz<3����!u������<g�O�1��\�����Sag�E��AK�1$)���[�"�)g��3�z6��ॢ�N�9+��|γd�<s-l�%|��o���٘G9qE�F>�i�.�!�A�n�����)7��Yh7n�h�+Kmz�Ց!!�l�."uqͻ0��y�:#~���v{�4�E��_ߋ�з�����,hΡ�q�H�!f:X�3�4.=���oѡ�:��;�I��(�y
��Gգ2|�mh����L������p+� �VDᔲ[nғz������{a�^�hWȻ�4Ӯ_�Ŏ���v-�����ܵެQf�?�Z�%z�zT�kew�0�C��������v���69Y���e�/_��O�e���y�NX'�ݶ���ސ��'/�+�wΟ6XqI��
�q����D��nmne���o��֠N�t�E�|��-mWo�4CY��8g��4"����~t.���a��t�r����ԑx�:Y"�7�zȺ�z�	�0z����{�&�ôr]q��J�Ay.%��}��0�X]~���u�p^+w
�gǅ�|Օ�ţ.h��Pl�N^$+��ޕG���K\{����.�-/eN����r���� ��,	�9YU}�;�:�C'˞�=YY��L���!ˇ<�bTv�"�HЮ8�ޘ�9AaN��ζ�k������Ν;����a���m�"�س"_[haQ��F���jp+��՗�a��ɩ���c��Q[뜬�P���c�]���B�L�sw���R9�N���(�b-��0�X���Į��NA�١6v_��	�X⍃e 1˧c�3���LbT�����ztą;�O!�������:�
\㉻c���{���$��\�u��d^K)x�Ñ�Q���j�,,�Lk(l�r��c�w��;6�Ǝ���ĉט
��܉8�u� ��R
_aRuܯ�gK�m�}S�hW{�K�۴�H�:����6?������nϝ�8o*F�8���
uoѡ�~�}�ܣ�#뱞z�B�_�{�}��Y�i`6���8<����Ҩ��Jz}��!L���g�����Σ��8���r��U�*�t�_���3f��jA�-�ٺ���6�w�bq�<*���h7��j���krr*�;�̕��6�a$�;����٫o5s�Tj�K��p�PyR#����q���� u%L5t��]�F�KC���o��(^�,2*���]�%i�+�J�toT�'/�p�*��:pX��#e�.�=ʤ�ٙ�v�Ƶ��������������ᶻ�6޾H��^�s8�l�(��r*`J��[Ɠ���:ᷔ��!�|����}�l�E��Q���J�u�~�y�N����&��,�!5JJ:[҅���W-����5��wਣ�1?9w�;th���K?M�>��@��{���2�y���l��lOO-�`̒�^� ����)ԓ^�no������<�K�-��%O��^���4�l��=i N�WΗ���x��%w5&L�Q�H�1x���#b,�P��r{]4��9v3W���r�2ײ���<�B,�=z�����񧾗�!��������U��,��/y�!�u�k)Q�U�	C�42���r���/K��+��J޲�R�}j����۵��v�j�p��
��T,�LS�y�wǬ�$οrć�nh�[n����+���B.��{�\��F
��"m2�lϊK�O�;j�вϑH霬���ˏ��W+L�G��w��F�>W�e�[qD%�0��xn}�	��:%w�Aҭ�5��e�ی?�pk�m|d��\Yh�ݿ�n��n�H����w޵׫k��Ы׫mk�&l\���/���^kYpIU��;??��.>�����C�LO����>{��}������~�>���\�̽y��^�X}���������g���B2�L�%�遏����PLm�͍���v-���4� ��8*{RY  ���.��Ζ�$M�th)v�r�84��Y���d9-�߾�t��AS�)Ik�3��K�LG�v*�G���m��(�5��w�So���z�wҜ��}C�z�2RV����|,��
����uo歟=�x6~]go��O�4t�k��̕8�Ʀ���$e.�$NMM��E����4P�e������7q��ɺ��%�+]�C㵜,��ʳ�Ri�Z]4uVaR�T�b���w�V��mEs1[��F��{r��J��|�������ￇ�u;s�l�qe�����x�z���"��M8���P�rX��/��}���[��Փ�;���ɲbS������=�Y�*�{��/=��-�y�F��"��[�Z�ߎqDt����"�r�������:˽�W�\"�Q�W�d9FFp
�%uuF{�n�Z���o�Ӷ�4Q����q7b�,&A�*S��Ki���7�C�F.ZB�Tv�P�&-�T\1'sPF{�(��	�\5t�-����M�x���g�#�0�qpB��އ$���Z%m��+����"|M�\c�QaC餂�0��3d0f
0R�a�`H}���C@����֑���]�7i�g�%0{AR��7
�|h�y�����в�P�_�p��d���{��'�Q�Nw���]Ѫ��}����pcN�Q�yt�OP:Q:�*deS	i�,��[�/�z�T-ڜQǝ"O~Č�E�������ܮ]��t-=Yʌ���8W:Y�.�V�p�r$�sFb�R�4>���2��9��a�c��RI�tʀ�Sq,�4��>��/��ߩz,�����`}#=]���v	�^�X���|��~��X^�iw�\o���A����v��R�nG������u��q�Ͻ�%Li%'�6_6�侜+a����rO'��I���ׄ7uI\W�u��k�n�۷`��l��yWH+y��a�����܋�2�.�����x�M>�����|hy�w�_W
UK$�:�J���y.l�����z��ˏkЋ7�)xS���'�,b���>�;�-)s�6^��W�����m�PG�hUs����~6�F���t?��z�L���*���da�ka0F��3 ��@��]���<���|���(ꎺ������	^��]JY٠>r��/b����>Cf5�5�I���t�|�*1x->�y@
��OҪΕ{f���Vf�3�3"���q�t��9���H�e��/�M���ޝ����m�kG�u���*mY��i�6�j^�s��k=�K�KGZ��%	#��1��܊��*���l���	��<�8�~nv{����l��\�9���F'kd� �q8�˷g� 8����0�qd�84_(*�g�Vo�2
�R�6ʸ�f�(�F���|K�q��|�ûw�������G�mwn/Q�Ql>y�E�޵շ�?k���aV/��`i1C�a�/�����N۵8X.vq��u��j�Z.���׿��oۯ�E���q��ֶ�+{���nO�hϞ�h����u��������s��g��!޽ko�����<saI0�����q& ����kB�(:��8�o���m�n�7�'��8X*��֬.u"����Gw��v;v����g���x+�BxWSv�p����������{���఻>8�o,!+\��/�LG��^��xѕE�AM�Ƭ�G�
�t�;dj9���`"7M7��"i�Y�t�����_SS�`��K�5�D|���t��o����㟯m���'ˍ���txR��*�r\�4qj�|���dQ�)|K)J{���8Y|�0���Y����{Ri��֭���?|�>��8X�o���|������S麘A�0
a�KGE'�q��5�+W�DRz�`,';��8s�6_|k��uQ

	Ɋ)����H]<4��<�W���+�}p��t���<������@���!�R�QN���"0�KN.5#.s��Ͱ�}�5����[�Gp��������҂31^��Wi��ތ�e}�9�eS�^e��̥�þ�r��Qf�P�p��?�`9��0��)���eƓ��w>C-�f}����PT*b���%tq"1���k�U?���: V��O��g�Ԩ�U���<*i[\z'��3�9��:���M��SWݵ��>��uPS��>!�6�`Y=G8����GZ��Σ��D��^�6��������Q�ї໹�q��y�Ο^L!y{�k��k����MZ�{u����^p��1X��K�2*�){P�{�Ϝ�B%��qX�4����;�歛��r8��nm�U�^�_���F[5{�GmZj�;q�G�C�P�D�i��⺌���� s2�
z���V��(��zP�����"�A��@��	�8�:����8w~�<=��07�޿�>��a���G�6�Cɶ7Wۓ�?oϟ}�6�_��mү���!����9�$Ō,5��O8Q��YI��\��y�jT�'������]s�������ͻmhv�! �{坎�r�Ƣ�>��%��Sݳ�W��idC�g]�G�2�N�}d���w�5�g�E�q�:���#=�"77�Ӄ��eA��9I*�>�Kq�y��������Q���m�NO|�=�,~��2��pF�۰ku9|���j�l�K��|.~u^t�Mҳ�.�vA	<�ʅ�\����{�x�#Q0��u���,��x���-����b�Y�R�' ��<�bwu?��7o���J�+��X�ZuȄ���������^!�6`��}���	z�����h� NM������`=�w�ݺy=Ñ�|X~ձrΧC�v�-.�F)�8�G��^N����@��n�\���^.��Y#W'K�*āCL����+��+������<M�zw�TדU_��\�����h���ɄC��<S��^9˼��#��q�8��J��ߓ=)��HSiVN�.��`{����G?�~��ѝ�^,G m휴7o�ۋW�	o���΃<��$���9����z�`�6�s��߻�>���������݄]�W����q���~�>���W8X�_��lɵ�����6��]��X�Fg�=�t\�#ĥzK{�e����ً��8���8WS��W��Ûvv9`6�"[�N�8�'�<��}���V}�V/6�=��nP/��v}Y�߅�5���gfQ�Us��$=�Q��M�ݎ@��F��z�����ݮ@�˕*�nʍ����u�{N՞q8�Ќ��RiDH�m��q"�$?�G�$�������^�+�����\x���tI9�^'k�MR��ԍ��,:YK��r��o�������N�������j{������C�
�HT)k�8�E�.Sd3E�*H��
$���Χ ��5���dO;���|�>����o�Źئ&��
Yt��	ht�`� Ą�q��0�N�����@~��8�c��!�`����y
��=����ȫ?7�si[ӑp�0�S�!�W���=��j̟Jݡf `��%N��v�\&��]�����+�ѡ���d���S[�e�#� ��� ��Ȑ �`�S.+P���D�f�i�#��%E\'�:6|nv�-/L�����ʂ+�4j#`� �sZ2Gjߍ�w)�L�7{����c���a�n꧟��~|��7@:R�p!�+��Y�ԣ�ﻙ[�4��iQ�R��g���l�(�U�7�%a@P��z����!ޓ�-�A1�+=H/�FQ:�����Xķۼ_L��/춘��(o����u2�%F �*��sA�@ �H��g	۸�����ѥ�OH�e�eUyK�
]Yn��)��4�&F�߼;��e����֦�ֳа[5H�|#FM��]��
<s�Kñ���?ҷt�'�[�JS0��z���>��!�}�{���,r�-���������@A�'G;(BWd�S��,�L��z:r��<� p���s	�("�R�rp���r�Z�v�z�{'����rh"09�kc�m[}���
�x#2P|Z�����']�@��]�;�9���/⤹[��-v֡)@1\��3�O�+����ԣ�L6j�`r�!����<ql�C$U�6<��eㄼ��C��k��A�>�k�����mj�J���|�~�����r�y���_�W/�h/��v�ހ��ل���C�.�˧���U�c�&Z�8y��,�T���hx���GENyE���6�t�-^��fo�+�8X�����&�.jMMX��B^����;���}ܳ?�(��,T2�s�2�2POq*S.y�t������i(?�+[���ڛ���5�|�|��CJ<��~��R�=G6����ꪄ���Z�O燺T���ϓ2���=�����b��ha�wI��Kȑ��T��%�խ���!+m�;T_����D����[�Bc���%
-���++�|��#oFVBG.�}�������:��5��m:���+K���һ2[�~��uJ�p@�ܓDc���.G��|Q6���%�;�q{�߹iهcJ#١�n'��ܦm�Eo�O'�h��\]A��id�2����70"g��4F%J6�S�ݝ-�񚋣�������ai#��Vlw��Oe]Ki�q~jQ�
�-u�\�G�O�A��	�R;�9Y6��&�rx�+=�`��1��"��������HV����t$Я��"h��%%yJz�P_���$�l�s|����_ŧ�h��A6)�q;O^���1�����o��O���9�x��/;ck��j�}��I�����󗯰at(+<��{�A����	}��nAW1�gڍk�miq���+C�:I����ן�����k_}�U�o�А�.�_Y.n2��:�	�a�ù���q=EG����yt���i�ܲ1���O����E{��Y����Y�H��X�VؠDg/�w���.GO[��TF�Q���
5�]Ɔ \��^�ؔ�
�=ϕ	֓��|Ĩi@[�R{��/�q�6)����0U{�t�fgfq���`�RީI�q�I�)�'�i��^�U6����B[Xp���8�9O�*࠿k$��Ex)���>p#	��~K�G���P8Ծ���9�.v�6��U�#}'=�ث����6
�Y�݆�q�uaq�-��R�ԙvK���s<�H�Bb����i�ɳ�Ew��7��@�I�����d1{�ڵ̿�}�V[���Dx�5�it��޿K+�Q �b@ky�*D�aK6�\��\5�dh	���P����A�ٌ�,��a��F�Z���g�9_䩷����I�����D"J�Bڐ�`����<����X<�F\X�"��3�l�x��r��u`׬+�)�&�΋�j|{�4XA�}=���%hT���+�S���R�[�� Ͻ,\��lA��jG�&�~A�ZK�1���w�f�N�o���0L;<F �ah`hd%�3�RM��k�4�Ʌ�ըD	����0�������L&߸q�ݼqa�0�������$�T��B����:p1[�%мP<O��V�cH�T���QO���M��J����ӫ�J��xT~�T�(�J}wF�u�9�(����I:��C:��EY�Yס��������O�_�;H��G�T��gw�ٲrT�H��)Ћ'
��B/���UWʁ::xs٧	F���O��௎QK  ��IDATq�������9�!=)о�6Px����'/�sA=�'\*W*AQ��0�#���K�o�J�+���_�_�N�u������ѹ�$	{���gpNf/Pkk�4�o\_n?��G�������>�8\����o^�Ǐ�lϞ}�^�z�ܼ�Eq�/�{����F�Ȳr�Ļ�MCI'�sHǑ�.�i�ȋ�j���U����
���g=��ѡ�p����A�O<z���u�N�t��Nŋ�p�B�Uݞi�9�3`��K�+^��J[�&�x���s(��<�V0�ҁ֑gt�<fKq𭑏㤣�#��!v����b��L�`D�a�G4�m��'�=�� ��GS�ˆ{J�w{��S��l-w���~D�)K~HK��V)Oz����ܓ/(�F����8K�g��g��k���ғ�G2d24�&��zIk������= Ҥ "@ݿ��G��s�c�	{�@�.�)�r�\����R#?�0���v�`gSa���
���l�]�`!��5��mnm��I�l�{�W7���@��^�v����ZYY�^gӞB饓�!9�ݹ��y�
�H�q��FGkc�;L���:_�K���f�{�|�=g%�.}�um�;T6#Η�ޫ����\��c�л�q�z��=�y����b���ɋ�S�K�!����}�ױg�V(�ڐe�8I�6W(��{/�3��>�9�1}�v���/�W_|�~��_��_}�޼|�a�o߬��_?i���/�8X���͡���<�o�Cߛ#L�C�u�\�g�O%��cgOF�z=?̽����a�>�M�:�i�{�,��������k~��v��݄{�������������Ç���k�=j|�a�>�3��O��˞Y�FޒW��ءx����\kd@J��`|����Gw��:{������D� �r�q�#���}G�yB)<C�ﯻ�2�w�O���A9�D,�{��.� ��� N�@�0ƻ�*~��F������z��~�[�]gE=�!��S24�zNH	�ჯ��%pbLq.��=#�W�_]x~��{����F��Z%U<]�줗]��C%d+cة?*=8	��ĳ�gT���|8�a)���+��r����5�ff��s��e}��ιr	�,^��ϙ�ٕt�)��u���.��c�mɩ���P`�5r�����5>�B��T�k�Γ�qȂp���Fo�څ�(��Ͱ��)�/�_����5lzj"�7����7u��q}�-..�U���v���Ί]��t�ۊ�9��u&AU�����'���w!Zν��M��>E'���E��G�q��^'8�dn!Fk`x���h��O��i�[��Sldqx!t嬣������q�:��}�}2�縘RN�,�'��r�\��[|��S/�z�v��{��o���š�]9V�V�Wŵ`,�Rm~��w����a��4n��@~���P��T�9L�t*�����׽��ɕ��}Ց2�{��r�6B�ۋ�l���ÚN0N���P�ym���{��I���ғmw�={�M{��q{��yV8s2:�u��0u@�!��Y�p5b�)6��W�FN9�ԝ��BpXߦ���Ajc�Ζ���l�B�xK�U��������'�Ԏٳ2Vƃ�0C��WO�U߅[��*c|i����!n~���^q���:�]y���R�)ߜ����ur�Õ�p�O��ĕ6?;ܖ�sF����$w��K;m��u}�^ҫ���a`��:��N�y����s"<��Jv����x�oF��ݢ�G}g�=,:���r�Ꝇ}�xw<�ϙ�F���q8���#��i�*�����ޥ�+�N�b<e��>u��k�:.�a^�п�ח�w>��"L��g���>a'?1�pQ狺���ˋ�p�zI��=:`摡\8\��^qb�b>4�,)�i���D���9`�-/���3�mn���>�FOCӼ��g<���W΃_��L0	�se�{y��:4��R�l���钏
b@y���u{��y{������r&#f��딅�32�P4.��e�|B�D��|0��2�.�@�f�f��{H>�ۛmok-[W����AF&�|�5���o���g�|Ӟ?yڞp��_}���'�~���o/��	����G�>���j�>��S?%��u���5���W�wP� J.�Iq��?NZ�Ƿ�	P	6jHS�S�ɚ�^\Z������k�K�������|�`���8d7��[�۝�w8�"�u�ԅ؂�f�*���ὡ�w=΋s�,$������;����{�p𤻪ԍc�������z�~��;`����K�ڣc<oJ���┡��RƵ�`r
~�%���9@Gmw��lM��D�8��U�*�����"��`(h�C�Q�;�@�J��Q~ϑ�F�@�i����}������O��ud=<>�[	9
��\�0��0C�K��++��W��1�=+b�wΖ��B=�#��4����<O�k�s:8-���G�dY_{����1q3�ԡ�qf QWq��/��k�x��Pt������ᄇG:\Ё��0:q�}8F�c�j�w�t��ҭl�;��"'�-��k�
M0 �����U)�PX
{{*������`yi�]��Ԯ����ׯ,g� ���V�@q^��&h�H�UO���t������On�V��w�zZu�h]��@֦��g��E�eZ���`�� �� �pq��Sh$��fSL��P�^��z]W�T���V9{(��8����ws�+~���4~�A�<{n�����4N:'˂p�q��>~S
F��ܣ+�?���ʕ��߬G�q{#"t�@}��p��7��qE���eJ,�/��M�G*�+��sz␼���{B�MՕC-mX�¡���\����� q1����63>���Xj?����'�{����m�����o?�e{��EsOB�29���iނN|Rx������+�˞��Û��ݛ��ˡ����Иc�2������>3� �<����G��s��9�`��;��v9gì�-�ĸO}[���PC*y&�ro�bV�!n9Z�)��~흭�QW_���+��?�mV s���췑�c�� ��H��,��Ļ6>�߆�l�hm�G��'����0���ڑ� `��ܐ�a�P������V�-��1���������.�$���O�W���rړ>����s�흢��� �'�^|}^'����[匽������9D�к��+q��b\iܴ��8�䥬�!�]d
y�E�8����z{��M�����A����ٳ��9�=�ܫ4=z�-,�ht*"O�+t@]�ц4fɂ����{�І$�)C�=��f�p���Z��Y�e� �T9PU@y�OL+�T�~.��
��_��7�pj;��l��������}�Ǘ~C}�H,r��AD�i;�Ό�_��]�Uv&�v���Oo�\k�<��}��G�����+�<���K.���?�gz��d:�E�\��k��7���~�>����/��ӿ����_��z����t�n����.�<Fd����;�O���a5F����o�^+D�s|+���z{���W���	�F���e�S��@��s�i9w�*2�iZ�yա��{�lyy%Ι{�:�K^�.���3]B�)B_�oݟ?���<�gޝ]wR�*��}���D�Tc�6DQ��9�0g pCw�<������@��,�)�M��  +���MѼ<�w�c�l��c�y�Se͛U��|�.p���o
��r�7�obl���IPEd$Ev%	,<�����*Y]!�����#�@�����yũO��a�}	iI�*B�D�Ԫ�!o����0z>��R�A'�W�+?�[r�#a ��--ε��Y��eD�o�u����ب=_86�j'?^T��w8M5+�r��B��N��U�r��h���=-N ���r�^*�5��q��r���q��ګ3fD9YYT���vL�@zv����^`�1�C�ܝ��Ѵ�/���l���ZY^û�͙�G:�r1��R�g�WD��Q���{ƭ��PyE�r��H�g�^'D�`�\jD��( O�Ϡ
��Ī!���+φ��{��Y	Ǽ��X���밸:5����C��[G=������۳x�:{���LЉ�3䝟�'pa]��4�xf�m�բ'㓏<F��/3���4ĵ��������p�J�@y�E���М��[y�t�7]=��yU�c��'{ڪo�t�<�
~Vg�+>JK:V=�:�UGܐ�	�j���z�oې�����βK��6=v�ݻ��~�������v��
�~{�����i/�~ն7ޒ�XBc�W-˫Ѥ1�A��, ��SҊ��3_��@R�0ro�5��	�rB�8iı��{rl��0���_�ly�<�b.<�O~��j�+���Fb|�О~���k�*۸OUN�t�����3��Z"�ԥ%"���c� t���!�tHÿ��Q
�S�>��Řj��6��ۆ���� 2t�][i+�m~�y.ȡ����ެ#�y�G띛VP�#���z6_g����B,���|�3{�Q^c�ϲE�AO�)r�2hL��׹��}_��JkҤ�Q8���^��|..Iב�GZ�����U�ڋ�"m2���1꡼��Աꇋ�ӄ5��0��;�E��ip�|K�n'�ffo�:����C�Mҏ��`mmm�����}�ʶ��J+eg��3��}�����.��1n)���!NB?��|�cJ�� �K��sq'��7�X2�4����+�?L�g��b����e�����#�8I66&RlSe6�[SZ���q?" i�bw��mn�dናC��F́6;1�޻{���?����W���o��i��Oq��;7��g���T[�ž�!�fo���Y��q�^={���o����/���o��Op�>kO?n�8`�a*���8ʌ�3eP_�w�H�wqz:NiR^�oz=�ԃ��/��r.8s�I�v�|w�'�I�]gx�FpԢ"��p(�C	�z2>�*���a�5��8luzF�L�nq��¢�2gK�LG˵z�B]Z�'�Ͳ[�<���g}	z����u��>���(�y�?z�Hz�=�y_�H|h�$�?r�D�~��vHN-p��*x1K �y�s����R���z�!�d}FW�|����ŋ���_�/���}��Y�km�홠[B�1��Q�rD�L�aշ�b�� ��a�
��<}0��B]_����w}�쨸|CeD��g��s�ҋeK�p���W�Y�u�
VhZS�y�ޏn������Q��Ί�S����s�Ĺ�-^�w�k�,,���t�pXA�F�C��QYxC%��Z�%H��Bޡ����;����J�[�s�����B{���&�cEPqV����� ����`šw�U�,m�:��!'�祌���g�'a�0�=h:r1n"�J�i0�Z�B�]G��L����l���;t ���=qI�:�g�Pk ���,��x�2F����y�cp!��v�`OF�mnG�˵�rt�H'�V�M6�L�MmX��<OPQ��B������u|�U]��//�	GpByK��CW�#k�{ST	kxh@����C�w�-}�x{L4*��K��)5��V��9:��1NW��j���O�:����(�#FO��x��Ψ�1���֐gߺ�_KD��-f�u�B8W�8"W]���e��h� �?���Zj���}���v��|��!��ɗ���~�^>���WK�0�@�cF:M�k�`��K%��T9S�4�^a5�|v�SM��-q5�jX��W;�?x���>$�!eE�B�Z%�:��O|�E,u�з�z��㪬�+�JZ��F����Y���Y�|␆���?rdx4�}�Iܵ�`��8d��u��!߇�r�:��C'Λfz�c��>u�<���#.���~�׆����@[�k7�'ۍ��8}�M�n/���#�q���G�h(�	p��-?� �hJ�X��r�8xn�A��u�8���X9��8�UWד�vV@��.T�F���w���T�2�?w��(�"�����4����)Ⱦ,=��ųj���@pVʫh	Gpo���
��l^���Qx��d�mi�$p���}B��!� Y_�4�0=�R���'�VtEE8��LU�׎x �UU�i����IO�J���!��Źn�/���wR�Ѳu�Ǫ|D����_�����:q�lr�z�H!72�	�F����K���AK�!}��o�����/��#�|��K�w�Se�N�i��q���꛵���F�ElA���cK�3��of����������������O����>m�'?j�����G�k�~�}��G��=j�?�ۖq�\�����~�����i{��)up�E;K]f�H��dѡ�[���l�N�t20��B}��g���r�q=���<�_p"��+a#�}��Q�t������O���D�"]���[�6�CrO0]�%�5~��e�@	׷`��ɸ{��u8�v�s�Y�V�ӽ㿇�[�.:_I?y�i�#nF�����UF/�F&~!�[�|�,�F�Jd����$.
i��M�SX{Wm��}�����8.K
�l�L
>[]C�Ϟ�h_|�e�����o�s�d���PW�qxL�� �;qc1�v�t�僃Kmg봭�ﷷ�G�}���{��zZ�֏{=.8"�w��!�}�>ɕr����!+ZUV�*XQŏi�C��}w�v��վl�V�/��Ͻ y�[-_�.O웟q�V~S�U�ۃ5;�P��v���5Wtq�x>WԏHӐ��s}���r�Α�cڕ��y>��]F�G��A��j(1pZnߞg�:M�snL�W `�����-*�K������S�>:Qm˧�X�.ء�S�j!��3<�?�&C�:\���q��L]}H��Ri������/��,��	��{�[Z��H�<�I��&�B��@�r�i��	�.��^�<��-��X��C?��%�Ic��.MV�H:q���L��+�NM��sh�? .����/��h~�)��{q�S��k�Y���a���*����
��K�vNwG�������,َ���BYP�bS2�<t�/�a0�r�/��a&���!���&�n^����Vp�V\��@hB)J���"��[�/��;���G�ٯ�f*�x_�m�Oz&S���8R:oY���Ҹ���8��^^=m�s��n>��ngq���`g�=�
W_gn�eh�ޯ8��G�t4x��>�#��Q� _���`�KE?�z(�}��z��\Q'�\#�Wfs��<osKmnq�ML�a���> ���Ի��3��_��]�#G>�'}D�_uPG�c=� ��`y)��t ����[W�|�����0YW6F���#
�!U� A�ø��儕f�҇�c�:��l�t�HXR1�	h���@*�9�B�L�>��G��hR���Q��u����l"gz��N��[�qP6i^��؅x�**��{�{y�V�T�����&q��>���m��T��i�}�����@!�����/��$�-g"��v�:�����C%~kq���q�Qh�፵|���l�����|?:t������$:h�*L�q��i?r�a�
.n�C�t	��%R����_�[:h���.�e��C�w�&��.������Q�F�=�S����4�s2>��e�yǩ�IvaС��ş���`�� �r��<S沭J�	������܌��se]�(��Qp']�g�az�f-��l���������������8�M݌�9��͡���76�g�.�C�^r�iז��nj�d��AJ8En%1��S�v����g�����dA�͛7��"S�N�y�c�z��\hZ�+�{%�:?\�J/x&�sz�v|����x���6���<���րϺ�/d�|�p�����t�?�#��!Sڕ'�Q����hk:�CȜ<h?���-][��k h�9�Ÿڂ:��DH�Om�M��Z{c��j��N�����#a.�L���r���|^W�:;��a������Ш�V�[]�}�0�ځ7,�U�ːǹ�Y�:�^�A'�}�@��lF�% :XCh[��pV8�p��lD���Q
YN��$	f�C&3�q]K,k�l���m����A�֞�x�s�U����7{�S�D�}�,��M�iK���\�R�Q2�S��يR�G��7*�J;h�ӶIw��v�d�"���*-��+x�l�D3�R�8�X�/Cȇ2K|�����:u�Y�,`��HDc17f�v�'��FG�g�z�`�;�!|f�ʲC��̌-�|)�%� �1���P��q����ش�����;�@p(�l�R����D.SGؠ>a������3߅:,��4��L�xJ�g+l��7�Y#[e_\�M�->�ǚ��4�%v���cݜ@�����l�X:@K�c�i��»���u�]���@1U-٣�c�oM+�u�|�g��RB��*ϝ�>d�'��S���{BuDs��.v@ȾdI��6}�K�F��g��(�#jrٗ���|{vܟ��礛�|U��J�UYŇ4,>��ʃ��9 �X#�lB�⯧W�w&�8*����
�c���*?�C����`�q��0]�o�8�A���Cn<b�!�
q�T)�ƪ½Jy�OB=n�n�\Y���#��zh���0U	��Ea��w��\!��ϥ��#C����X�s{�=��ݿ���w�mo�m/�~�^�`9K:t�n��1�O�yE����,g�3�sF���xH%�ux����뱮b�'��#�L8ϼs�R�b��/��9���6BL�ӳ����ٵ���?rt���>�y�Q���� ����}���޼ho^>��z�:���)-_j�(��s�෣�'��E�ޙbe/f9�i>��P�O�f�����</��{�%YZ����4\!W]r?��Iz��R�k�(Q �l�,�@��Y6�%3����q���{�����MW�p%۬f�ux�/���+4�B Oˣs�P�4��O�i�}�t�u/K�D_����*��8Qf�`���Y#Pg���δ���������s����E��760�gj���v�_���n��������Y�Ǩ�j^rL�k��Bw�r� i�lao�Q��6���ԐDt-�t���B]jåN�8��dp`Z�!�1})}K�հ��a��GElp�
�ں
ޕ�r��$}���y�:� ���lD�nC��l=??;�f	�J�Z�$pK�ص�ߴ7o��_���"�ɸ v�B�أuL9�[{T�0��1�o߸֦'Ɛ����-x�e���y�j�]���nݺVj�rǛY����tx'�'Y%�y��ViQ�L?<������(H2���5��,{��)��x'NV��Z}_�6��ԛ����l�O���Jg���#�w�8�А�q�86�P��{�J{љ���{���i��:�2�QWKc;Ю������KAK�_ �Ggvww.\ǶJ�D��U�����O��o��7���S���p.-��u��߼N��=����t	����w�Z�(�j��;�cH�����V��D���og����߷����_���h�W�~��_��p��?�r�����~��������O�>��g���gq�LW��aS(��2�Qy/�N'�+g���+�z�M���G��g��o����
4ԣ��Y�����p��%���$z"-�WH���B�A0�c+CMp�c��a[L���<����,a�zn��gy'[8T�2�-J5g�6�W%��J�Q�{��08�X���n��ؘ-|m�q�{q�"*%��bk�8v��mq����&�Cᄛ`�qc��l��|��r=���5����cp�9Sn�aB���5õ�L�5�������� �{��Io��5!�C�?�(�"S�::��:O�ѡ��mx�E
����e%pm�3ޝ�Ȼbػw��P�y#��r��=Á�hP|J���r�g�\�>{�;�4���ك�u�����9G�SH��=WʚzK�t�iXU+j����}6�����Y_�8.�1k�Ű�	Ұ��`�0N��������0p6$�x9��,ʚ��Ї�0t1��yN��}�I#W~m�H>�r�gu��j�B�^����v��J��f[^��������œ����mk����(��'��#�{[=;z��,�/>4�b�1ҀE�؈�CV���:����򳸡2'�:2�1�#���4�4��y�3�� ���a��*XLXV˅�*Á2Y>B�	�Ӡ������ޗ��Ƌ&퉈|<{_4o�gA���+u�t�\SN_��t,�K���ԓ��.���n�N�-��.W}�:"�	t���Q��1�I�=z�B���x�ۇ܎�b���}�2/g�oT��6���D��Q�X��x�w�_�+�J{儊oeD䃩�7�P��7<�Po��]��]�{_�<��u����O�������49��U���t��m�����0����^��v��}?�toϞ��4���pC�V����Q�;���~��?�U��n
�JI@:��k�ɧ~��]��L�j#$��'�7�W�Cy�h���������D�
�6�U�_j�[��ŋ�훯�`��>�]�aY�:��hp���m :�i˔���p����K�A%�q|�/GR�]�N������'�M���ա�6==ږWfڭ�������r�ug	gk�ݹ{�=��������/�տh��_���G?�4+�@X����:�Y܁�_iH#�sr�g�������Tw��>�/�����τ�4����+]��J�\'�P���S�<�AEO#!��"4�P�_��4[�b�SO�~�+�ځ<��j=���y�-��U������+��(��L5\�:3�#@Aa|h;�S���G=�8�:��[��J� 9{�kE(������wB��t�:O�<i?����Op�~�ӿ�\,W]Q����N�W_}پ��ӧO"�$|��������n�&^@�Y\�?AL�_��x�?���?R�� �۳G�Q8���aB�J�^J%!�LH|�q��
2��U9T5T�k��D`Kl�3ӵ*)�Ҫ�2H�΀.�'/��,�3�^�%-��n���d~��'tε�Q9Zn>�ӕ�)�Bd�+��
p\�!��ؽ�Ʋ���Ɏ�hA:�2�-_*%����KY�'��z��1a }�w�X��ťᑆ�.J+='sh��)�\���2��n�q�JQ�4�Cj��3��2�+����y��$x���Q��sH3u�NU�����hg�,W���_�:8W���*���-?�(U�a;�!��.w����:ZM�ђ�o@'y	GWS� �\���?����3o��;�vߜ�w�*�k�dG�V��ay�dN��-�Ơ�UFU	FC����C'1�1bl)��֡9Ҍ�.�d8��yo�i��徇'�s׽�V���~0v��"~gw��~ήy�4�g�yD _	���
RM/�-j����n�911��nn�XnK����/���8WY�g�Mݝ������m}m��{5�
�1V�Ȗq��'��8��L=���l]�]�oz��-Gp�s�Hk�uC]X�>d�±Û���?p�&�J��?~�S�]<��n�ҊSxW��xsNH� �'=ÿ08q��\���"#8g1R�vN�>��v��S�6D�@��h���x��q�+�:�:_�2��x*�GHW��lVŕ��y��NG����cm��1B��0do�=��^�,tQZ�q�<2?��O�ٖ��s�v�g�� ���hO�M|�7�З84�Wt^<�<�	$�
^W����o*Q���z���K�u"��&'�S��#eo���8Aoq��oެ�i�oW�_���{���3e]���2����M�=�E;�w�N����ϒ�����ܛ7�q��#i�7N�Y#x�ui�W2G�O�N��%.��(��{gͣo6bh��)N�+W�4��VE�%<,������;��l�w=��obc�dy���1�wΕ� {���rE���Oфܛ�/�G��gO_�����h�"�
�5_�{M���ȩ�Xx��3��̌�����?p.׿��������6x���mV�s�A�J����h�	�{{�����u���;��C���9�}]�~)��G��c�#��~���`��n�yN�wI�<f�.���(�M���-���>iro>U����~��K<�Ì���L�<W�zt�(�����j���"�Eɑ�o�;�W�����d���oڳ�x��(Q���S�ӟ/����0�]�� ���F��X� �T(�L�;�TeQ�*dg&'��k���۷ۭ7�˹��:�g��P�����!��v��F�9,le��ԯ����s�r��;�#d��q��S���V�+m��r��=ikۻ���y9\||���� ��h&ҳ�՚��<�q�H��ڸ�����Ec�V�Be��^�V:k�����^	������
��dB���r�%�V���H"Tq���Jf�VG��C����̕693�&'Q�CmE8b}�.�<�^����_�o7W�/���f�x/�>L�Cm �j��\�}dĽ�t���U�hZ� Y�=/2���w��e9dg;�l�?�\
ŉ���[�l��'{������%m0������̼�h</:=v�BU�+8fەg~��>"/���c`'�ԫ�):!�&� �:
c�������s�B8u�AC/^k5�4�)}��E����X٥�>5�D�N�b��;Zk�����:��?�B�j'o����v���yh�I�mAR��_±2=w}��Ѧ�*8��S{s4��������{�%�d�0I_�	�|ؕ#e�\\*�d�|*����*��8s�W7t�c���z����nR)�T�5y7�=��e�k|�5N5�<q�%�Tr�w�،B���w�������-r�� �g-��=�i�'Y�i5��8�p��	 .q�aX����o���#)I#3�l����LZՁ�q�q�5ih؆��_a�K�^9iC��C0�c5���K{���v��T�{s�-͍�A⮿~՞~�Y{��Y;���D��@�}���P��vLY6Ťe���C�"ژc�[��u��(�����U��������Z��|��Ρ2���m�tq����6;���smy�Pe�6����A���r|w���?z.�Cǵ��מ<2��9������ �O��12������o0�_��v���d���F0ab(jp�H�3�<Dj���Ro�i@��M�8�<��T��hU>)�a��NG��� N�����B��f��ts�?��|/�V} �s�n���G��T�(K�(9Y��x�^]J�c��$8đ���3��'�S��+ī8,;%�!���֗4#��|h���w��ɀ�U7DJ<9�Ά����֑!��!K�3c/-����
����;l"�y���n���S����z����"�۫�/��'�5�G�i{��9��K�l0�HmmnfZ���z�u�vq�Ї������54�I�G���~���V_��/]��Y{��e�X续����S��\ViHǪUw�����Zbޑ�0s��N���!���vZ��8ʝL�'��:%���z�N���=��՝�(�)o��W�)��cGA�NGG���ۣ��o]kS���@칧/_�g/^�յ��k!2�W;��y��}7H�RאS�G�d�@��SZ����>cT��.��ݣ]�2�͛b���XM��1O��gml�kj���ܾ��l��ml��P7�G8M�EJj�W��Ѻ���mbx�{�q?7Z�d�`Y���Q��=K��#�S�j���Cĉ��z�a�3Rv>&�`)_���%v�������U���"Q�Rپ������G���Өm]��T���K.�Ws�6��re�K�cǂ�ֈ5p �s�p��W&�l��^[a���㛄�z�,*=����z����#=��`+�R�rV�Ѿw����㟿�ў>A:'�G ��\Ԙe,@H<N�tIoU�L��ڈ�#�7�Cq��h� +L��J6����������G��[7�go�7�g�I�g=Y��%"����>���ܾٖ0�u��L�R��p��Q|{��o#Z�F��o�̹�ka��'cY��B���R�ܓ4?g]��&S쪎
�k����Uq �<��͛q�}�q9wF� ���>%���$B{�4$i����=SxS⮡B�� q�Ǔ�������0��΍�)��e޵���
h����n�wa�珂F�At�ԹJ�K�OP�8����$hX�ٵ���ر�c�C�kIe�BT�ll���EA)�MT�J%fZ5|��+��&[�;�H�_�UG!	
/[����=o��L�����������#�U���e!S���)��cG���E�Q*����>�ƭ?��z�AU��ސ!�&�Dt�x�NT,YNYZqq*{��kՇ�]`���H_Nh����<-���DM�'�֜�	�x`��2�K�s$J~�fŶ������ן��ԛw��^�(�g�+B���Ojl�ϬCWc�A�޾���pP���|a��}OV��N*�I�4z	�??7߮_w��kY:V'K���g[7ΣT>�C���'"�F�p$���3�R�ֹ������!	YC��T=�[Ґ�X�3H'�.�ʙ�S�A�X�z席,ϴ��W���4
�][[}Ӿ�����Q����9T�H�}ﴫ{j���K�`���0aޫ�䇌$ �2��m�#iE��M�X��T�w��B�_
��)���c�o�힝]h��Kmjv���\|l'�V�˫>�譢t1�������������̷��o6������}�#������M�щ�~���L��Q�д֒���;i�0|����~�(i$X%։?�a]��|[�11�I/���E���a�S�l�P5��1�4�b�P&���=�"��7B���f�ҹ���^(`���H��@,S�}A<�8��f��4M�_|�����N���A�3�~��tȇ�c�S4"�]�/�֙�u	������is��i왾�dO���;��m{�߾��/��gO��gϟ�:�~��,{�:�S�&�ʝ�>Go�
*�W͗�L�Ԫ�S8]�]�Y��^�g���Y�;�F��g���j �a��j�(�T�i�;'��)�w;��P_7%�&��S�� 	�ԙ�?�A��8k��w�he�zUzⅵ���	͗n�vJ�ڛ~|���p�][�m=��>��.��r�	2�������r��W�}����i����6�La �2�vY�����<�p�c,t�����t�Ƿ�8�n�<�ݠ|Mq(N�%�X����[�= J�<8q�$n����g"���L<g�l:�6J�Hi�3r�Ls�|�x�@|T|�}��m/(g�aV	%ZO�JF���H	<�i�jă�Ҹ8��U?����Ȩ���,��|f�]d_���C�lxY�t�|�͵�ohQ�i?UJ��2Wў�Mi��d�װ�4�^Ҷ��.��9Է<M�	L���>�w��q+����5?���H�<���n�����ʼKic������7k[����;YY]��N��S=YT��!��dQQټ/�sntD�y��H��*�U�0ʯ�������8X�[�������`9Ѧ���$�]��<%�Z��Ν��G�ڇ��n߼��g�c��$�֎�Et��t BY�w�p �T�mm�b���������J���J�����L���7`v�ߺ�9�&c��p:s���r�WM����/�%��O�R�ZO<e�\�~$��iAq%�A7~�=	F�p�|6��5�9#�2�iSR�J��^��v�=	K��6�/N������4��t��T`�G0��\07���K�a�,�q	�����/!�[��@��t�lճ����T�w�o���<B��4�u��)q�s�;���+��Q��Z0�#�}7�,=lm!\q���ev(@�i�#�d��"\���՛e��'+5_�iX��b�P���g�Y���W֖A�@Ed˱
]G��ltaE��J��k[K��R:��0�O���tr&�rB���W��p��i�#��fU�<��d��ٳ���қ�G�&��Е�sNfsᬠ�*l�d�d��0e7u?���LR8J���ܡr����Z�R7�R\�pUං�?ǝ[���;w2�cy$CS��鐞�Bb-F��E�EJ۝M�/��j�-U�1Ɣ��!
^�eW��s�/�ʱ*��������<WA^�����Ơ��*�k��ɉ�8Y�Sc�=n;[m��6F��Yn�=�s����������2Na~q�M�/���9��4��B5N6wX�(���S�B���LE�_	N�Ys��
��
�@���Y�@AY� )����� z@'krj��Y@��"�u�}�s_AJ,��'������H-����츐������C~�5?����z���ϑqo����u�q..�=Gfh�iDԆ�Ǒ�B���|5+�e��BE#�� @�e�����C��:��5�����Y�״��)V'�
�z��@@�����u[|�W�^?K�7����o� ���\�jxur����'z��.=�@KT���~�Z�x�x��<v�r_�������<���3����1��M�]�"_��^y�|*G����x�ƍ��������w����r>��V�r�-��#�����Zk�]�j��G��:��^L�p����yL���*y9$�-qw¯�s�d�u+�dQ"�%�+o��칑��1��{��8O,�s�C�Jz�٥-Nu�\N]޷f3�)��ـlϜ${�$�8�Z�O�P�mH����qfz����v��������z������W��g�ګ�o�Q�`�����Wf��p�:�6Rh׺���qv����:�:�=+P��{�m��^�Qz��յM��^F���) �"��S�����c��g�T��D9(?�'AK�e�չ ?%��.��P����=X�0��euA��W|'?nKG����<�C���f��BVe�m�nn�g��k>ˠ��G}����,�Z}P��z�H�|gg7��ʂG9׆%�Cp�/�X��]��������B�?Q������;��X)r�.tV��9V�ٓ�6	q�p�P��1�o��E'k���У��:Y�"nA� ���ꂇ�d)x�0�@e<5�#>�Hл�nA�T��+�\����o�wC@�Ric�mn~�- �K�*�-����K���������}���{x��&1ګU�Jtll$v��C$�����.N�=Y��a���B���Z��]DS�l,6��T8���w�,�r�.]�=N�ۮ�3'F �E'+�"Ε���z�����`	#8Scc�Q��ؓ5���898Y�n�;=���YqX�*n�wը|��uZ�҂�bIK�1��9X:I.y��35צ&p� @�z��KY�ۡ����C��dYo҂t!��2�p�Ә]}�&��a�
]�MM』���(0�"�\�q P�S���bb���5�$�J_�J��Mw���� }ˣ�5yCz0e���`eu�8Z�d�p���杳�����N �o����
��U<]h��t�'���v|���Zg��h���l���A�g@i�\U�Y�ђgm	��H?�Ȋ5T�UD�Y�ɓ.T�rE��S�\l�%���M�g?��x�/��|,����(��+�t��ϴ�0n�5���Ke`�<Wӥ�Y�r.��]��<y�r�--/Ei�H��%j��|���_-�@ha�^"�a&[ 3N5F
iȌ�K�8G��ϪB`��蠇�sɎG|�LqA�A�!���YW��1x}vf,�4LO���Q��vE�m��K��d�v�f�y�n�{�A�o���nsm�u�A�~�n[�q�-�\�67���5�&qp&&�������vw	{�	pOil�ИU�:��!G:YN�W	��T�5&r,�.�ļ���P�5�I���'�!��z��|���o�ߪ�8���󛳫��9���?��z�;RW�u(�.6߶�/��?��%�d�_�S�l�	�kk�6 �^�B����ˁJ������8�m� � �	#�E]ڠP�|��Qd�������� ����F��h�G���r�Fy[J�%����~�m�|�\�����B�4V2�����_�AH}��7�����G(�w�Jc0�t�����9S���a��S9N��d�Cu���2D������-�%|8����ֶq��R�*W��
,��!WԨ��ʅxv��A�"��l/��s�WCU�Q�g�C	��7T=;�/���q�8Y�͉� ��Րf<iў,j���fA��ɲ.JT��<��vUBxT޷�ӻ%��K��M�b�!��a�9�Cp����Gmiq�}��G�~�Q�}s	��洺)N�;8n/_��g�qdq,�w>k���QO;4�a��{�v�sj/�۞��{G�)�Mc�I��e�ņX��\� ���F{��e{�-��|�y�'O]�Ì�%�9,������!�O�������pĩ�=��A�D�¢u����|��t�z^�͵���x�ҡ�9���T+� #w_�����nm��>�w�ߜN>g�� H�\\�$K����m�Z��N`��o�;������������@���ٽ�ԡ�����cx����J��*�����5�3ДUW.QwW�[6��M���/�Ѭ�]�F>��5�m{kFSY����8��{e�p�Îxq�,-J��^���˨ ����ПK��y�|�ƠG�s^#~q�W����"�U��>��]#��H�k����U ?����8�)�%H�1�BE)(A��N�����H�c���;������έ�1ӽ{�H���	��\[_l�o��PQW��:���?h�~�i�����'h����䴡�Qʀ���0M��+H��t��Z�,��͌d�n#���R\Jg&��g��To�;�]5��i�GB�`����R!��R�.����|*�ll�S�=e�A�H���\���d��@w��x��9�л��8�V��,ᱤ�TI�o޽m/_9��
mF�g��J���1k��r[Y^C�C��^��i�\��
�4IKm~vK���� \∕�=w5!	c�+���k���f��jG.GK����alhQ��8��ǐw��Y`�GBe�3�<ذ��[�:G�N�q�7��_�� ɹS(#S[�XS[/��s�L�(��PA��m�W�/�D(F���B{�nb`��
#��3����C�@��������ýsΥkhL� #E1NK�*�Й���.-G=�<�������k/u���v�S���?n�[f\.*)�>K�NQ����Pk��u�2%=e~$\d�
���ǔͫ�FY�C���+'��l{��a����gT]���i_z|���h���5���.�^c`��#��K������">�(3�Iん~m�b`��
�x�@��h���)��5����rj���əv��
F����S:��g�}���矷O��i�䳟``}�>��3.d����ƽ�Ɲm�ֽ�~�N[_��V�60����Z^]k��kT�\/�*܎�����C}r-U�[����^,4HP9T�oi0}�W����~�ԛN7�Y��\*%��U��G�W�#��=��4_ߋVu��>���� ^J�	t�3*p[oQʞ|۞?}�vw6c�L�RhL��MG�UHT(�A��s���m{�(�N���Yf��E��(�$
"�2���^y�x��_��� _��v�p�t]f�	Ƌsd�#Xе��9�F,�+y�4��2��U�#A'�y���oLK#�O3�)V����mr�N*^d���T�2���Ɔ�k-��
p T�[\t��r�0�(WF]���|S"�qQ��ɬ�Rz#�:�]���7��n��P�R�َ�ؙ ���'nL�l�ڬB>^R񦂽����*G��@�R
>�Klܽ��M����J�n݊�+�%��8]��*�F�S=��t>#�4�!O���2�*�]������\NCe�	F��c�Jy�'����F�t`���֙r>�7�9��rmn�Ѣ��Eq��u39y���]o��?���������nz\ݎ���N{����/��4b͓r c2�A,�&yZw�4�`P]PO�6X8��r���Mu{g��e�V�Wov���_�o�}��y���'�믿k�~�=j��wt�#k��\�����早�Et������ft�l���|R�?��<S��������u G������7��z��;���aœ�	��l�OzJg�7ye���������@�H^�NJyQ��F����L���4�����L��5�܅S]�,Gd��|F�4��A8/�65���>I���.C�j��g�P����.��2G�4�=~�Y/��?�l@Ddo�يKO@������p8]��q~�;S��T��y�gy#
�{n�k�MUf/L�p8t��#H>{5nݺپ����'��O�O~������;w�D��7iR/zpD>*$4d Mal�+������9	Y�x�Ĺ�y���A��cB�i�(sW��Qѳ��Nط�@�@��9ժ����
A�Zoa�h�l����n �b�:_�ic^�2ho�D�����£��!�P5�&h�9�l�s3��Q9t�������"^�>��C�[w tv�`��>3%Ĳ��Jg��;]z"�5O��6�����D�Lb�Ȅ=õ�" ��w��z;.FwC]�}�������Ԛ�ݥ����P+���N_�����:?�gx�/0�.�w��������>��4��+�#�s�Q��lx�F��{?����o���;�َh��r�B�tV>GM�\Ew����Y`@$H�!���U��vx��W�8��^7��K�ǽ��Ӱ�� {�UlH$aL+B_�z�� ��(�N3��������g���/\�{�@Wː'e1�`�4�6��D�i��U��R�)�.���F��p���Ԟe����ٶ�*o#e�r�g���/�Y����_��O�Y����	F��{>i�����J�6�H�9OD����R�]��:��Ɩ�
���'?k_�������?k�g��}��?�P���ݸۦ�Q�����y�W�+C�A7�p����/�xy$�jMƔ����!2=�{��c��u�}�K7J3�R��5��4�k�������zB�cܕ$�s�g	�8�{uP��nTaϬ#�pF���!���Z�fo����E���$���<5]�yV�����K��[�F�J����A�D�nzF�
�

�	ak�F�h����U_�H�����1K�<�8Sb��[��ѯN��ڂ�������Jd�i���F��@�W@�2�O;�=>�SD,a�H_ʲ�|cG
�D�K�/Υ��s��HF�z}��S0>��pj�A�y�_�x��R�NR�s�y�����Q�s�J7�ШR	�L'���z�w��ͽ��*���:8OG��>��ݽs���E�2�EN�����g�}�<x�ҷ�r�"�j���[X"i$���Mޑ7�w�/������������5��hم� ��ĳ26�?��p��b����q�����M�n2�L�~C�N=���kcS�Ғ�����C��.^U���t>�|R��1�w�r��+-e����b����L��}�}������������_�����������������_��_������?�M�������w���_�_����髬��S���#�|��]Tc:H�aי:bh�t8��f��b�l�L���3�:�^����s$�s}�����~�8��s?z~x��;x�t���� G`�����q{:8?_�W	�����+aH���t�D���\��~���|�k~��|�8���7�߁*����C�jI֤���@��Nz�xE�w魂pPn�םW��)�Z��;���@�|�*SZ0�>����1�����݀���#S/(fPvG7\�T}����B\�a@��!~���w�";����L��q�n��W9U�ʸr�F)+�Ù�)ϵ�Q��&7���6����Fw{������A�;�L�Rxv�ِ����Fష=�=_UR<��N� �d=���\[vD�85	L���C����Îf9�"�I�y� �h�S���Rݖ_�����A�G�o��އ���i}6��fkd�����e,|�륷�EZ�Qn�����ي�|�#>_���}�ni	IWC��x{�T��%�(�F�`hq�8��;���x׀:�fNU���'�Q��u:^�Ff�~r�iIN=Ҁ=�p�k'VG�\(�x�wch��6�L��)
x��H��.$�k�y��}g G��}��%�C'�E��u	�>u����(�weX�0Z�G�q�����J��O�g9����;�>���pFِ��k��$����5i>�=x�aJ����5�Π�M�P�i1�Z�3����M���m}�5�B>��ݽ����'�����>���v��Cd魶���r�!5�Qum�ܦ����\�8��R���umj�ML/�ə�6��֖�n��?h|����������������'?i�o?hs+�9�r���鄮��ѷ��M�k��
���k�u嗎�1�P�O���)r6r"F�8���2V��l*D�/�z���3ސld��Dж�ȑG�ww�2�(�=����rƆkآtJ#�T��I��\7��l&ah]ww33J/6�����:�҆�S���9��)K��=��}���x'��!��Ea��a�5-�R���#�5��M8ʥ�g�a�ᨘ�+4/��L�R3���5�~R���]Z����/���wNx�(B~!�ܬ��+�B��FEޔ�5��ąy^�T��w��A�]p�_��d�Q��eӶJ�y��w�y������+��{yV�����}
��&Q����df9J�{�WWW1��/>�I��O�����,>]&q���~�����O���O�?F�Z"��ONR6ׄ|��G�#�$G��t@8
�r�i���Swi'�!�Ұ|�O���}�[Е�v��ɰ�A�k,����Z˄���P��A���t4.��^퀂��{G4��t,/�	�W��_�L4�[_D%}�څS=���.R������sR.iE�_�8�0�Q�9��r�b���?�����;�2��΅�=o�}��}����7��7�=o��l/��n�^�m/���־��1��ܭ>j*i�n����m��H��{�CAj{R�4z�5%��uM=���#���������C}ׇ�8���f�f*���u�X����mW���G��y���n`����0�ʋ2�z\���K�n~����gh�|)�%���_��_E�3դ�ϥSׇ*��J'�vڎ�ݰ`Q�$�����6w�~�K�C���E�E��H���I�a ƞ	{�*�\(0 ��ap	K�vbvv�-,��<7(=5Ǔ�G#�F��^X/K5���8{�_���&�J��_���p�UWW��F��K��p/QX����+�W�g�"[ڋA���h�,woqq�S_�̎7���T �;�R����L_e �
�`�F���"���.duFnvv"S�W���r[s+yw9��UN`>�+{j���y��u�X����P�E��Оl¥�R�%l W�BYa {��V�}�;x������R�y�N��A;�C�2�Y:�6��»\�฽���}��:�f]e�F-4.-xp����F��jJ��a�k�z�ϩҡ��k���+0�;X{�o<{*���D8�G��I��X{���1��r������s����%���=�uZ��W���fo}
�Sp�]�y/N�έ�X!N�vM���r�$t�L�]�H �U�G�M�iTy	��n� �f�8&��9��|Y�[\�?\U�35v�d�P�'��S�o����T�a٩�����ܾ�������?i�Sg|�n޺�Luڏ�̐�9 l1��]s;t�������N�h5c3��1�ÏMεY�[^��|�Y�􋟵O?�Y��ӟ���>l�+��t�=�0�:"cy(m�E�(j�ſk���үýB_�u��5�k�4�����H�Z�^C�ý���{��Yu:��7�W��y�����v��溚ׯ^�W/����M�9��q��"��rP�;-�M<P��*���i�hl�r�b��s�3���k�P��Ew��{䛻���-RwKmzn�#z��I����J�dMZ�AhY莏eh��.n��B��������u�2���?o�ZK�mue��)���HY�,�#vӐ��,���R��B��<#VC�x��C��;8qdZ���FW�J>�2�+~$%�,�yM}�4^�ȏ��xc��Y�|7m�f�7ST[-�w��i��ʹ���v������7n�V�e:��S���ǟa���}��O��o�}���:;�S���-��Y�t���:a)�*Á��U�k�����c��bi瑣r�1��"7ĩ�\��F��x:���艄1�餳NE�0���Mg��||d����tf�NC�s䶠u������N�T$��*ߑ(J$�u��0�Qg�ܹ}����������l���ߵ���/�_���]�7n\�n�̗�������}����)��.�x������^���6eK�k�^�p
zm,�	����M�&��;�6�}��?�~�I�����wVԏ��u��{�t"^�G�]���(���΢���i��.5P>�]�h�;Ȼ��v
U{DU�GeQ����@:�0	V�F�(��-=������=цt*v���(�%2�d^�^�"A��q���?�~" ��^ɸz�� �x� �޼��K �Te� 8:�'��ˋh�9d[ʵ�m5@�0!2A2T�4T���l���_gZF�I��O��\�:1дU
��Te@���nc[#/�a��Z��J�-�\k$������/_�gn���Q,�lyM[� �|��H�M�ku�V1u��s�`*��"97;E��D�����]�]g@%kLi���t�߆̺S(J*���{�	��qT���IObK��U�67�p���zvQsZ�iF���U�����a/�
&R1&|MjFqU� |]֩�|�������Rw>Wr�K�+:M���;P���P6�W6�pO�cu����9xַvMY�@�ҘB0�x<��3�v�B4�e������p���=N|�Ph7ց�V�m)�8�i�
� ~v��u��PB��=�|����� �U(;%k3�ŷi�Sʥʭd�J�^:
|�J:�|�0I��N#W��7i:��뛤s�z�m�"|���tF4�'�AGA��_n����.��k���(e���>��ݻw?����ih8�1B�;�i{ns�2=C�����fX)������)�O����9�P�WV���w��~�>����ǟb��E�Z�I��)�("���R���8����h�F����vS��ͷ٩McK%"!�ͫ|8<�}�g9+�z~������|�@^q���P=��흽�*�/^��ܳ�����՛��>bj|ˀ�'�خf���v�-^D-#��+�^�(�!����!�\#�����x�ݺ{?����{H�=h7���v[Z��Z���5UaVq^F�_��(ԞKxf��U�,���[v��	tz���Z�_����!�Xrf�<A<׈h��^�:�Z×���T|�����=�ն>���&,��u���@=D~E�SDܪ�پU�tg�q����J�U���m�Q|� �A��	O�uC����l��&Z*��4�i�-�Nml\o��=h~�郷o�&���
F�<��3|v�n����w�d
�mG6@���
�%��}h���)��e�F��2�6�2��w�,S��yxq��R���z�#TƩ6�v� ���U6ڹ`[��/�ɝ*���;�n�Q������[ګ�?���(�	M.�_���9!���8ӼR����,;nΠ;r<
�f���������������m�����������?i�}�i[[_K�dǬ#�v\8j�R
0������*hW��Q���6��m����k�k�_�E����0��C]�R\������G~^G��v�!.�������xޙ�pJ;�.��W��kD�f6]��U�M���s�r_��:��OG���R���_k�K<_�0��QG��O��*x/H\� ]z-We�i���m�A��2jNÎ�O�����˷���p�}KLj�FO��a��k��1,M��C�A�*�I����L%�1��"�*�;L�s:�J�1\�PU��BI
Xw�����!�����E;T���ʤys��%��|���a�WzC T�������nӝ�.���y���18����?e��P2ˎ�^�^��m=��*?��ZeTyBl���x��l�nO�sc�'=�ƍ��R8�Saq�G?�ɝjt6�3nz�q�����یv?N�(	���]�<�Э]evO�wW��
�
�JP |E���<����}�+Fpj
!��H}��I���薎�^�A�.��2k5��@ nIS��l�dgA$��"m<6�1uk�ḻ����	��V.Χz#���Ã�]0{p� ?t�$�r�f�z�J�u�y�|�<�YYS�t8�1V_؋�ҙM3BG�-���(�2r��z-�pd�6�8m�p�XgІ�qr�:�ܞݭ����-�UbP��_)��=xi�� >��8�`�5v!O���*Z��Z�h#8�r�+1ˆxeT���t������(�8�-�O��,ÖQR���0�P��_�h������%��l�mxwΎ��;[`��!�bS#B*�ES����.x���,-�7S�-;"^�p�à���ʵ�#k]*l5������Ӕ1��~���U!M��>�|Es��;�׸r�����YþjK�Smcu�ݾ�����޽�>x�}���о�D8��AD���'���lT�Z	^kk�9^�r�Qg�0i t,}���+�W�r
�8�Ok�k�;~���Gx�������F8�1*~"���˅Үi��s�3�:�� �g�����v�\���T�|�_s�z3��.����i,~���$o�<o�|�����w� ��Z�Y���)��@e�IG�����8�[7��=8h�F�	��p�B�tj�#��(�+�nJ���{��a��Ï�}�>��c��P��a`y.ܭ���&F�+k��.̟Gn�{F�J�� sF!�{qn�g)/�6��l���/*!�ą4O�Π%E�)���.�Wҥ���+u��A*���V��O������R��Wq�>�/Ʃ��UnR���J�r]� ��c}�w�Nt
_$͢e;�\C\��|�CT�8 ^Z��.�wJ��2B����k��.�Xow��-�r0Z����^�*�Ϊ"j;q�֭v��ڷ�Le{��I����,~Rf�c��]Y��C�p��$���Y��g��M=�a���j6#s&�p�dwC`9>�Q�,�l��4]�B��3��t<�,�E�e�q(L�q���+7�� �c�NFhzv�ݼ������:qũt����~_~�-������N���&���q�Ip��S����wo�?��/ڟ��/���g���e��O��s��[��wb�Ϛ�t�Y["жk�M܈{���v���v떣�����9�������O��W�Ho�&��؋h�_���W�+�	����Z>����Fǈ~A*�d�.�U�����*�@��I/�9�û2��)���������o��su�����4< Ĥa�E�\Ӥ�p4gY9���g� �Q���t���0x��vd00&������F��}BQ��zLG�g痲	���������Z�2ݼ��ܙ�����o�����O_���uuwA��H�*����Z{�]/�H��� Na��W�ͧU	Ѹ!{rrv�Q
γu������;�P�����d���Ϟ���/�cm�c�!=*䄵��!ޙ�b^��C�� �4%�������wA_����{���)e?��s��W�%���{�ih5�g��Ή@U�Y*D��/klz$��a�P�8:J����_x��9�Ps�% ��s�U?Xxq�S�{�����������=`"w0�@A��xO{�4����߶�ͭv��׎$N��:�Q�r�����@ڛ����y��H��2сkx<�rP��_n%����8sچx�$�9?'��==!�创�7�đ-�E7��/?Հ�	{U|��L�O�����mc�F�ԙ�_?��W��Px ��b��[�
ʑ'߃�C�3X%�άA ���W-P�:�( 4�<w?n�*��6�?�l��w�1��O��=�4D�T�jJ 4��]�۷���P�Qd�*H<�kg�;���z��H�`�&0�]( A��[���Ma�?��X��¾znP����6��S��H��^��kI������(V�P�ĉ"^їQor�&
�i� d(dS�i\��"_��,�񑸃&+��h���M �86,�� wj���ZP���P�yH�ӧOi�7w�rڟ�/ʲy�/*���r�jRTed5&��g�7�y�d]K	Lb)x�Pv�t�x�AI[��D~��4ʹ�N���D���L]�o7�r���{�����w�h��ǵ;򵽸�ȏx�l9ǟQg��iwgĄܕy�NՕW�d��(¤��E`�ȅ�a��<���i��:Q1���d�2�?��m߇RB3~�(�\�&���2��_��0\Y	<�f9\��nȴ@��X�C�.}ӼC��8����f������W8�Sh�hE�:"w�y�����������m�yA�Ӷ03M�5M} �
e줬��ȁ.m�_Ǯ��#
��xQ����}�i��Oʹ��������}�>���Ï������v��g�~���m��C�Hϩ���u�m�x�6n>hk���;mn�F�^XkS�m
�b��F�j�f�A�P�t"�N�;{�\�9��K^r�Ƒu(�ܼe�����cTÀ��9B�q�k�׮���o��;�0c�;�DeD�Yw5��(_.��q;ͤ#y32��JN���/��m��R݈)eT1��-YRt�IK�'�+�,�p�Ff����lp�#;G5d��;s�����nz�Y�O�?mO�=Aw�F��mk��m���������˙Z֊��N�2?�/;g�M-�Զw�.'k<0ލR�|�s͝xݘ����]��.{�e���Z�{� �%y&�(ԡh9�|ls�kм�U68�o���:e����R`3���e5^�y}�-"�a[�t���������U{�������P#m�"�vN#?N��X��=��i���Y?��c���>ո�^�+P�m��3�0h�շ�t����S�p���<?I��|/�{�o�4�V��2����v:��v�ڣo���~�е����"G0�C����b����}�y �$+�S���(-�WhU�
�52�C���$��w����-�<��Y4�_�8I�u��+���N�qD޵�R^=���|iǲkċg�+w��v.�Q5��(WFG�D�F�tL>�n҉�����^'
��� y���I��C�����fjD��v,�k޸~�ݽ��u�zpiێ��o0�v��dadm�g�F�J�#��Is7:{M��]3� :� ��/4��U�t2������'o����̑��l��_��헿�u�կݾ��ۜTn/򡇻��+
D�`���LNT�;(I-V�4�<<p��ɺh��'�'5���e�OP�-�l% q�ʺ,��JN�&�k*Vda�w�}� r���-N�2bэ�R8J���1-�|�����,{�����*��۫�*Ij��(~��OF�h$�d��(q�m�a�^�j�l0�|k���0f��|/f��6��N\M#q���~���2.Eo�9SB�Sfu���aPѯ��d�K1�������Xk�o�o�5��U�%����r���#X��BY��� ĩ6҉�`C>��� p�w��Y�b���H<�A��{FF	�/���n]*D3���|M�[�1�
ש#�k��q�>b���f9�B	-�*h��rW^���V��3�s�凂K��7�uM�k@q��(�P���Р�^f�s�.���\�����w�*[���}⋋b��$(Q�?q�C�H^��<��g��Z�\U?�㡛��#%�o�CY
8�Z�`5mP4���	Nw����O�5�ã�=�^�|�v��2,�����ڔ�S�Qa�YJ�b\���"�Y����i0Z^�
eGm9W�"�m���;�-�7�<�X_m�n;bq/���L5�G������P�)Õk�����Жu�}��K��o��	��R����?��`���1^���7g^�q7<�`48��j�0��]9�� 6���qJ�#I�Q�6]�#[��ɀs����/�"��~(w��>;��n�(p�ql�Z���l�۾��79���]��!��a�j��4��,x�ze�y\��j��RR�G�Hʘ.PO`;��7n���?h�~���hw�}��w/�9��PЗQ0��餱d{"�{f�#)Ό���g��f$k�-,-fV��Q.g1��Pu)o�yW�;�/��S��S���}�΁=#�����S��$U�R�>	N�5�	)��T�taV�/����c\x���F�� �3-�{�3;��ݐ���=�a[#]�b��x�8��(i�J�S�τ�Y� �?�v�'�7�Ӂ�״-Է�O��y0�v�R�r��u��ӧ5B�L/��(�ԛ�����G����gV�ӵ�W\(^u����-;������{G�m,��TiWǘ�\��cN�âq�dR�G�d�i���C�f��ԩ�άO�!��'k;�U�����aЍ��3�9����z�]�'��>�ݳW/�k_��ލ՜�r��$L��YE8)�wtңen^_k���n>����Ci&����j�����7�Y^^h˫�muh;n\���C��2nݺ÷uxf^���w�!�����0����z)����4�`�\vWo�n�<W8�Ӄ7�	7�Hg��r���K�E˕�����^�6l��fgJ�Th4��S
����u�8-PCI#JC�{g,e4U�t0���AN�tZa��9���C�֨X���X�pI*�˯�7��aNz�
6ë^�{������)��B;�cY��t����:W;�b��H֏YVm@"+�������\��\��xcA�+�ʕE+�qqwA�=��s��L��=z�}�O�7��~���-V_�����wvbيt����YϾ���4'"(Z����4����kmw��t<Y.Σ�����Vo�
��-¹�,Sz0��G(��5�?	����:z_Dn"*��QQGF�FΥ�ui�TZV�J��B5�Z(��P��ux,��L�Q&��=�XEӑ��RJ3-��X�p�}�9�aC� U�:�#���J��G�4�k������hd�7e<Ӕh�-8	�X)�L���Y�`��Xך3
^d,�C�ȩKKKp��s�W�j`9Cx��='2�F��=s�-8�%�R��b8 GAd�7-��	��k4BTPl�4p��x�s��|֣�!���(�Y�K_�ѹ믎ݦ�:��r�j���sG�jK:I��I�6?a���� �+!�˼�Koe����S�qJ��h�cF/'5��1�,G�Gx♆�U%��W�YZO��w!�=_����;ӤR0ң�ҭ�/&3Y������N�>UP��2��Y�v-\�pw�LϜQh��A�2={�=����W��@�T*�H�Dʛ�t/N��r\���w��P~�g�U�UI������ ��g���Dfz��\�B1�sc�ݻs;�	ܻx��4��6B�A�gd	��yF\6�_��S��:���\�RJ�AU��l=Y71�)z{yI�Y֙k���Jp3Ы_pߒhn�w��lCjǆ
+��l���H^�"��I6�+�j���j�G���P���5���J�N#s$,�-n�Rxz��^<{Ծ��W(�_����6�r����p� *5ă�Q�J�*�z�,iԩ�Q$�'m,�9r��s�N{�>����O��}��O1��$�f[\Z'OG�<�{��딉��5x�X�2�g|:���Vc�^\w�\A֮��y�N�!,V�`�ò1�����tӌS�f�z���<&b�;��w���W� �(�"�R!��=�+�*>Fo��s�����v��Gŷtf&���N��:�B�߆ހ��,:2��5CY5�XGm��i�4@�ӈ�'�Ƨ��)󶥅#��J8�D�S�ˑw�;�w݊rj���� �#���&��~9��iy�U�	�X����B�5H����m����,���j:��|�OED:��6��!�+���L�f݂���It�b�^��,���U�,��HG��wӔ;�0hn�A�l�Q�|gG����	F��o��� ��ԷxO~��t�)gye;�R��0��7V��;7۝��(/� MFG�@�yH��3s�����r�u�F�{�V:�����k|�0�����u�	����;a��I�  @߿6��7ߴG�����]��?��+��4ܝ�v�<Y��I���^�jd�OC�B� '��ԓUFB�]��0�C�z�K{��N��.� ��\j0��� �q��׬ݲ��3k�	�8оr1k��T��k�`ɋ���-zx��=���r�e��\ԫ��Fɍ���׍,ٖ������5���ک)m�v�v#�LH@@�"#Y(�Gܖ�E��!"�LF�j|.�����)9*k��s�����I�Z���oޤ��7_~�<���}a�<�����]���	��+�K�X�)
*���<�

@��GG��=C`�F�.�,��G�*�
��U1dH��5.|JE�~��*)�$<I���w<JcM���7ed�h؊�Z�'�%�6�`Z@��Rf*Fd��4�*��"N1�vMF�<N���O�N�SC��J��[ O8e��4�j�E\�۞�/��B���J!��ң�B��ŉ�q�v��FV\`�Bd�N2"���C���8�bd�~	#��0�>T�э��:d�γg�8��V�4{��\{s��ow�u0�pv�S]�����%P:�Ttl�T�9=�1��.�!��%uuI:L��y(�P��)�|��ЏPY�d�t#k0���R����΂�.�Lߴ5�����@��3h�����}�xW��'��s>�H#�z����c��|1.��
pJ�]jOyZ����+��+_/F�5�# �:~@>�N�(��/�0��m͢� k��a��I��⿔��Z6�4@fM�6���k�\q���pV�@*��7o^��8
����,Wdf	u)�_��\B���]�IT�N��x�t*���v�6e�!ʅӭ5V����H�;7��}��h�?|�}������пk�Dn��&�:b�h��*�*��*�ht�^S%�7d��y߁��U��)����Ha�C��,l����Q5l�t�:6C�a�Tʷ
�����u��x#���!���xa"��]Z�a��3?�K^��*������需J2;���K�������j/�߾�����_�7��g�2
� نEiǻ}�)I��S��F���!�Giy�X��>�6P
?l�����>��L�[\\oS�K� q�J%���Gd�������IT^y���v�9`��ʢk�4�f\l��)��RA�#�B9it�8rڛV�lO��Ҙq}�U���]�2k���(��kT��_n)��h�H��d��]�Π#{�� ��{�2��\Wb�`uW��cTYt��I(�1�/q��~"L�1�!�"��.�x��|]�e���Dv.,�S>��A;�m���6�4ܽO���ݻ��.ϳ	o'_����7�����Wt*Of�	G����
})��v�`2�9]FF�����`t1׿jdY*���*�s�d�W�?g� *@(��ˑ�� p��������ݩo�)��@��������Oᙩ"�Q��m�U>k��>k/_���U���G҇��$=Y�6�F`ҫ�8sc��ٸ�,tX�G�l������v��u�����;�2v��-����>�G}��q�Ȏ�t��Ϟ��~�~�믁�u��C��қ#dVZ�$`.���.]�m��y�)����*	�;Kb9�Ȫ���*a%c>��s*�XF�������u6d��	��&5�9TDQ^����JcK],�hk� sÌ��L{C9/=�Y��Q�_���6!�U�^SR��o�_:���'�9�d/�'D~:G�]��Ŝg/�ٱ������
>��?hd]n|�Q\��,���
�>��O1�UxU���U��oń2�1By*Sqn��h�-c �08�e/�g4�Ý�W"3�L*㺦K�teO���R�7�pj��5
�h���{y���ȝ�|��jdQ��l�,��*F��}��B�ϗ�]��W"�/�E�^&dY�4�Xeh�t�-�,�)x�/f�8>S�P�5���AA"��kd��۫ú��k;bXٻ�i��3]5b�4yH�̜DD��BW;����<���FE#���v�҄� 3f����קME�V�����CF��P��o�U�D���&`�n�j�z�����Jz�j�jk��(/N߳!Q�Qq��Gq���������4��*��s�S�����a�e3���3�58/�,|�Ry>ɯ+�$ië?��.���h���:����邎f��)�-��$e�AU�-W����	�<�X�fY4�2��-� �S>w[ps��8mЩf~K�(�9�&}{��{����l�+��T�(���Z>�F��Y镁e�5����B[��x6�*u�Ϊ�{���b�_��^�����P�̒@��(�X�u��q��"4�]0}�N��Y�޾�\r:Kd��"�T=uA���g�7�a�.��p�T�\P���}(*���9�\o93y#�h��m}e!�'>h�|�Q���ڽ{3� Yȿ�H;j��:�4'!G2F�g��F|��2N��t�wF�U��$<�p�J��@�gG��j`UҮ6��N��A���չ�\�p�$�eT��I�K�!��[H�D�L{�PR��;!ͻ+e�X�V�{�x��>u'�6��i9����ڄ�9�gϾk����l_��o��Oÿ�(��� 1��/�g�rA��L[�q3��/����j���������ڧ���}���{�?n��7��y�`P��'��}.��4@�kd����?yO>��L�ƕ����lOm8䜝Q�1���5�ȑ���Ȓ�e��T�+��O��@6��u*�`y�q)����K���:j⽵d�ا+��T�]���F콯x
��b�Z�}gۣ�ԍ,]:����5�I���eu#F'�� (�z琰�s������
핇��'?�9Y�anx��L�6gh�ʬ�����d��ƍ�m�]sIC%ϳ���c��;���Ehd.儔(�d�k4[�^ݍ,��f �#]�d�&k^�0,�SM[���x�c�+K�Ȫ2�S� 	������Qߑ.jz��]y�w�C^$J��J2���7�>��~���=ʿ�p��1�^�'.1y�<���{��>���j����^!lN�U_�^Ż��Ƌ��`~}��ٸ�27��[km�k}}�{)�,.ډ���q7�Nc�=s���'�������o����˯�G�3�rO�,q�o��ů��;��JVyӟ���B��]�X1N3��2����!�1+˒�|���<23_I+�:l��-��;�F~���8��H����N֍�2�j���z��W֡�C]���:z�kȍFH��8���!��Yߝ�]Nx�|���C�W8qi�}t���R�$p͢:��"��`d9�%])I~�,OO�J�_<V#KZ�Y�#����"Z�ӣ4_"��s���6�0}[����!{8e@	����շ�V(.�޽��:�u�`I�A�4
b�]�M�*F�v��C��h*V#�����GV��&�唏�hsdS���e.�3�<�3r5��AP�)��Ѭ���'��MyU�bl�Z���1���Y���S�OPf�L����E�{����c��9e�:�3G}���u#-�Xa�R�G���!����������:?ZC��@(�����^N*�^�}���&�&���œ
٩,/�/�_
]RL�	 ؐi��(ݿ{/���Kˉ�bl��Hj�Z��Ű����"��!�4�ҋ���m����Iø#Q=C$ҵx�w�󆦦�&�6	�J��[�:�A��6�As�W�,�u��ed�b��s��2��;�uMZ�"�G�?4��)L}YwQ\�q�F�7�6�d�0hkb��^�q�z�'쉛�%�N�3��J�Z��l��H�,��׸���
[�\�X<{�<��ሎ�@�mc��J
��*҄��O���76Lҝ4Hiм�%�ɺQir�)�ko�w1��f4�5~�e�
wt4k�|���M.t)��}�\��k�Z�g�C��^��kF��x�[k��͚��W�f���B{pO#��.k��)�9�U~#5U1vTB��;�% �OY�=���zC�]��	�䞲SO��2��8t�Q�wG�4�4��U�4�FS�8�!�F�I[���B[�)2�E�{�ʥ����on�eY�+W	]��Ӷ^�qQ��r�H�so��%߳���UvK6ȴ�������o0�����}{���=d��#��SG_��A�+}zUVɧҏʝ孩\�$��
[In �L�_Z����}�����e�^��^.��4@���fٕ��M�"���M�o��w�^�_<_(#�z���,�����h$��-�k̬G���zv�8�J_{+$���:�'hj�歬�N0��J�~
�N�����?�x��
�����!��xϡ�!�C���2�#�ʣAz!���ed������M��4g�[7��Oѫ#}�q����r>��g�۳�χeﲉ�W{�U:�{�]^��՛(�n�TgG�<��9�=}�|-sꕲX�1�g�m�t����R����z�ʺ<�y�,����I]�62
�r���ӎk�b$v���N�C\u�c7�J];������X�*T�3�$�i�榑y���{na�B٪���)n��������8�;bd�G��������N�l4��ϑ-�bJ���!���E��ܼm���8e�X�L��f�"ry~����e�4۲n�����o1���o~�~��7��k�F��y�]���TtE�U>�w�}����ҖĐ�W>�3��\�!�//N�s0��+%EAϏ����a���'��1����R�c�ռ�(G�I�5�U>S��p��U�^k��k��j�)X�����q�M~0�ղ�,[�������fΑ��2��7��p�=t}u���8��-F�L3�����N�.h�}��%�ӫ�����o�#~
�K��;��U�)~�L~��Ͷ�`�bJ���@�"�Q�@E޵fo�<D�Bm�ܿG:7�"F�ʓ�)	Vnz�
eqc��wt�`_���u����3�
u�U�����tk��o��K�y�'_�,`�C�ۍ,����B�ˆ�j� ������(�1^ciciaq.~n�w��)�:�^���w��b�8�3�P��q4G��r���Ҙ��zU�n���ᥑ���� r����I�*�
Sa��ф��:�0��V(������>�B�Y�4����zM;�q#��F��TfQW�r��naXmmncTc`�:�W�I�r+aϒ)c�^W��o������c8lm�Y�F�4FV�s�qz�#=*0T_5���:q�A�z����#+S� �#���}��D�5�􃐄ХG�
a�k���M"4rU���*�$��^����"�E�)���cHf�I� J��#~���ܲ�v�2\2��8�<:(I���c�����KZ�&�k�����Le-��{�~��q#�0(�̳
i���i��� ����Ls"�s��xǩ�ـ�X�R��j�(�	�x #i?��/W�
S����<oI�.`Ca̡*so�g�����X[�1w����!JƇ�;w�l��&�(6-�k�3:���N��;�z��ý�s��OW]��~1H|�a�{�)/7ո�� v^�wV,���Ec�9 +�ƈ��p�̽� 䵝%4�A�>;�o�q¤���y7�_IS�&��%�ܡM}x������8�D�	��k�_>i������o��=�e;�ۤn0��͞m�V��(WN�b����-5-L*��m�Q<��O%����_Z��)�~��v��'me���@0G�)
3D����V�|)��!3�'��������pM<=��s>��h)�
��xN�>�<IX��ѯI\%FGl�˗U��7uvL�idY�c�:�qh�Ѹ�"�:�Y^G%xG�U{\��>��-iR���ZF�;f�fc(�Y���^�SR��ik�?�N7�.�>#5��ـG���mB�H^ֻ�s&�#���ſz������]��˯����W/��W��&���em��lg��W_}��.����G��'��~��Ǐ'a�N,���ʡS ��U��F�A>X�v�i�;+CC��,��iP���1�c�E�w�.�d+��8�<�ŵ�4b��9�_5���9S��n�4?��w'��8}6�&HǵS���@�a��	��pz���n{������FF�m�pR*�.p��#Ó��K�mn%�{�v@:Ϟ�l�޼A�?N;�:W���v2�:e�g��#�O�%�:��3����2�n���W��oem����z�܌b��΂���^���*��kj;:�2�t;��(�y����7#�	�ːX�K{���D�ߥ/y�d�~yqS���p:<	#~F�팉�.��UU��YFV难�Z.;� �.�|Z�f9���ma���|W|�������e' g-�e��t�h�{�ux؁�T���]��=g����i�&��$P�0�:N�UhX*�2��)ZA�;t���o��˽���A{K;���̯�V �(��- B?���*�(X�z3r���
��֋˫���~�ߓ�p-�ɷ�]z9�7V� �CR�<\z%�K��Ҧ�r�qvn:F���B��n��633�jnf&�=���
Okw4�-{�4�l0hh �Z�UʱxMϱ�_Z4�To{#\�������3\0��.�u#���6��Թ��v������6�
ͬ��@��^�Y�%����J[[Yͨ��O���6�.�vʽ�ݶ3,��Y�W˭�5�l@z9CWօ��a�C5��BRWոW#[
\�a�Y�H�˿\�j���^��#�P�PA�货��G��2�����.�� L1t.��@)��W�p�U�Cj�!J����Ǝp�o�u����\�JW7*��%��//qD3}����Xc[��H"GJ�6��Q��������g<�(>�װ�K�kk����F�QvGx�{��u!�4-��EuM��l�8�T�����+��6��l��-�"�ݕ�b7���s��ٶ����\_˦��~�Vyh��1է�ѯ�U�e��ҡr����4?����*7z��(P��}0��Ebzy���V��1�i�V�;��~V:q����
�=�����u���N�&J
��~;��j[o^�����������;����v�:�ה���
��g�CZ/o�EG b�O@�N��zWe���������ۯ��o�l��=j;�Mg�2zR|��c�m�6��ۑ����I�(t�S�\��,�յ��޽������Qvt�Mբ0#�-�)I{|Q6��>2��t��\b�c����
�G9RyH�A���ЛHr�c��-�g�����M`۸�ͮn��j(�c(�*�1p�W�IR�$���65~��!�g������N;�}�i���>%�4,^� ;R�[f���k� ?N��2&�f���>G#�F^\�-�htt?�xe�48r^W�-iXZw�'t,2��z ���Qu�7�rX��\NW}g]|��I��(�{X�f�h���eeTE�	�w�뼨|Z��qqh�ҷ�$���[��ʄ�J���G����r+>��22#����9�s�%��:���\9�C��MC?���Q�FR�u�]�O5QƵ�u�hG�����mz�H�o����G�@��u��aϳ�(g�m� �:��3�¬o����q��7��_����_��/�_���׿zҞ>9h�^���Ϗۓ'����^�o�y�=F�[gȨaX����4��y�=z��}��wY����b��̱�͑ϖQ�\>&���q܋�~�^�W�iQG�.��6��C/�u��}�}=�9�+��0vr��Vv�׺w��a����hUu\�S����8��ώG���Z�1��,�������2�
��|�r�������Z��&|?��R�]D|�:n�;�dix�.�b2eZ,�l|�9U�d���P�0��D�A�Q�W���EM<O�v�A������ �0��C(��!A��]"�k9}����dg�̻w���P�1����'M{�E��s�����9�H��=�H���X;��͞B���h1!����1�sp|
��/�Jb���#Y����AF�h��
�=:u�г@�~�J�$M
Y�� ���<J��%�~zuu�--�0�9�����p7OۯQ/-�ŊPU5��wZ)Z�Wϡ�7�����u\��q�$6(a(����|���cq�?��;.p�{�IC·��(�=N��:;5��+7�����%LE��JO��Qۇ~T���j����l���iD��z,7�@��2}�"Ho�=�c�3{T4ŋ��2���X}$�t����j��{3ZQ�)���wx��Q5	��e'A�_�ȕ#YNt�K�v	�<�s��+WƅW^�.ʑ	4�1���'�0�<8�̩e��������ɚ��njG��.h|�c�,S�yz��g���j�L��'�P�C�i��+�a�r��#Y����20溭��x�Y�,{��+�˂a��K��4T5�JG:���)�������G~�nު�%\����.;��9Y�"��\P΅�HH�J�ʧ��O���c+�E����W�(�����y29� *,�mq~�s.�?��=@~���=�2֡�\�4�B�y�4́:�ZO�\�������E9_����Vu`���|����n���#7�Ⱥ�Cٶg���ꈗ��Hx�ڨʠ��v{�$��3ʉܰ����rʺ>��b�%�)[R�A���Ϻ�4�'�t�R&�aX�;=�����I�ۓGߴ���b��b���MO�!g�Ń�N��T:�E�r�o:
Tr���c�K."��ե�����W�{>��ɷ9��vQ"�3�X�few<�i�T��\�����������vԈ8����X�X;�줲�f�!��v��<��-S��tʸu`��	�F��c�P���|a���-W7�H���,H2�`R ����,䅆�W��P�%"�-��&��9��bZ�Ok��[����[d/e�CD��N�JW�oh����<�1)� a{h�s��9�c3�[�B%7�X\r�7��F��}�V֌.-�dѻw��7s$�ŋ���o���7�;qa�i �Kބt4��u8ݞ�C�b��n��K:��/�r{�v�х��t%�b�BRo.9p�k��$@���D�`�����v&YOv �L�)�L,�Ӵk�WF@RQ� ��&�o�h}�9�7ӡ�쨹(
8�wO0�޵��`��p��a?����N(����yq�M�[nk������[[�{����C��i�^�k�_�n��>�.���m��`=�p��0�����G/ڷ_?n���ߴ����=���r4���E��@�y�[�����f�������pQҧݔf�#yF{#�ţo�����˶K��� ��N�O��T���t�}�Q��"�ֻ/���n��P��'�E��w��A�,�L�(yx�e+�^e)�ay�!��>uaxcV_<�s�W���"���3��Q�-e7k��6��#������7� e3 �2� �l]O��$�� F(�1T7����k�a��h� ��Ynwy�˰�P�}� 2%r�&g��V�;�����)=�袱�R���'�.&=�)!��ǝ.�-�1��^1���BC+��X,������o�^�Tj}�BوU(��Նo
�X�Xx�,ù�e9H"V/���p����i��Dd#+�y�)U4���q�A���L�t�
a�UX*� q��@����1�kd��y�E'�<
k2�ArEq����{�O�z��;�8�uA3�>p�ؒ{�\���>&��Y,!�Z�b�e}e�U�jgw7ƺ��;<��`�
�s�=�%F��*{���r[^�vz�����A\����r� 
�Ą����S�7�x�U
bD�0�z�_*W�&���`�us��W��+\h��Ҹ#R�|����4��J��+@Da�4h#j�J璚�n�ۛhgF<6>KC܍,{�'f�a4���+�NѤ`�����]�a���K�n�:�=#Nʜ�ߞf�$;N�?�o��h�����遇�Q��_��%H�45������ۃ�[���۷(�Y�qpʎ�TV"T.Ç�����w0*^�w)z ]�2|�ڼx�C]���Cc�Ml�v���%���L�}s�}�ˬ���ǳD����T�)	�T�/�}'|���Z%��I��{���zT]��K�S���(U�ͷT-r�u�h�#o���N9y_���Ϩx��;y���>�G��X�1;N4H��YȀJ�YS���E i面R>SO�9�W�����}G��lٷ7�7_�l;�޴ͷ�۳�(t���'O�A�z�B�a��+dZ��=-E1��y!�]0��ԗ2�O?��3A<���݇����-������yHK�cy���[�!��{�KwE��><Գ�����w�_��{↧��c�eBN��}x�Mi��#	?�'��@��m{���Q�*1�:�r}��	���)~s&L�keWW�C���xx��U�l��Cr_��������Gf�̸�8Fҏ�H|�]�z�x�D��'L�{�S�(/��C�*�Q����.�(�v0��k�4�ԑ��a��v�;��Q��R}-��+1fl�^�z�cp������.��D{��a�N������=mF����N�½�b��Q����t7d$N&�^�*O�VFi1\�#;��>
��[�|��)k^擯2�5j���A>���?�{�}��Ӥ�샶�83=��<hO�j_}�=�x^N����C-yu����������yf�g�^���Cd��1z���V{2l�����ͷ�g��g/��7n���޼ގq��ɫ��W������׏��ܿ@��٣ ;��̴=雼���F��r��m�>���{��ы��׊�'�p�I����?���4/�L�w=����e���P�M����#!We,�v�W�`d�ܧS+�����L�]���9����^������Ӂ���#4��4|�.�7�Y�	����l�����P��L�������_��i�����z��u#��%"Lcl圥��F x��'�ۣ��R��mأ/�,�T轹��"���IU�j��5�]��,wɚ�$=�DUO˸�(��9����W�͋W���ghn��b�ݾ}�t6P�]�f.�=4��V0+ x���0�<��:k[{�ed��yA��`�b�5f�?��y��=��)*�cZ�Ƶ:p����e��Hl�<£���ѣ�����db�*��g�R��.�dz��S�V��9���Xm�;�g��;�!��"q��Bם�S��i $T�Je�pxG�2J���8%�c��z�@c��w��
����Q{��wD>��w��s��p�F+Jjqd���@w�n��_���>:�J�;�8�����������LO�F܅�
t�؜Bۇ�}���uL#N��`��@#{� �q�2��O�ۈ�!,5��X �)5V5"�C��YxCD�!��8����7y��Y�T�A�w�cb�R��#���f\�0?��,h���u��5�"�dҞB�m�	[��n��;w��G)S<���ژ�?g���f�����O�jlyL y���`9�ۻ�z�mM#��`O�/�4��d6� '�Ĵ+�eɶ�(N��5{� >��;V9�?C��t���y3
U�(�!��Ƌ���ۃ�c�8�)�6

u���D�K#����Am��Gi��Aҕ����t�����3h:unX���U�x���S��q�<��gj�nt����<��u���o^�h_|�Yֵ..,�wZE�RC��q�F�g��9�)uF���W��\ ��N�ū<�{I8�{0�
$��+��ڮ����N$�6G})��N!q���f��ߎ2.{N`��G��␦����1Y ��<�Y�Ie%ӵ�5�G�����
f��#Q�%��7mw�u��ポv�tG;�� y���w����;����Ѵ��E�z����������٣/�c�����K�_��o� ���	�A)�^�\�@�譇�(ևp"���$H��X��Ǹ���[Z�����w�����p���U�QTp �C��uV1Bʇ�[�a^��:*
�c���(�>���<o�cG	QT���{肌l'J��Ó��
�r�ΰ��َ0Ng��k�{�/�BI7�n���q|]#�N�
&1$2�<�hn�� �X����Q��D`;^�
�n�A��p=�4���,���)��\ۭܰе��1�ԥ���l£��{���v��N��G�B������Nw�s��k�w1D���¹˝��e�(��9��J����{�Ƥ�n���7ߴ_����7_�޽y�1xď"ʽ-���C��ѳ�ЅrC±���\�k$��bR9���E�u��k�5�;;f\��Hо�f�T�gYS�-٥mz��'�m�R���٫!��g�!�k u%g�l����?��}�Ž���Ǥ��q:�4m��̻��o�i������ͩe�k�..��,�h��]n����W٩(~��<�E}X�Ʀ�w���n3#�O�>mO?mϟ=ko_9M�%�/�ӧ���� �_��7�7��㈌���n������1�7���k"}[��xoۖڒ��z>ZE�%u��NI��Z�"�|��uO�	�SКzf:�m+�?�|Ƃs�fuH���Ś�� ua�zW�������$WV���>��)��ѩzxγ�����U�W�5˸��b���{C��T�����U�p���D(<	�ptXt)7�5{��*��s��αi"^X�֠i��<��
=jh���D��
+i�JEr	+'��ʳq�7\�\�h��K7��K!�z��t8�x"���T�<w�vk+��ֶ#*#����

�U���wﴏ>��}��G�M�]�T6N5?�{a��5��RF|u�).|�,Q	"��}��k�*�u{�ep���C����j�`�S�U���x�6�'��4�#p s�=m���Ƭ+t�X�-R9ѫ��b�_�lY+��a䆇�+�Iy%�(�0lz�^�a����8쩴!�fC�qw}�p��������48��~`]L��c��Y�0�@���{�
�=���DGto�v0�в��`@ (�?�*��K��Ͽ�u�Qg`l'Nz�-�z�p��8����8� �q�zx ƍ�1gJ"~#�i��9=���(��h!�.Aky4B�C~��G�T)W���.\���S��uxiF��+�V�//mJ����͗k���|[�?�Fyi�ttI�s�j����p�_�i(�iٽ*�����Jp{�b�C�9�c�o��ap��T@7H1���E�R�F8�T%�����2J>s���x��}�*�JG*��(0>?�l{�� ����˳ma޵����@�F��\�./Ei6��d�3�3?������~�3L��C�rN�ŏ^���CX��O�o�w��?�Q	z��a5�1���p����iED�:%	�:Q�8>t}�����c��oړG_��O���Q{��Q{���O�iO}�}����W۾��_����?������ڋg�b|?jo�<k�;oH{�6�8�_�Ǥ5d�J�5��k*��v�Meg����I�\�dQ��i��vR���U��v��=�]��67/o�Y I�zW�WY�>uU�ׇ����?�E���|5Z�������K�\�pY[݀��3ZS�P��j�0�;y֦j|���_@�mee��@���NלrD�?�k��A�gj)����<�#Cl��9r"� �I_\�S\;�lyY�4����m���E�����QJ�J���t��R^&?#�����z�������޶�̖8"���52��&\k�s�k�Yy�h��T܁�sE_�A�۷��SJ����P��o�'��Kx,w�WX���Q�^�F�7�x�^KIu�kɠ�Up��>����R�����æJ~���/UuX���|`<ۣ�,byyØ��6]z�������kx�9|�?����5۶���vJ;��ʣt8� !�����ZF;!��>exG�����{�}����������ū7�՛wVO����o���_���������_}۞<q;yw:ܣN4�-q,Q.��6y�� �4�"a��:��>t4��8*G(�%>����{.�~���O�!J�� �����{y�(X�T*���x�	��J��K����G����t��Uk�φw\��/z�zA�k���M���2�v�K�U�S:��
Y.��n
�p.[��LS/�g�kpV� �?�6b:!�)���G���2�JwG��u�}�FxI#���@|� �I�h���>�����_�Q��?�'��)��#a�^�-�a0��m��$�@=I�'A����U
SAn�*������y_��?��$Ja��f]A=W��7�w�o|�bF$��B!�]����z�e{�hdj:�
�A���?��x��ސސWa���'-_�?�V:iڸ�3R���%*���Hх�3�5늆խ�ݭ�Mj;>G����ö�#|s!��{���F�ì]��|BXw�2>^��.H4Z�;[m����)w�D9u4cCk�M ��~��
��h�F�Q���(�͉�T���k����t��|e��A���4>��E��^Ư�)���]ml�$&1���J�)�p��<�g. ߫���4wѴ�e�h�1�ܦ}z�C��Q�<�rCc�2�p�#n�%��|2�f(�]]��\����aF�����"V�Pi�] G�Z/�IY:�u厉��ޱ�[��=;)!�ӧ�]y%lN�y��M�Z7�������c��}d�%OiG^,�ғ7��RWUG^V%CE��d�+��k�K�xw�@1��b1ݖ<��^m;*2J����͖?�%��c]�����?��W��L7���u�/��2K�Uo�-;8��2	UE�s�X�Ƨi�3����A��C-稂NҺd�gM���Ѽ�)�;���ރ�Ͷ���l�A޼j�޼ho^=m�_=����Q{��;�������}�k�/y�}�z���w@����Ǌ�!�/�����eg~ 	G�F<hd�S�<yH��E�"���)`���uڼ[���;����meu��ώFxW��{&�+��r��z�����{�cXu?`?^�?�{�0�����m�m��8�X}m2Q�k��P��}>ǳ	Ɔ��nf�Z؇gO�~Y��3E����-y1j#@yT؈�*�؈�N^�'Uҝ��aä]�W�KeK�V�Vqmҫ>=�[z�q�w�P2�t�{�5�q5άs7�q��J���pY���zJ��I�bj�����4v��*��_��C�$�'���3\M]��C{c
�6��u�p�iA�v�S?g�2Ȏ���.�9i�Qf��!��N�IǶ1�h�l�TVkW9�,AN_;�.\W�:�����E���0M�5y����0��ڛ=�^����tpL�_vhd���t���/G%fj�2dw@�4�y���4��v
�C���!�r ����`��>���(>:D������Gg9�-Q�tqe�.����`Vy�Վr�D����84T�}���߬�T���9u<|��YѶ?�U���?iDMx֢�2�l�(ע��W��?��]�:�v_a�>{����iy4�Ee�xE~���Cc�y`Y,m�,���\ﺱ�cη�܍�j�Y=�@x�(���B`\�KRM������n�&ސN��Qx� a��R�+=#E"�j/0�܂���-�)$�A�(s�#����>����?���O��?k��?j�|�i�w�~�Ntg<�*�""�mh�%n��CA�Q��dd�_���wW�v�w�~��˄�J<U��
��r[�h�r�E\�h��J8�TC���&�J㉣<
[��&�0M�.�L��1��>?6���9ep{��WX����v<S1�Y���:(�|o20
��yj�=�h�#,�6�������+��ְ
�Ӷ�u�9՛Y[�v�����V���&�=�uBx\�Y�*鵌��@o������N�H� ��[�ڰ#-�L�� x�I�%~�IsҪ9�
J���(%0�SI����}�f�w��\��F+W<��������tL��#�'g�Q��0��O�n���U�-�CG�����<�%��'n�в�H�#_��f<��y_���]n3X��+Z�4`�(3K��iO������TD��� @�2�J�C�)����5��߇�A��`\�rY�(-_�_����]Y�k�xy�Ma���οj��\�VQ�$ňw��7o�F�H;�VT�Sv(�P�-�[>p�,�E:�8�0E6��a�W�)yP�0���鏮Es��Q,��l�N�#{��p�r1�u�v8MB��5��Q�R�*oR/o^� �P����w�����3z��Uc�C����J^���k5��Q�&@P�ENS?�ě w�������f%�2:�qtP��$*iϠ�ϸ�*H�����)�͗�57�ᘚ �s�]��-d�;����~���w(Mo���䐽�/�io�	��|������Y����Q����sn��4c�x�]��r�/C�zw$��-eKpG�0T�WVs����:�	ON(��\�%Gɂc.�+�����U��틮��N��rUy�,z��Q i�)�¼���r�R�[N���)�8��&���)�Dw����Y[@D��L��Sm}i�-�`|����+ϩwG���]�k�ҕ.#���i�y-��\ʣ�bmx1��5��B����]}��������)ys�}9x����y��E�O7�qꯛ9��X�L��޶[٤s�v�)2R�='�ֆ,�Y8
N⪔�7z��'L�I�?@
�xM[!���R�ۗjK�j����1H4Llw��N�s��08�hp�L��[άv��妝�rB�z��� �qۛvD��\`2KF\��&h�Ph>>D�o�Cl���J;[4��R��)�k��w�'�D�t*�z�m�<%.��F��L���O�,���E�N�^@�҆b$:�c
���,��@S���
�>F�#�Ǚ�vŃ����gۮ�U]y��N�y^�����Q��=\����Е���ǥ^|Ï�F�m$��R�u]����^��u��K>��Q���ϻ|�_\�R��e\%�ļl��bܙW��a.�
���y�ݑB����U���n��|��U�0]'Y03ʝ��}������n '*��5Z�WN�R x/@���y�}�ͷ���Wٝew�u1οD	"�,�;�Ǡ��/������'�~���?�Y{��(K���Z�l� �Q�3��
��x�w\�K�"檋�����e\���D�û�-^��G��ʛT~5�u���Ŀ�4ˠ*�jh��S�@���<��pOOa�|�]8�1K^��t(�0R9���T�F� C�S���W*/���"����Në�u$�s_��i��0�-��_����I��q�#�a `h����c���V�~}o7#c�P����պ����oo67�[���ݶ�V���;�o ���ux��'(U�CҴיpW,����Y�̔��i@,檱��	P>�$eW��Gb�`'���v�KӞ2�֦�60�n���j3�7�5�/a��e��m��r�w
D=�#V���z��h�K(rKW�Za�iX9z5�Q�y�OvL����v�m���;�4����/�|ax����W�%�� ~�,�qd$�!
�R¬`���|n���'>
��4�䳪[��`���F|m�A�(�vX���W5���<3]d�L�E��2p�l���<�@/�y�/ �ƫ:2�P=�n~v�-�a(L�ޅێ�cT��y�ω����M)?Ey�ptw���uU'=Fխe���*]�]e.� N(��8���MQ�3�8����Խk��G�g0b���ѐ�.�N=��
w s76�w����&�a�"??��I�F�(kk\c��Y:������h�4��}�C��vq��"�s`��p�I+�Q��Q��_8��5�-Q>���Dޝ�@��ɕ���֟�K��4ďu�᧮SҠV�Ӡ����R���\�wC���|�d�[]����:�����6�\r��%���ep����D6��rƢ�P,�-�g�����x�X�l7����"�ƶ�v�"���8m�[��:��tr���Q��͢/�� �.z�H���찛0�����t�ٖ��Zp�����{ۃ�����+�2��p�Pb.Ҩ;~��'���ڊ������L'�;��1T�euT�>"��[�2�c�
���q�FF�l[ԉl/�3�q��U� 
���{�ѷ�P�����A�Q��S~Qߡc�;�s�C�$p��\f
7F�x��p-;�j�*�.�\[��"��'F��5,�r�E�`�������P�mw�T���F�g�f����*ʏ]3f�����P��W���>x<$�cp��t���gl�����j9���%�.5N��-��ȱ6�K#JY�Ⳝ�V��� M����"|���b�C���~e����^ڭwE��NZ'��8*�v���Z�:iA�M���K��ۡ=�������!���\t毻Q��ȯJ��a�G����zƙ�D��7�88��w����C�o�6�]��G�����1I� &�
Xn�<|�����A?��@{5��+����j(���x�T�K؍�����r���_מ<y��]��A�逎T�����t[[�hwn{���������
�j�_B�.�יY\m�|�7�F�2au�yŏ���%%�G%h��陇�������P���F�������D�_=i
��٪���ّ-�MLGF���*�̮���X�u�	��ȩN�#�>[���]+ۗ�1�N1�NO���Y�p�g�����8��2���4��"M�ǰ�S�A�(t�P)>��m�������vH�n��5p�����5���n{'T7w�"^���Թ[;����"��}�ᾆ�:JN�7�>�yJ3*6�~)��MPCK��Vb(�*LM��'���6C�E�N#�M��h4<c(gQcSE�@m#K?3wc�F��Yo�S4���[ �y%��~X�o��	�<CZ����<~A�A�k��8>I�m6�x8�A��(,��2�֥Q�<�*�\˭83.����pE�8��y�qoPq�S�dZ�ѽ8�XO����Ty��oC^qM^+[ª�@kY<����d����tyX��v)^ą�ltR�|�2 �Sdq|��R�U��\'���ʄͷ�Q���e���)�M��D�`|��h�Pg(
�3iS#�\ULL�0w|.t������l�q9��2��������Fh�]�4�܉�\�LwU��oy�6��b�P�T�]ˣ�Ɇ��q����Ŷ��B۰�]`�b74���*e�p��T��e���1?�jD���s#��,���B��?oͦpQca9S���M^7�����Y�K5:��e���ز��� �ȲP���E������A��1���/�լ��ʈZ��a\��.RG�15��	wω7p&]�Â�h��;��,x\��j�+������� ���TM�3�1���J�|C8��,) memz�I_��[v(5o2O�L��ȶJY��"r-a��1l�@#��݃0HO{�~��β�J/��9��`�էb�9�/_�h/�?o/^��Z+�ގ:��Mx޽}��ʖ�M��
�#m�ʬ�=pi����w:/֡����W7c�
�ߓ�`�<e���:Ix�^� K1�r��x��c�O��0���h���`���o�q�#�)���ȏ#�5�]�r8]ؑ-�\��)�1t��)�{G�g�CK�s�<�+���E��GR�R��#2�:�?�)}�i�N��F0c��^����v�DN9Z��#�����F�G<�ѯ���ACK�s4�YJe��O��{X�e��Qf��h-C��2rŽ���m :�������n��kp^�����K(C`e_p�:��w^;n+m�E/���4C�q��t}q�^ٖߏ��9\��m�z��[����廻��n/�eY$���؇��dy�?Ҽ
@�,�$t�9zu="/Tz����-�!]�UE�4�]8 �̸k�_��j�����_���y�ER0�$�픅ӡ� �`<��i�hH�����92��I 5}��k���3$|Q�(��
�^ȯ�ǯ��z(7���A���t����6���W����6��|��T=��i�t*U���9���h8�H���ʢ
��m `t�x%�ț�uV�06v���v�|��|�v<]#'��wmwg�����u��}
���x��|��V�t�G��n��������g��v��v�w����wӛWʌ�Fp#�F��� s���;n�����Fik#����9'=�0���}���;��04�G�MX�����M~* �h=�cg�[�G�4B�h�Q)q����\=�\��f��~��P���uIc�LO�wW"����U����mv�F��g6hHn�����O��	l�g�a&��!e��uK�5<�s+|#�����޼��.�t�xi:����|��ǁ�G.����3�}�/����T;*��+?�k�]�zK+Lߗ�ք'2h��2�o��0��RQ0[a�>�@N}�V�FSX�i�� ��)/i��]��w��P)ܩй��;4�5�����y��,����mZ�?7]��9��T����M�*.�ĘY����ww)�F7��Y_u��y�T�xO�=d}UބG�F$)���L���
?��R'��O'�҄�g1��%CJ�aǓӎ�:�G?��h�蔈{{G�ͻ���՛������٫�����������f{�f���m���u}�ny��ce�A�}�i���o�v2��Nm��n�S��,ƒ;NcNP��U�P�Q��Y�
:���<�mn��y(���q�C��S���n��ҕt:jo~��˧��븘l����G��u��+�t� �knf��)�Y��c=���
����%����q�NQ�YG����
Fm>8u{|G��T��5Хmy_ݢ�s�t;lepϟ��#�v��h�aSL�
<N}8K��AI|�<%$�HG�)��<�	�Oĕ���mul�$�g`il)c4�]��ٳ�C���7����ޣ$^bd���܌�e�)W ��'2цKX7~�*�� �rN!���V�ӂ��K��(唩�r�z���_�[��3Yb�vy�.q�:�M�Ͻ��d�/#�¹����y��٢�:HY�j�L:o൩Ye�4~&rbfa�M�-f���L�9h���eMç�x6�B�h+�լ-q]���4��Ye��Q$��9FPFI�{Hy�b�aT�X�o��k���G�F�W�㈕y�o�.>uJ�¯�cA��}�)��R4��C�}��t�s��K�Zq#����ᥑ�/����KLo��jR�&���w��p?t����z7����\�*9h-媲��:ߧ#eR]����o�l�����r*��3��7z�wy}��𾬼��K��h�!�P������_���/�������=y�m���]�Q:E�d$��1�^�:!��H��w\��R�nx���A�h���8a��2+�z��b�����l�o�Ziy�ҟ�K��G�V�k�0��1x��Eé�嶻�g����F�g�P1MS��"��h�4@%rG��]Oض7�p�j���q���i�N$j�zv\��
�#am��׉#Y"{Xʘ��� tE�iOs�@
OmS��ɹ&m�#�:��w\��Ȕ�`�N� �w<�ct��˧��$�ْ�2��Q��=¨Ұ<�~�]��y������N���k��h���TA�ǘߋ��4V���r�Q�0�W=�*��K�D�wۺr��}�N{�EW�5�j.�|�?{�y� �lI�F����;�Z;����(��׵qwE�H�h����B�B���6���~�w���,`���o�)���^z�Y��y`\�i�(q�c�|�^)`������IGA
�Wxs�p�����\��Kw����(C�6��kh���E�ėܩ�Jl`����K����5 +|d��&�RE� u�eeWon	ͣF:�!��H;�2e��E���nW��D��m��N�_Cq��g1�ڒ[�#�f10�ә~���*��Occ�4j�VS�IW}����u=�%��`B1|��^*ߢ}饛���?���Q�u$K%��k)]�z��Oe�D�ӻ0B<@tn	�
��]1!`T�kٖک����Hו6yX�F�퍾66C⨑F���tZ��ጝ���������Sm�99�h����9@�"�4�4���N�V�*4�q|�������(�n�}��� ���v�EG��Iе�oz�{h�р�� ��C]���+��wy�[&�օ�λܿ�Y�!r��W^zt��/T<�U�Tm*cO������&g2��Y+++˙
�z;lX�E��`f�w4���M;�EU>$���Ox䈆��%��.z�;ro�#��8�.k�[KZ򥾕������6�*ePf���k�e�2�Q^�%]�V��6�'� ln6a��wn��'�Hl:5���Tp�O}H���N���Uة�x�c�)�,4k���
c�W��z�/F|�p!ۨ%��9|�1Ky\\��8�)|��M� �O���oh�i�ś�J�X#�Z��-@+�w�ĸ����4��#�̩��C���B�];z���"ӄ_`�4Op�b��i�dV�����:�A�8����u�1$n$x�-��+&�q�z�ތs�{��>�:p򮌭�n�etRc�khY�����2wإ���V���CK��F5L�WȚ����{���n�X�m�|��Y�uw��i�Fpy_/�?8a��g:��{?-����4�����7ߥ3���*�^��g8�c��o����������u񳗛��.)�!�+2�ev��iF'�@�3�O�YyG�ԛ��i�TŔb�y��������l��u4�Tһ���
�ǳ�V <P�<�qJ�/+bWМ:�I41��'C��ݽ���y��m��=y�Ee�v��D(��oj�Z�B�k	��w8	�����*B�)M����e�a^ޏ��� �K!+�S�L�P1���FAE0�hкum]�y.�0MӖ	�&�lP$:�$�ދ*G~��K�z�T��A �ô���q�b��VF�lP�9������9�:=e
q)H��F{�r����&#;�A��]8욚�o߶7o<�ͩ����ꚤӳq��8��u�6]���!�s�r��0��i,�#�;p�wr�$�B#��fSsО[�����t:��%���AɈ���
Wo���i���pp!�\
���撄4e�8DmO�S���0MҨL�Ш8���(NM/�!��h8¨�N޳N��]wO��s~zz��i�+I2e"\Ѻ�cᄫ����H�*H}����H}2���4��
/��bt�뮩��Ё^~+�����|{��Kի�Y*���&�#e���,��U��v��Ͷ��E�z0�["�fk��ݞY�7��>L�Bt�䁴�w��>ߧ|�+������M�,d��9�l9l���R������<$��
9fꚖ�嵶�q�-�nP��o��b���c��`ǿ��<�:�G/t���^X����~�c�5��<�>��<�{#�����������}󢹥�9
��0�2PN�R�1�y��J
�%���9���ѡY�_��|�g�yX���휈��Ȣ{;u��ն�>׮gk�U�_�@��su�� _[����n$���u�`84�Tp��8����L'�p��q'5�I�;eh�5%3�/h�3�����+��Ս.Tg�mV�~>|�4ո�v�:��a�̌qAR`z��VWt�}��|z�:L5�%҂>a��3��p��R���^���݌Fjt%=ӗw�L;��͝�������}��!���|e�K���w��4�i"~|"pl���z@�-1��� ہ��G��`0`�OY2%��M[i��&�T����!<m�G�C�keNr�ܰ�xa~Z����>Q:vʿ�}��b}m-��We�F���޹�n���͛9��%��n��3��[[�ѧ�[LJj��ݪ'E��۲���S���1�o�������Ae$Y�Y܈7u?;�(Kխ2���ND��Ȼl�E���T�$���	�R��F�XYZjwo]own���GH������כ���뭌2� ��̴��vD���4�Evh��7�/�U��*8�s߷V��Đ�V�p��R��|�E�N�7���D^�$yi��7}��۸z��U_�&���M��ni���u v�Sqm��)�����I��I�ڦ�j�4*��h�b*���`�:� �|��G��x�r��p#c��T�<_���p��k���/{���H y��^닗�Q���$��n٤?��]�J�sfޝ�]f1�6F�8}��F�y�F[_]��'iîYo������	����I�xR��t���~'Hb+l�,�d�!G�P�!�_ˌ*�2�ƚ���0��1������.��x��5�F��59e���>:��J�vd;�st�r���}���q�w�5;N5��
 ��TF�/ї75���Cȹ����I.ɏ�|K|��R��(�F/F�r\y9\�;�Hp]�&>�`H�?���(�S��38�<��U)������1�������k�@�����B?ӽڣ����;�3�XeQ�*%���Rw*�
N�/�1��P<�,� k�� �,��e�Ɓ��9J�.�w�G�6�����[�ҵƃ�?�a|���;adm��<c��Q1�����߇��|.G�N��%�d(�|�H��� ]���c_#P��ʱ?���q�L����K^F���|P��J���� ����S<Ә9]�s�<�#�Cb�i<yࣾz�5
Q4	�i�n�c��l�a'��y(D"8S��%E�x�"̡q�<�y;PB��"%b}�>�(shFz�>���z����;kRa�j�R�"�訦F�v#��L�w�-�^h2Z�̩xp﷌��`:k+�˛��p|uEa�~�"a\O���k��͌t� �N�	���'��?���E���Z��\<e�:��C��)�ܬJ�|����V���<���IEMY�ڂ�I�\'���U��G�D��K���P��%�ux���\ç8���>w)�4D^f�F�O�?:p�%F���m����a�n����� g��x�!X�����TQw��|z`���/����
8WNȳs�mqq-��~C���v�ƭv�
��{�֝{��������n�^�n�	�����]�8[XZ��ښ\E�]�((F��:0�U��Yy:�!5=k'�YG�S{�]_��-,��(�SQ�]E��4����V8�p-�puUq�|����&.��z�����)�
*�|x��w�Wm��s��>x�\�Ϣ�n��v�����p뙀}��QÃu咴_y�f?*���Ȟ���]{���v��H�sڭ��gv�#����pV�
ra�6?���E/��S:�0�Ż����8z�5Mȟ����,�^lSm���rg#g��l�P�Cy'�bt�Q�G}��޽߈���ҨҸz��Q����dT��'r*x�C��=>���A�f ]� Mݐ�HN�����2�T�����Ω\`vj�r�8v4U�hd�zٙ��Cئ����t4^N��2�5�s����v����.@Gҿ��%(����ͻt�-�;�R�R��)����!}���]�Lҵ���Wy'����p�Ǣ��O��봮���Y�Sv���r����IOY*=�ҐN�+�ZI>?��5P����V��{Gz!%>�n9�\�S��p�)�NA����M;�u�2�>�dn}߿~��:������0��3���-~��䫔/_*���;�7� ?�xN��G�Q�:<��,���xFy�f��ϣtfB?�ಥ�zS�a�?�YO_�m�_m�m���6(�*�"O`Ul=�$F��4����KEt�$L�e+aY����O�^�Q\Y�ј_���bYp��j>n��������������ѓ(�O��l/߼lG0�����;W]D_Ui��!�m�?�Ⱥ �����59;�(�ɒM%Ɂĭ��"ˀ��|xg��R#+��}5x��IJ����ʗ�Jr��{᝛����g�Js���FE���k��(꒷�I�
�-�:���Gp���i�a� ��,b�/-��L��������V�I��B_�і��ڲ'��	������gQxHG�P��:0Te��)��aίA��eFzrҊ�2_���C��zh�g�!m%�Q�e7܎]�3��x8&��ã��x�v+B� �����y��0OBc��)�p��5�0����?7����=h#�X6��4�jX"�g\�*;�(��=�'�Ӕ�!�b�4>�˚����FF{����?E� ���� Ҽv�(e��^k4����EH�Fs�P&�Z��i�i��Q�\����<~��àݞ�w:�B�/�ݐ���_�y��x�$�҃�p�i�k�O	.�z�~�HϠ��>r����6��*���,z�DຎO�<�>�Z��gz� ��P�TpI�N�;� i9��~��ܸ}�ݹ{E�F�%9�%���x�����՛�c��R�B%D:L����B�v�(y�R��n>-��������J�S�g�-S��ȴ;+�m�o�(i㮱�zp���ru���j�s�f���'Rɨjh����Rz-�"��\@\��U�l�� ��e�3��(�*��{)\,�#�B,��'�1�3���wo���g�|o�M��	��q��F?J,��?���U��Yo������qۂO�0�U�<�{�d�G#hC���v�at��öz�N[Z��Q�%��ŕ�6�l���i��9��Ц���mBܵ��)����6�r��w�|fM�����7ﶍ[��ƍ�my�f�u�N��8RF8�f��s6���).hG���8����7�O��q��z ����@:���J�9`�*{t򐼦B���J�o�?��G|o�.]���28�]୴C}��Ç{mk���s�����n��z��dl�5�5NƯ9�+)���H<CQ�v���)j㼟!.t&_��D�yB ܺ��Q�e��J[hK�T�rz�F��IuNp�o��5�2m�B���v�)�<(�����CǇ\��/��-�,i���6[3v��y�ċ���Ў�)�ې?}�4#So^�l�{d㒀m�{pzq���M{��e���/�W_������Y�j���YF�qQ�1�)�(^�i䒀�3E�����dV�u�*O��q�F�������ǥS��>�"�wV:�.�v�m�m�-����^;Ǐc�+���i�[��n>�������yC��z:�au�6�v�+d��W���|���o)�>1��=W��6T�m�-'�G�X���Ë��z0@XhH:J<��0�0;�
^���&5�ɁV"7��L��.���֥.��i/�9�ʽU�چ�_���|��N�jE�<�B�:0Ե����,����4�l��.Ǩ�1a:�)��u�AޫÕqm{D��,\ʚx!P_�~{�*��<�ʻ�',?�ő�w�s�w�xupB���W'��IE��N���t� \C�PF�+"Tq*�#7��|�9@1��������(�-�[�hK�q��������?�n�=y��={�.lND��ȲV�@(�9p��ʝ#Y6��dY9U�18��	� ���<B%���]g�r�qQ*4�Hd�*]��E�o߼i�6o߽JźɅ�~����[�^p�#4$�ps`Q��@�~� F�=j;�\�Q�����z�>���!�z�[�����o0I�eX����>�zmK�^*'�gF����;�"P-O�X\�\T����C*I!�����^w�r1��W	�����myy���jX-~����Z]mk(5�K�W���_0.������J��9�5��6�گm�;6�!�����SO�.2y�G8�%�32q\�)��b��Cx�#�F'c*��t�E�bd�}��C����mD�E,kHL�c��c�*�)|5�ݪ�.P�il�4��(��e���tZ�l���N�]%�fy0��)c<��H�I>|�l ����Jq�u�/��.�;%8Bx�(�*�y'.b�&^5�YS_�ȼTRw���U�+'\.V_e���
��PaH�J��J/
�t �2��f��W����mw峷У2u8�w�a��9"�$[��x���v��W� �$\�?��������.���Hw�t����/jG�w�2ꙩ5X�4�TI�x�FQe^���[f�����9�l�99�i<������t[Aip!��rI7�٧�'�?����FD�7k&X2_���葯�8ɥ^�N8��������-y�Ԍq�_I�4�g��Q��7m�-�%���Oʬ�-�j���	���J�I��]c�c<ogo���97�XY[��qtJ�
#����7������kX�2
&;�IA� aZZ�UO}�C^�!��b�����f�a��B�[A^��9�г�j��ŅUd�Ӌ��.�ۘiU^�h�݉p|z��-̵d���Q��4GG��%��hP�7��,��S�.�!��*�?���/����KW\Z9����kh1޽h/_>���i�t���P��΃+��1�P`0�4��Z�X�E�5NN�AG�`�]��)ʥ��
� j��Cg��A��#2�}��*Xƃ�L��}o7x̣H�a򬲪���y���]��F���9e�|�;�._��l~�$w^��z�^a\�ƿ������?�}���p ���D��r[w;�i�҆|	��i�\��g�%��3��^w�}� 5��>ubg��f2�e���:$���#[���q7�R|��(��<H9b���:�ϝ>�\Ȇ&�M�[����v}c�}���v���ɬ��R��p��m?y֞�|��W�k�\[��[X͛_�H[泰�L�N���g�R�z�}1�u�:�=
�-U�ֳ���#�J���r>��e����x+��e��kn����]������͑�Q9�^m��#�x��u�'�C�g�����,.����?�z�����4�=7��w���\�gn�W^�W���G����*�S3Z�sҡ<�q�W��(sS����^��L���w����Y����e�@�^�	��x�FN�(V��i%M
d�x�p_P>�H����w������r4KEfA�����g9O�/���M{Ƴ�v����*_�UD�+�jyz	OB�o����\�p5���!_���˼#��+^zCno�=�~{�x����HOЅs1,��u� � a���n�w��Ƃ��԰�Y�;�~��@��;�c���߸��6P�W��*�V4�P"�=������������0�mG ��Z���(+Kd�P)��%��*}�ՠX���2��a�~�qt�����E�k���=7�p1,~��S�3�l?	]y&�[�bT��x>��щs�	��pTõ�*b��{���A e�:^=(a�VZ�U�W��i�8�.�k���Z��}���	Ң`Ԣ���߳5�S"�4~�0�ή���|�<�.�'�������s7��sP�Cb���G<�e����?p)�D}�W��5����0��h�ʍ�@T�(c:M��)��^mF�t%����~�?*��²�t���l��EƎ�cٸ��yk�� ����*��f�R`�$����� �ۖ�Q���&G��v�P#�-~��/�	�߱G,ds��ls|p@�"���L�Y�˷�`��T�U�7�k�K��y������V I	۸��ׅ���RE4��M?� A�a�H�|v�]�,G��M�hY��:�݇�~�|�i���΃��Ɲ{m���5��֦	;�Q��6���P�R�Ge��:	��[-#�I������P�:1�۹�j�͕1��tCK�:�q��A�s���'?k�������=��s`���qd��	wƝ�j�V+r*�P�ze�=ޒ(��$�8�h�Ƹ�<�i�u����j���p�]�U�w]xO��K#�x���cK~2|�#߉�wGw��M��0Ң�81q��'rN�쌝-T#��q�iOCFM��J'���U<
��zVgp���)��/�%*\~n}W8����k�囊l�Mǁ�}�N�c��m�hKK���]�*ۆb��i�/f���asw�~�ݷ�7���}���َٝhq{U)��"��E��RТy�Pe�r��C����4�[X���8�.�u"~v��GQ́�h���U���zȬI��;���r����tB �̴8�9zZ�瑻�O>ƹ��:t꿻uR���S�1ϱt�*�����*b�=>�?���Q d��vf��V���M%���2��eG�	�|�.@x�a�G���S�����UWq4OmK�;���h�=�H'ue�\q�ݲ�;�q=eK�q~��.s�{�QZ��ΈE��!�R��U:��`�g�������v��^8�M��q
-:V���_����Qxڐ��t6�p�,��|�S���/,��U7|>���?~|�����Rё�V�*��xGx6O!5\z鈗Q�S�܌�-�߾����S�G���O��ׯ�d݌��~yR ^��[�����r)I�W��f�8G�fѻ� 9�W�pQq��r���]O�V�cS4�Q-� �tlHI�+���.�����[��~�-�m�����.Z���
{
?�F}o�� �n,1kϩS
��]�T����ɩ6�-�η�9�5G�0�V�Zw}-S�s�,k�kZ�J��i�<;BQ�(�\_gcⴂ���T���i�&�cx�ц���=h`gg?~o��6��j�@a�z��t|���ܖa�X\�ZL]f�UwlT��a5�rr{�Y1�d�"���K�ݺ
�wW�7�x�sh�7ý��i(4����y��؎xl.²Q#C�r�O�1�Χ(�d�)�鉣�:-�rfwC�F]�P���QC`�-�49���N����e�'���),�F5\��(@�b~��@?�B��3%��r(�G>ǥ�������
͊����ȬiK�;�����"��-�O*4vDi�BRJW~��2��C�����b�L^����/G�	�1�n��y��cҷ��V7p�ΝbR�x���"��;�C�H���z�����}.��F�c�tz��8C����=�%�/9
���{^����L��Kv.9J��Lr����buz�Gz���m\o�>��}�����~�>�z�O��;�����6���!3�e�� vX��ï��ѹP�.Ȓn4��p�������.}�M�dN"���77��U��Q��g������>����އ�����x��AoS��8�6���f0�ww�}��M��ݎ�%�L��Ѥ���|zP�xѐ#�Z���*������j��?�Ǔdx9���w���#���4�(!��=�N#�K.g:Ʀt#�s��F6|��90�QP�r<���wҘ~��7�W#I�z}c)^ʐ�x�n��o�oyi=�u�}��k�� *k�|�ѳ���G���ӟ��=|���W���s�C�Z�h���#]�"��I\�Z-��ZZ�D�'��f�2�rmM��H�w�"Ũz���������� ��=>�م#���*���Y��f$F�-����9�v*9ҙͰ��%�EƑՄG# �G������킗w[���ֻ���C{��~v)%�d�<t�.��%T84�  ��IDATqlzn�_}�-�!?����w�IO�+p׶콽�tF9i���_����6<��X�O��9��!^��j'�0s%�ZrK�:ǩ�����e�t��⦾H�c�����U�ߣ���v��~,�{��X���W�$~�g���q�{_.�?�ų:�m���U�ը��ͦ����G�Q�<�Uz�ͨ|9I�*"@cjp�x�w�WE���p��]�h�?ËT�A��P��u:V���9�N-� b�ʠ"�-�3��}�=��Q��+{r�k�0�j)dEZ�*1t�vv�˫a�s���G9q9���_�7_G��#���v��m��4�ͨ� T*�J[ao/���.w��)�=p*��.��n�w�sʤʁ��MO׎U��A}���4<����Q;��S��5�4����W�2uqu��.��:�НH���9h��ϝ!s�(vm`�4F����rS7ژ�:3���nZ0I�'��1���|��C��r�=66�x ����F���J��``�4A��,�
:gݹ�2��G�
a|jp)�:�� (@׿*����ZN}Kb��f5FT�*o��Ե�#{�a���2��[�В�ar#O�����U�2e��X��?��pvV�h5H���%5�2]}��O9��J��eY.�v����,s�-�������[�o)#��IEhP�ڡ%{J퉌�BL�}�Gvx�R� 1�K�R���_e��.�#*41�xo�{{�;�>h/{���w�y[Nm�fʧQ��U�v�ቋ6��83��Pp����a?�a�*:3V>w����v��|��Q�
��?ěa�v��
�hT$
*A�k�нV��g&����(���y�_PQ�8����VF�Ww�;F�r
�S9U�����4=�˵US�?w��7�g�֝�W�ۭ{��Ï>n~�)F�G�ƝY���f � R���ȕ�����W���X�g�_��q�5�b\9�`xF��vyu����ep��N1d���/n����mf�f[�q�ݺ�1� ����� �u�ö܋kmc��}w���x��=�*�v*�`éG�R#�����Nc]#��aT;������3��u?r���]�@/?j�ȏ������@G��㧃�!�w
���G{��~�8��8ks�����|C巉����E��(T�t
�B��ŷ̊ ��:��'��r���5��_x�jq]�m\��w��1ʈ/ck�+<���ҾƠ�?x��}��'K�?D�l"��{X_|�Y��O�hc��v
캳LV����ǲ;�;��'�|�>�^�y#k�2H^�*p]��h�ޑ~��%�(Ep�b�/]}W��S��6�6z%��'��%�=�u��� n4J�ugGȵ�t,�i`q�Զ!��
����-�����.A-��X'�͛������������[����SE�D����i��`[^�t歄{yG�x_R�zU�UR��羦
*���5�2�ԫ�U�B�E��#�^G��&=p^�1̜�t��:J?^��W����.����M��:����/��r_�H�AO<��;fĝ���\eݐ}`�ƣ-]���7y�|n�H���8�yN�hp�VH#h��b��x����zA��D�)憋����5�H;|�?�����l�G��d�w����D������rõ2�BZ���(�FE�� ��Xgh���9�!�����L��.E���I�WG5�*Ѻ�K��t��U�-���t��� .ar�ӡTJ�ϲ��.
���k���U]��d�2EI����+��;7W�d�������Gޅ�(^1f�!i��y���:�m��v�2�[/vpF؃7^�q+�C��(d0�A�4~�W���:�*\�:&���}��(D��!+�Du�+��}�SOc�`
�嫸��)�H��lݚ�\5Ν'��E���
�5��~~��	
,i�A��aY����+����w͊�6i\x�50SO�M����� ��1��0؎ ��'d��	�y�sk��/��`���*lUvK�j�f��k݇�X�僐 �4�4�e�ԕ�>�|��.*xOh��\bD��lRC�i���]����b���<�@�~�Pa.��G�����Cۖ	�����t��U���ǹ�. wj�d6�pm�
�<�m�3��z���NM���a�������;
\�������q��.���L�y��eF����o �֙�G��{#Z��"��St���-Ͷ��X��ܺ�];;�����z7F�r&
0������bhR٩ˆ��o�)M4&�eX�U�z]��`�������0�H��YiC�)�ᆰ@���j1�4)���������������v��C�"�i7,�mnt��v�h\ihy���w۝�;�>l��=n)
���1�4���)�GXe>���-�pR��8��F�Ѱ¿�Q���ÔK���k�ِ��U?�S}O[�,��SVR��'x��Ņ��N���޼l���Y�j��4O�*x���-,䬌�Σ����6�XWe���P�mĽ7�2�2R|�'������������v��vU��o�d�%��J:�-�m�<�N�zv�#�%��iH��k�|�d�s+FEw0*ޭ��j�r��qy��\�o������I}�EB١ ����s�>���?F�,�P)��s���Hս���Q��w߷�������_��EF�n޺��uҞ�'���3u������숪����]d��G��H۔]:��5Y��;:�t����Кt;��1@S_�����U]�YH�߮Ê���B�Y�A��a�+ω�K�^�kT9�C=�"79��}��dbd��wn�����}�كv��z����1���n�����_~�~�������� ��-���A۶�3h /�b�^S��-�z�@�u(������B[��<�w�2#�ґ������b��6��4H���%ZCI}���W��L�c|��_�NL�d��U�5�l���q@��v��
Q�!�K�t1�I_/.�Q�<;	lk���h��W�ګ����9��\�&��VEn�Q��:��/�V���{G��Y�RM��e��ޚ����mai����Bn��=tD;�]7�17�⻼�QuP�����ǿ�sw`{��F��	id�<��K1�"�9Yx�y��5��ڧ���
=EPVl*&L
"��.�T!�bk/��ѵ� �J�kl�3����'De˳d�rP����찵��� H���.�&$.Eh�F��~�3�v��Y�X�`Y���������r	��%a��⨻0�_�^����C��4��a2Laj��r@�"9~
E��ŏ����0)�'}Q�h&$a���껼��#<�\�xI�^����W�#z�����?_���D����r^E � ;�5�0�|�T��R�]��1̢��[���Fɱ����Uc�ú��*l�X��}p:�1q]����`�C��OL���<\�C�@���@¼<8X�d$(����q����JU�B���D0<u��jgFz_)dM�{*��E<O�:�l8�ȟE�O�P*���+e��/ �{���������ˀ#wy_�*0t�R�������é.Yu4�yA:��S�B�0�F���i���N�4�6��k�t�2��tp ����\�\��skӨ�bT���s��7�_���=����f���==�M�2#�"?��R�hT!����c�g��/M�1�����c�XGm�r#"Q\�S���D.��<��
No��$Zq�8�<�_�2s�:a��\����X7��GO:|�l�R��~ޗ�!U��kf�f�v���W��K���Y���"�id����h^�T�=��39�j㺻��o�Z>O�.B3(r1�,������0*�0=��>��5�0����2�<Uf�,�.���Ub�_�*������4mO(�r��y_�Ig�J�#ȓ��:"C%I��N �er7B;y�P�b(Xf�xŢ�Z$���mX�Y����`���B��ߋ��
G�,TB���ݝ�(�/���+x�-b08�-�?�TF�AZRQ�'��5���Z�!�|p�^��?8rc�9|ސ�v|alEP��3��������L��t�+#݁Y��ȉ�>�V7 �*�7��/�`�0j`!�ҡb'��
���&�Q�l�
:�ϳ�T��~�o��ۓ��e}u�X�Ћ8s�����v���X�o�?9'���'Y��4�Uz�����N�s��`�˳��ұ0�Iͅ����%Ҭ���������*����-�Kg�Xnha��}ڰ3o��@n�%|k��o���u��fڽ�w��������(����5F��߿h_~�=��c�w��zlh�B��N�/� wS�����RՍX�@��/x�)�y�d�S�O�1����x��D�i%�KK�)�T<���Q)G���2��3���^#��*,u:�
��J����YR���I�i����_�9'�5�N�d�8l�ď��N�|�h��&��2s�=�r-Y��7d�+����^��0q�`��e�y�����+���M�,q�}}Ww�;�">'��r���������� �����t�{w���R=!=b������/�z����m�È���ҋ.�̊J�F�FS����@z�$��K�B�"S����L�C�]o,S�E O�
����?�p��^�8��i�햱k�򭶾����8ٓgx���D�1�#�lﹽ{� r��(b���j�:,]	.��s�=߹y�Ȫu�_.y.���U�;|��N|p�1\�%nƖA����I���=�2�:�+D�s:5b�����{)�~�@u����h�9��&$
`�N�3-�Y�`�@A�"�
f�hQ��2h<E/ՈV��H&�Ռ����\����g{z31�r�M5�S0�pQa�,���յF�7��V�X`TaQ�S����>�۴���X��k,���T<<ߦf�g$ht�h~��g,�Oy�p���'t�/��1螪}ӫ��S1����W�W|�6%�s��/|��IOw��4c���w�K�W�Y�h��*?����[/k�����H�Y�6ZY%��'ԩ(6BF�r����0���rZ��rgG�\�ptP��$)�l<�8��8����$�o��4C<GI=�hmu5�qT�����O0����Q�Ĩ�R�� �H+g�z@܈�7|����"�4��S�N��n˓mmq�-�Ҡ"��sW-�`<M*�\����\�(�x����&+�L}��ț����7���� ��p�UIܺ�5�t/6#ϹZz��*$�%Q�e�po��{��h(��oQL��o�e��!7����(���+���������{my�F��_�/g�چP�#�S~䎰��U@�E�Q"�L��ӓ�J���w�,�'$�ʫ׍��:<�2��x*��xGz)\�lGʫwٝ5��H���HE�xEM�r,c�n�!�'�5 �[]���s?��w��g]�J�����N��~Ӷ�^��rZ�2�Q�sq��t�(-��J��{)�v�z���'�,�}t�Q��S��xW�-��jsT���LV���P��V�p#��<UNX_I��@�e���}��a�
�h���YUg K������~�$�mw�?�?�6[�����)��{�i�t�.���n�r���[+��d6{��Q{��qvBu�e��4�	���;��vZ��]�F|�����Ա��;�Q'mKw�G,�vy��	:�9z���N��]hw��"ݞ���#�����K�iM�p����������{�?����=Hک����>������#y;Ќg˩ש��L�,(CKޢĔ�db�_n�⡰¢��h���6I�r�P��S0V[+R���M�2��A:���y�Ε��o�*�V�2�WF�	��(y��S#�<��,��ʔ�-5Hqgg�cػ�3BLKK#V��,f�Xm��@F����u��<[ש/�u7<��
���:���M��;x�����ܡ��@�߼NFḦޣ�\T{��0I�F��M��Ъ#9������M��t�ކ5���7\�P'���M#+#Y�1�<��	E�{YD��P�ޑ�o�tA�� ؅�O�~�0)\sߟ�����J���Y!V��#���Uo�I�C؄䡁e�ʰ�QV�r���׳����7P����>�	��g:"���5O�ߦ�[��mg�Z�?��,{�F��֍,�-dRB�5���檑c���Ί����ﵫ��䭟�gaW�fx�J�W�O���(����4B�R"��'^܋C�ʌ=Y��ѬA���rӮ�F`h����\ݥ��Iu��V{�)�V��W8	�� ��C�2c��*�5�<E&����UZr�@�~a~�-iPa�,h`���id�>��B\\��7{c���a�t�۱�9P�n䠢u~1�|}��;�1V��@!�	B��iP#����R�X#�`�	��I���T�XVY�Ey��Z���2�����z���C�+����OOd6��]��E؏���0��2���=�Vq�5�DHã��4p*���
��_�z�CW��gY���/̟Gmc-ߙ�q�(nM���W��d��4(����Э��]ҝH�R�ćN���:�� d�_y���1��,�t�����(�N�y��i�:��<�M��)�;�t�[���#y�W/e������t�bsm}q�-�S.���vz�Ă��*#+���ف�;��u�Q��;; l09 e�H��un/ݨ�.]x���է��5'>��*W����S�f쵽�����s�W�p�:E%F�N	Þ�)�xq�FsJ�����ZX�/�pq{�񴄤�ڤh���rk�Dq��FlV��G�Sq:�ɵ�yx֍��/��Η���l��r��t'��. w��uh(��`�N�WG�R��Pae���d�g0��ݦ=�B6;���C����i�os���vt{��K���P@��c\��i���k���eƨU;a�4��z���q�C��C�'�>���;5��ed���.���(w�qv�Ca�I;k9BɈ�e�uT���,%L�]+Y�g�K��v�?�t}�s�;�i�購!�ʹ����߼~���|��F�i<mom�;��C�� �ۣ�*��y���k�|�mF�mÝ�!�Y�~���*��˱�v��'���4�AN���x#��S� N���Y�
V/�'�s���EY��7,c��(q�T73q��8��C���n�������<�w�}��'���ն�<�v�5�[ۇ�����/ڳ���Ӹ�܍i4�\[)�A����2`���Sg�-H�<2)u���[*=hXe�ᣮˠ1��Ĥ?iJ2m�1�}����F�P�@NE�%�*%�$Z|^��d��#�齭�i�0�ŕ��[w�{��Ҳ�Б�m��G�	Io�Ȏ��.�l�Zm �B͹��&{�,<#��׳�q&�Bvw���[^����b�>(0�	>��j�A����mk�t`mH�,d����������M���lT�8�}�F�{�v�X[�D1���Y/�l^Yc�d �Dp	��F�h����]G�D,�FR����}1��x�qW�S"�<N�G�(�����W��@!׊V���<����j�~}�ݼ�$K��{*%��6�)����`DX�-����:��R�������x���2�pidU�r��kc���g7�$���_z����p��%��BOC:���I���q2�:bV���4�����(��ΎC�x~���޽�F��"��i�7�����Z�tp(�+���1���ᷞRvJ'��/�pB/G�{�S�(:���,w#�/̹+�|F쭳w��j37��m>ȡn�r�S���(7�r<� ���j��l�>G@TR��<>#X�Y1.��T�0+��X� ��H/��9W8[����w�\�y`���ױ���n��$ʬ�#J�H$G�ǣ��f; ��w�95��ۙoչ �5h�.�[Q�vǎm�
�����(q��ףXM��7q�S|��P��m�U�
@M�_�h��`0��턁r���,\�N��x�M�*�Jy�r�#���45M���_�_cLW?�*c��W)(�����GɚT���%8�MeC!4w�A�T��h�葳Y�Xըu	U���Me�aU�'u��:���x�.��¥^����f�ݝ�9�!�����L�ҭ�������;ajC�#�7�����miq�-N��IT��[r�Ǻ��-�o.3R�!��9�(�V))<�i�d�$�������LڢS���m�C���W5c���K�U�
���d�&~v|��w�
���.msF�J����v�L���"�����mq����'�VJ�N�΍Q#辰�nj�~�)�~��)b��Ifzkm����Jo���v�6�i�7t���yR:���wڋ����˨��)#峭�����4���#�Y=޹$VW������n{��U{��U�e�ʚK3ؖ�U�n�����}��I;�>�a�ussM۟�dy�N;?;L?P�2�
N�Nw+�UZS��ヤW0�O�w,�.�ٻ��  `tp���e��w2�^#q��	�f&C<��e�����qxY-3��e�\�-�m�l��a�	%�Q���9ҧ�^Nk> %o/@��r�hX����
����G�ly)�>
�����y�&@�`}��/۳�O�Y����GWoxR�i�6ү,{��o��ԡ�[�Ħ���e�y]�F�3A���q�`9�%�U�S�*��r&�TP�_�w�=���tV�.N�\YPE�UL[[�������R�&Fiڑvpt�^��mϞ�i�^�k�G���y��hG/T,;Q�Q!]����mS �?�Vy��սlOgs��k�E[���=��N���E�q?τm`_%7��k��\�#��i�,q��J+�]�]��Y�*�V<ҹ�<��}�C�zp�a���h�ŷ��^�K��7����C�*��O3,_���z�Y�_c+d�z�L�������Z_�	�~�*�c�z�b|�<w�&��p�]���8�A�Q�&}�V�.�A�'p����N�#��hӓ=���
JVs/50��_���^�F����|���s%�a���Rnj��8 ��ܷr|�Ř 7^�nx;u �`c��F+�׌� L����� �B����$���:f�+-7?�Xmm������e��iײ�BI�O�pc��ݐ ��9]@̼��Ģ�KDj��ųؚ)�S���:]u0���¦���	XNBf�
�"�D-_��7Ó�#"9!q�:� ��G'Z��=�._�D-�+ґ${V�$P^���D�VY�� �K2����}xt��!ԇ9��ݻ}H�e���
؎��!a���r$��,�*8Zf�\¹��N�:*y
/֟��� R�S�Y	-�v��{�fg�9Xlk�뙾��[F�BaF�rI�#�rg��Q��r�	Kۨ�y��.q<�a�׵{�.' �n�d��J"�uqZJ���:�>"�'Zި�O��,�B��t�Q��9�G�P�:�OK{XW@�f�ZF&ൂ���U��Vݾ.^y�K�g�	�������۾&�%@lօ;��Nz��_�H��U�e��WJ�?���#(�S~�����K9}��5`�c���!���[^|�~Mdu��(}�}x�ɛ�ӎ�n�>1=�;�.�^CG�7�%5�<�z��hn.N�O�s��
�xb�x��^���兲�cgs���ڻ�}�=�a!N��ٔ�_�dMLg(_�Ķ&�(x?2L�/���man�m�-��9�J��Y�q���5F� �B��R��f�Ą�{G�et�[f2�^6l)%8�Y�e�,�i�x(�M��_<=)]����l�DT��R�e�
��3���2"85����vs~��Q�޽~����T~�d���,�ɥ�s+me�A{��{mq�Q�_jC��짠�I����0�� �Q&G�UT���L2�Fr�ρ:m��2��`U�R�l1hӷ�w�~�Ͽå�8}���۞�O)2x�~�Re�08�ʠ�����JHf7N�o��㣜ty?<@X�N�dϺgu��y5 Yy���_���{��>4�:��Y�z򯏭_��{]P�C��7�q{�vv_�\���ACi�h��:�oHq?&4>�1���w�R�v�w��ʲ?�/.Nr����>*�dǙe�ە���6�@%��I��K��yK+RW<�wy���Q��/�Z[P!ܥ��x�_ɻ�4�#ǧ�&�s�9}�P��9*���1��
�m�+�,L���O��y�޾~�^<ڞ?��橄��7
y蘃V.Ǉ��-x�7U�
�K�a����ʒ}�3�;�J�;0������,�p'+U�QgD|]RN"\E��QT�k.���<����b�s�!�CF�JhJpD���05�i/P������V���|���Z�<�Cm��)��A{�z���/n�Y��\x"�P,�I)$��0�0-=�����:�mΙHK��Q�R���=��7���vO�7���Dz*���B��\nS�q&�� ��Z�|ܽ����(��笙K��=O78����_x`��U��9� �����{����e�'/�6 ��aF�6�H�4U�	_P�A�S���QT�O5G}�-��H� ��O����^���+�<c�R;�OT��k��w�#gԒ{c���4]��"56�Y���2��7�߆���I�e�{(�0�w�?���ե%t���;??C�B�љB�
��<�����~�O�V�t����4zqAl��${d�/£�"d�W"fX�4�Dւ�>��OFX��$���� ����܁��`�I�����n��/�{�߯����>Xy��pz����Wl~�L9"���5��r�2ӘJb �T+]Kr�bMW"�@�+���(\�����OB�vQ������;�#��6�v s<j�(_*`{�._���<�a�Q��w�������E��m��:�s"R��g�������\�_�7ć��A4����	�g���,R�)e�*�BbW���q�W<;S�$h��+�ClL$݌l8z��dү�^[흶
���w>��M{��_Ol���>�d��3��z��
����c��i�$b:]b!bb�[���џ��+ߪ���>4�1L�v%xk��$�Ѓ�Y�F�j��X�2���;����{p?��Q���ˊ?������c�9☰�U�����Y3�'/�ב��r�y�m=��Q�h�D<�	�tI���<My��3Q�,�'j�w�����&�����ni�z�_nx��e{��ut��.a����'s�����?�N��V�f��e��n~J��zQ��t�rJ��S�*�5����;�ȫ������#D"\y��ji�3of�q�Qۼ���/odi�����t���.�^Q(��K��[C���%^e|�k�>��|�~h��7&�+�zT�nDyusV��.�͟�r��se�-/��ٙ���~Fd _<ms:��Y���$~'�;Ęn��]e	��q?}�W�QHZ{v�Eڧ��.7o=��2K�\f7�V)�|�ï:a����Ƿ1��C��S���*h��Y���y�d�����GB+L�Bj�m=˿_y�+����~���~ݤ�.u�@��^7��Q{��!�2���:��Q��y�iۖ���9��Aȵյ����ʖS��|g�=��NmVѓ�L&��o6�6��a�w���O���%��r�G��¨R�p���`]��m�`�Up'��A>�n��ɣU<��U7��$���B�k�/����/�
|B�|���5t�K�=IU\��|���[\ms�
ӣ��N�L�7Jv0=� �>]�*���'t�մo�-*rgA��Q����@z��S��
�N� 0�Ȼ�G��<�G�Q�qŁ�ce#�)+G��o��k����AP�.�Q�:q�*!�`���rr��<M��%̴T���C>*��x����Z��k�ٓ�[-������r�/P�u��y�[���-��7���6o��=0���k
'z�ŉ���>x���<�������*?�9�s}G�v��Kii`�`��ZZ����\a��k����<�/�տ��W��^�k/ߠ�;��%O�06z���I�B�Qe9�0�4�D����p�5��	7�0bC�F���o�;���2��&�@P��9׋f�?�+��I����J���\�92`�JQ�5Z�hXJ]�5D�S�\.x�����Y����N�S�X�S!4ZuWӬ�(��ٗ��g�c�����>�#F�S�Ѵ��gm!�^�p�R0���(u�fqOڱ��"S��CйH<��Ҕ51�A;���+��H��'��8]��K7�g�*K�TX�|s_@����Y!ʣ��F@�2]i�l2�c�)��b��s\6B�,�,��B�:�֓���e#=`KL<㦊�1}�7�7g�N��{��]v�~2�Z��2�LP��LV�rN�l����Q~�@m�u�m-���u�R���LS�sqX|�i耖2Kq�}���#��z��u���&�r�_�"nߗL��R)ui&������ix���;�E�O7A>4��w���bwO���&���0}z�P���R�d�Wf�,֔��
��B���t��QX"qGLk�'�AN%:�$=��#�&.����4~sًiz�����Ks�'�4����^{��M���%]��΄K �W��9
�;�±�������k���8?Ֆ���uEP�/3�T������*hK��޺�+�/�Ii�-_���!�����>�fq
��ӵK�O�I�Z��z���x���"�d���RWg���]��no3�2���9�G�:Jtfrie�m�\m���-�n�Q��^�l�k�͡�����H����vſc�� "�W�i~���"&ƯĊ�lG��v�����=5.#3��
gf2���������;�^	**�Bo�KFw̷��)aK��˪�:�ү�}��)��T�}���y���77~a�. �\2�R8+�g9���|����#{(b]���M�ǯ���P;9��{?��(����
� >�SKl�\�T�QQ^��/���GaD?��<74Fz���Gy,~�{E���qx��m�Q��{(:[��Q�<�}�;�_Aף�=�]�h�vT9[_['�V����Ͷ]Zvڔ�IO%�i蚆ߥ_ƹw�^�޾�=��}��'E�<� -�?[�'픎b������0�o�i�(
����b}Q��?�n��̏o�K�1�
�=�����S.�+�K����US�_*9/�/ ��`�{����a{��u{��eہVG��>⦴�-�,�;�fȑD#1���������C(+����[:?n�g����֕9�S)�h}���j���7O�U���S�����UW���_d�Vpo]�ϭZ��!�p���Q�錯qTv3�H=l?��6��,�s���0�O�קg^�L�Չ0�-8N[d@�Ft���;L��m�kf��+ۻl"
v�1�����V�
w7DL<��SiT��ٸ|��]Q0|�.�P�BB�|��F�'��)9�{N*�)#{5D.��O<������m����/2���F���Z�>{��^�l����� C4K�P.��)�JV	��=Ha;��RS���A�g2�3���h��vl�f$i����X9 �۽`����y:��ʽXވ����/&��X�\�xp�d��ߓ��up�WɺF�h
Ht�R��Ni]�� ���Ue��ړ� �G����"c>&���0�|I����HB�<+dEh7/:`�(Ȝ<*TEK%�N�h.��� �%ZI�KW���Hk��W�B�:��K^r���� ��eNuh��xB���{"<�W|sͷqLG���SB,�_�M��`�i�<5�Tkm���1Z?a%V�@�^巃�l�ˋ8�����㺔��D�(G|\&hy�_��2���̻4"����!�*Xl]�ggT���.�2�a)]������c��M��MQm�O3x�&�{$��0��}`*�Z�R�B�Sޒm���{|/k��wM��>Ĥ~�������=Z>�Hy�q����ζ1�*Қz�����w��K�>QJ��sQ�dVtp�t�X4��J��	f�d�|r!"
~^:&W����O�)����*��(Y{{�{fg�yȤ-?5�5�B���W�"q�tGpʲS��k����N��-δ����4� ߩO�I���Kc6´Hĺ���~.|�'�	l�Zª�kcĵ,·ڸ�0��Z�����)���G����-\Fj�����:Mn�Uf�NO�i#g1����l�}REam}�m?��m���-��k�3K�Be�־��Y�^�
�H��i��Bv~�����܅�o�\;�箼e�g��ђ���~Y"�2 :�;0t�3mye^x�-AK�f��i��}'?�`��n��o��fSe�ME{W���JsD�����z�޼~�N���o�	��{��G�������৸K���d�*��t٩�O��O���C��
J��AB�����O�F��	#ϡ��o[[��;ߥ��H�Yf!MR� =�-���C��n�k�����O?B���l�o�Qz�5�۾��B�^�Н�� �a�q�o�?�R��G�I���6w��9�k�~���Խ{�!�c*g�>�����'��������G�'��X��`���:��̓�ۈ�3�G�/OBQ� �8��M�t +�G'�}�eW��L�)YE�_���
��zLL�U.�+s��'!���˹'ka�\ADl;�P�P���l�v�FƬ�%�@��W�T*�N*6*��o�f���U���T��2H���G�����@��2=�G��L���:�S�\��l��HY���]�����%����]�P��,+2N�#]@6
<�~17?�����Oc�Bcs:�몌�ͭ���;�LO�O88pzz���'��ԓ�Ѷ��\
����c�����6-���Mx�3q�U<M�F<��{o�~]>�%�|K��V�q}���A� )������5�s� |�K�y!?hm�`�ॺAn�&����N}��m����Nɺ�K�NU�^�Q�d`$eǑ8Q� 6_H�(�3Y%4��#��:�;�i^G��PQ ��j�
D�?Lӌ1�7���KAgg3ra^.-���_J�DGb���AbKgZ
<v��Ʒ��v&%�v&��#���%�(�8��ӎ@k9uSO��!�ޤ�WB�i��y�ȉ\�9`�T�p
R�g ��ˤ����� ٭{~Q���_	�N!������{e�o"K��PuZ^�y�9y�UB�)����3���!��/G���0�4�2�N���A��������<QP�ʣ��#Ўg\<�HW���t���p̲�9LB�����D�T��q����#�S4�3g�b}/Ƣu�K|�t*g�\��:��1�3��awo�wV�d���Hǋ�+��JV���e�7�M?a�s���F��&�cӮi ^y.�!��5��4�b_����I���2&F����5a�s8�\���X�mcϫ�~��{ؖ�ֻ0��XO�]r� ����%sc0ZQ �~�T�7�Eɂ�m�P���a��d�7ΐg)y�K����ʇ�>�,G"K{d�G�rG֫W0�w�2�k��������*X����.K���1�E7�O���8�z�ٶ�0[�^ ���âdQ!�Z	��.�r�xc?���ܩ䠈�O�d��<���]fb��l�G�(����c���U+U��ߥ�abX�SG|�i��+���'=/���[&���woP�N�0^��n�|������mikj����4��=�6,�q���fr�
��0�1T�Jt��:�ߗ�N�[M������1}��rY�J潎��*�Pw�vw�禢������C�Zj㝂e~����>u�������l�O�*��|�x�7q̯�R��kϋ��Ľ�<�_;������������4�N�v[��-~���۶�F�i'��#���./T�6���v}!&�7KqS�p6X��>\�0I��`��V!:3^�3��eπ
m:�����H[\�C��h�|�%��)[��+뛙IX�\ok؍R�����c*2��(d�Z�M���1������ %�!��KU���}���V�G��b��Ҷ����#i���Y���v�@��9�0�N �:Kۄ���_�!���
7ɑ
V���d�]�N+��jFC��&����g���+�^���
�ɩ� ,�0�*X��:=3�>ޤ�mie>x����s�^���@T�.�9��rYNZ�t�0ȋ���u��BQ�O9�_*XC�**H
�|U<9�:�%�յBQ��c(6��"F��'b�d��;�bY�x�0E���Ҡ`#ܢd��@�y�o�]���&������p���\&��5����,��qԮΎ,L�*GE����Μ�'���
����vp����(�KT�Ϩ`Y1�Eᄼۗ��۵{�#X�o�y�I�ʻ������[lf���w�� ��?h�����_�]�3j�@x���
����"��J�;�W�qRמ��а� �!��'φX]qE�6J�F����3c����_�o����r��C4j��1����C�3��;(Y=8�J�̂e3.
B���]A�����anHB��@�%�(f�S3�B���N]v�Itn6s��ʖڹ�4 !@޿%Db*��NɢO��J���{�$.v���
��? (��T}���s	ߒ/�z���[�^������D������PH��%�#�,q���Ze��)�UQ�A|��5M^S,-j��
Pi�]x�D�=a|�7�Z�9��w��X�8*:��:*�8���q)���K9��t��e.��V�"0̫�FW��'
"q��raYd��VxF��Q�*Z��xx܎O��:E��jO�^%�����wf�<�½ c(���R���ɮ��`������۔��V-_��i檫σ����I������^���l�X�.����˴���{�I��W����[;x��e~e�ʿ�ݴՐWe��@��A?�K��/���L�������94pu�Q����)Pa�"���v��1⎩���0�ٙ3\��y(�)�����~ƣ��`���.������a�	��������i�\h�T��(��!)_��m�i�2M�
#���ё�631Җ槢d-���`�Tg� jO�L�����\��%���#8����7$u���wyeI0��E���J�7�D�N�C�);�h����ǂ��Pa:U6��9�[��x��!Ԝ����ɗ����{@������at���ǟ~�=��{miu��NΓ�D调~����RA[
�~��>�P#lw8E=��������2��'�w�Τ߉ ��.�D�oB־�W�z�@���^����vN��ia~����3��>����R>��k����M�+L�h՟�	� ��KE��=q��y��e[lr�;�<�ަ�~���E�*�h�y6X͢�d]���EW]�7gf����9�W͐�Pҷ�)��w��Ƣ@_�����	���rAK!�U$����^'㩡�^�?z����#y�{���fg� 
iM���,.,e)��B�]v	�{���<iR�w�1����"����Q�����h�4p���s�R|�A�p: ���d�Hz� zD�N{�"�_ZU�ͷ��5���`U�T�Ɋ!ܤ��Ƈ��<k�T�;�^�,��k�LP���U���禨̩\ -R���s�ˏQWQ����>>�ho޼�f�n��7�\877]_�.������<���3X��q����Qk�FPV�Z^�n�o���C�{봩�#i�E�͓��kЀ|�Qb�g����1�V�w&��{ѧ�W!r�}V���߫ +y���Zi�{�,�C��Qؿ���Ľw����b8��EX��~�+ҝp���<t£�=��af=�I��̖ף�=h�˻w�#4��6��=��~ܠ-hC�+���~�7�.&oXc�|7�A8���}R��@�0�4�A����+\�qŽ����盳X���V-�����Bu�y�tE�||qIa7��א��,-�F��d��=�����f�2�Rip
�+Yޑ5%b7P�
�2�{Y�D�"��R��q��T�\t%H��2�D����$��)b	�B@?zquMg@�ZX�o� ���f[[[Ɍ����^{tvl��r&�%�
�"����%�V�����z鉎0�HD���g��<]����g!�������:Bb�ʕ��ǷdG�j�A�:}�y�K�,l��W�88�Vǖ�U&35�i�M�v�J�}W���o^Ͼ-��(`��%6�(w�^�K�03ӗ�!�T�I���kZ�8	�����2\x����])Y�u��I�-�	�3[�},�'N�N�������`��RA�p$�%�W޽����4���������^�0L�m���_׶2��'�����3ɳ�!��ZW�֯����"��e�.	��t�e=����Y�A~�&�q{c�����ܥI���aSK7T�J���*) ��������W9LHEIa'�=�*әɂ�X ˩Pz�e� �����ʇ���
'^l���U�f%n*ԩ<�=}�M.
u�Oޒ��N&?ae�*�"�B�z*h8Z�R��鱶���87	��i���r�2#��4�_��`O�������tap����<�����2aa=s������F��Gy��)da��M�!�w�
�
 ��)��!��ŵ��Ҧ�J��/�}	�~�O�5mt�)���\�������wۣ����7i�iJ�@�R��i)���W�Xe�����30����~�OS��[��R���e��h��x��(v�`�l+��pf�Ã��Km�*��=�q6=av7�$������ٸ����3���>("h�L�
|x��y{��v���]_�L���]z�� ٗ�o9֥�Y	��r97�^K��U���c ��s�A��*L���~���.}�5JF(z��l��~a�6@WV�ؾ��E蕬�Y�U�Y�����ݔ��k)�'Ε_][�����=˴�Q
IC���5r����NA��HA�ԍrG� �U�ʻ�����w�C��yL8��Ŀ��Dq˄��/�Ox�	�� +Z�f_W�l5��Ds���K��r��N�MƀJ�4�4 ����ce�1`����>��پ5�RhuwE�����'�y"���2aTv�Ǐ�,m������,4�l�К��h�K3(OS(.����J�����O����q��w�O?�~��=r��6�bc���.�U��������{�y����e���+��5����2Q�����F��A	tu�4
�3M��Ӌ(gK|_��ѣ�?�~��O�~�G?n���w�ý,7uCE�=~�����⽼�Զ��2{��%��>����l�����~t��)߾{�vQ����۶�r]i�5��O�����S_i|������חp4�1�$�.M�|�{�IӇ7���'��Ɂ�y���Ꟶ)�9Q��F^22�tk*����~d�]��8�ׯ�ˊ%�����(����P�6���?�^���Bi��%�3Yo\.��,�Wg� HQ��+�X��d�X?��'0��dYx�`�4�V\ �4�]S�
�dM���7<�Wcn>#}5f�HOL��V�N!"O�w爘N���N�9+�P��e�͚d��|���X��zp��ux���պ].(�U�*D�`���HT�/���<tt�{���������	��tJ��v��mf21������@�n��ݯ����XmHgW$�5B^%K�UT�A�)�aL�aU�F@�\��!�t`�ĕhz�E�##(>x:f���o��B_1�����Na�%,�Y�jG.A�\��1�$k}�I`e��'(Ϲ\���yr�'/e�Ru��f ��,G��X����y�f�\��i�t�"B>�{%���w������f�^ԯ{L;�K=����?L૵m�ug�o���n9�3�"z�i����|�MA�w��Q`����燦�'�/G��������Q54�%��CF����;y��j���Փ��H�����J���2�d�B�e�߃��f��C�P���\ �������8b�h�gOړ'O��W/s����0<�O���V�x��:��_\w�Jf��MN����,�EB�C���d934�R�@B��;� ��3\��~#,�_�ղh�� v�]�ę��aҰ)ܫ�Θ6�
�ǰe�X�D�,ɇ����zAd��z����+�(��2���d�2@<�v�2U-�����?����'�i+��tf�W�-�[	Z��
�4NĞ�m)�<��C��]{���ml�o3��m	~Cy�$M��ԕ?d�6s����|,,G �rP`����Hb�7�����o6�~��*��?�-�\��<?�i�Ϟ~�^�|�������9��A���f�`���kh�}���K�lR����Vr����Z��|Jس3���Q�
�.��?��	��_�la�˙ES~��	By�]#푾.?"Q��B�ַr/(��]�P����iٕv��6B����P�#�e���� -6��f��S{���*�� �3��<@��R�Β)��yw�����^��Ʉ�
�TO�+.�ȒC�I�+Z����!�TfU��_�`B.���w�:�`:�����v�NE��8ٖ��=��O�a����(��Y�%�Q�F�ؚW�8�����{��ݯv���Ї����ڦg��##ȏȓ�(Û�k(4�Q���ݏb?��~u����E��\Xg1=D!��g����}����q�����p�'�
�}��x����3Q+k+(V+Q�<��JZ���;� =�^~�E����滲�'3{o�'�.,����0݊��{�<P��(�IM�e���b��,�E��]��xᩯ�N�J>�t�8�\�@��(X�Vg
S
��=؅�s�-q�*���~q�I��[o����nq���Jl�$�_)��{��r��{��#T�@RD֒�x��,g��h�X��v�����"k�.������6zs�F���d�3Yov��A-�$�,1�aA�.��/ۉ�0@h�,`��a�#h(�� B�p�C$�'g'��4�!04I	P�HqI/#�����<��\��0��u��B�r����v�d�Z�~
[�PJ�M-<Tk����J�nM9�M��QZ�lc�k�V�'�PW �		����o ���2� �c�D���fy�
c���/>���b�DX�:�3���Z^Gp�(�B��i�z��IL҈HL ��4�׭� #4-GK�A�Y΁�hD`H��U��~֣]�(���d�+�--�0��Xf��/3��P<QQ��^��¾��m^��RS����)��5tI���B,�(xC���i:�U�?e��W!IԵf/��J��L�\p������F�Z�Իi�n}������A��o	���������\�w�RY�f�%L�c��O���m��(}��6$љ��Y�`1��ͤA$��x��6t�-i��&�ry~L�:z�]@�Q�<��Y��Sg*���E��刲x���#nk����&8�`]lH�b~Μ/..E�r����2�{�6}>��y�|�^\>��a� �M�z:s��Z!�B��P�96VvL%�٬	��Ge��*ʈ�<��d>u��i�H��@8�Kr�-���x]�V���\J;��΂��f�\����~D�!Ţ9
���v�;���=䌂ʛK4����N�}���}�M8��}M>�mve�N�݇�DyߖVڃ�?o�>�N��z�F&h�R��p([ʣ��+Y�=���2�}�l������X-p�;mW��9�Z�
]�;1���ԅ�n;��e�.s��7�f�#��?[���;�6�[����l�3�O�X�v�+���ଷI�+*X{��+��'�|�vw^�����dA�����%���g�`	���:xWKt������d��C��u/�|���V�_�zdg���p�����?4���y���pES�!9܀���#�L ��<��N.���uJ��kF\�J�R���H�����5G�­	��ʬ<e���,J�/�����z����8|l�$߼���[d�W/r�������%�PMҵ�W��K��G~.�~��f���S}7߰���C�"���W�2�����˃�D�lk����e����WG*�u��{�֐�T�~�	Y@�R�R>r�a��1�3M8g��m���D����V�2���<%�٣�%�����1
ѣG�(4��S��?q��K��t΢�Ͷ����ų�8y���{�y��}����G@��B����y:�3Xmg�Ӱ=!ғ$P��3a`�:��q*��?VI{�&(xpBT��f��S�QI�.�$�u�E�_��<G��1���������u�Z�����W����w%�`O%��>W���,��R�ݐ|�[��y�� _����ޝ����5_x�@���0��/Qz7O�&�KSy�����c5��<�e��]��S�R�\�:pE2N�v8��+k\򼶲�D�By]�Eƾ��d���/w�\p��!f&���BQ�y!G�{��d_.�P�)�������.]ɚZG��}f��cT�Ѥ /�X�8�q��͞�/�s�h�N�������w�W�(1.�k����v;��u�=�rAg�r2a2�%���q��UV��!��n!E���K	p�7�3@=�H]�a|�[!��2�k[�d%|Ӥ�wg���e��6�l�Y&��hRʎ�"�.fKz�����[l~!���;��V&���B�$!�P��DȜg�H{ɞ*�շ�ئ.��~bT�Y1�~6���K�j[��H�3�#(��;9�m�c���d&��� ����:3v�LA�Q��iO�ry��ݓ�j+
VXz1g���ő��j�� C�Q�j�b�bBwM��`^�$N=��j���=��*#L�O��[����c@�ͣ�40����aꑼ�E�nX��Ԡ>�i�o���O��E��"�'n�Ѧ*=�����Jn��p����3(@�t^���N%���ER;.gu��
���� N�J!�A1*�*Ys��0�����<M���g��ӧ�5ω���i`��c�#�T����+�*%˓�܋239��1֦�xy??=��^Fy���-�SЫ#\�%� ����0���d�?4�7˗����6�^����+`S���0%�ɥ�0��=�W(��6�0W(��g��M��;������'��ӯ����=��S�:��S�����<x�m�Y[ۺO�["OͳN.�P�W�����D0��+@*����x`��C���~?���o7U>��WU5��G��|���N�������r*���#C�]�{���z�K���pwMo̐����&���N�B�&'G{�����o�_���]�愠���Rރ�J���d����6��`���D�,�
��Q��&�3&�pA�3x��X���"ցNQ� �W����3�=�6BKᬉ�Y��YTs�֦/�7������V���wg����U�Zn���sƕq��iV���[��׬��z�U���	�)C�Ѹ�g�h����>�z)?a�c�HZF�*��:x��իv��x	�}�M��2e�>���Ӵ�S�<Q�C�Ci�f��Jds�4��gy/i�R��_�<���}h~�,,4O��y]��S�tҋ���7�ǟ>n�����,ҡ�� �ř�Qh���B[_F1Z�Ef��1�"D����6�_Di�B�@r	��&vK�l���K�G�9���Z%zjj,{�T�VQ�6i���,M"�N'm�c͢��}�fjf&���Ч��\O>���Le,K
7����ʠW�,G�zx��_�(�8���ԑ|T=R|�˚�%�8�5ܵ������� g�����C�ߢ`��{%K� ���"�Sa��$�2q����?6��X_���7�q�����J��1�|o`+n}�_|W��v��>�;��M�6��.�d]:�V�q`~�앴(#w�7P�F�ۺ�ݷ����4%K�9�?{���d�x�^�ڍ�H�1%-��3:ͤ�%D|:� ��rA�{�����}��#�R��E����GK ��Y��!(dT�J�@�w㹄������IB���i`kb../�I��% �D���P  �H`TҤ��b�;����Al޷S�H��aݮAl=��1����<�SƮ�wt����3I0(��!��q!dWC�@��/#Y��Y�A���<��  ����ڬ�3�A�a��pW EY���l4�̀�F$���BU�Q~�',
F��v�X����b{C�a)ʨ j6.S�
G��%��]���x�H�A4O¼��@.ݏ23A��!$�P�so��"]{Ӷ��v��1��Z1�b$,O`Z���m�~x���yD#DB�Sa��0�||j�Yj��ޱ��&'y��ύ���K�"��p���������N��X}��F뗻�(]&G{�w*Nt-!��jZ�Ho�y�������/y�&J�i�ZU�����7��' �f�쿝��Ym�w����Kб~�uL��-��*�i1��f��N�F}��X�g��;Ȓ�8�I�h7�B���{~n!�M2xw8�}d
^�d�����["_q�&aE}�r����IO�`L����Q&^!��/���7�ٌm���081��'M*d�I]�H-s�_ӟ�my�zL�'�i�8=���a��e�����\9��/��d�8�B��-m��FǉJ5�H�w�}��=*Y����^��d��~�޼l��^����v,c�O��A�k�Q������n;=�){��"������}��gl�l�_��<�'2cm	��/,������eim�=��;���|��}ʁ�\��F���Cπ����4������V��Y���g����B��6+��٥�'�{a�QH�L?}�x��>t�M0ٞ�BR'�"`�tS�	�]�_K-o�H]qT^ �0�)O��
V?���W|6O5t_��p�W�޾@�/Ώ�/;�͋'�
֛W���J7x5t}��h7(���'�ÔG�G\"���L@�5>I{�K�V�p�]��Z�o�0哧�e`���Q�/���Q(�.m����O::JV39�	�C�5�l�*}��*[��v��X``��4KA�\AYayv�>K^�e肶�/:�&xl�CtA�;����k��!��E���8�@H�r�*a��6�6a=�f��v`��hC�< !*g�����k��s�#�S���612z�8���x-���5y��J��T���F_!�;����xr��Ma��5��=f(��JJ�q0ڡW�ʽ����1�`ۧ��ʣ��_�YW�q���{��?�n{�`���̵i�{�&�p�84���6���e���4�9��0�A��kc��s�/�������� �E���Y�.��[Q#聅D��/��?�*��XBʆ�n$�݋U�A֤�F��R茡\��2X�9kGǞxN�&�t	f_8�r��g.�r�g,83,];^�q�\���N{��E.����
��}��rI�xV]�AcE��z(WJ�l<랈Xy�4E� �&Mx�7,V� ����5r�{���R�{�xZ)]M2`-;ux�ހ7�!�"#dq���e�����(�zl�+��6Q�	Ҩ�-t�<>9�VV������6J��,�����d���.�������G�#��<
�K���733�;�J���K���HK�!�e�
�X�m�n` �� 6�R�)�a)~��j2��,%˽X��h�K9�2G��X�@�
�uǌMP�=YǗ(X^.zڝ.�L��(�c�-WU�l8�7�,3H�a�F$� E~����w�N�w���]\�I�V����S�lh�BZFD�J�{6|�����֤6qK	쐼K;��[ߪ+���-Aư�W�m]|5i[N����0X����X���8�S-D��%�m0 ;�K�$��Iqs�EsT/��R����:!	sԦ�9q�wpz��B(�Oe`�����i��l�	-�j_��c<�P�X��l~iFp"��u�_��O�wO�FXD�	�4� �J�+,6��Glq_����@T��?�f���%��?���?����� ӿ���Hz��'K_&E.���fo,��X@W�btk4�`U��i͂���ވ\�6�3���)�Q��!�Dɂs�� �����H�LZx*T�W�&<�ǿ�����y��K-��
��8�S�L��˗mw�]�{��moS��[ES����y�B��i�knz��O��	�]�A��i�4=�<���|j?�H�ߥFvY����;���7ue,@P�FN�����x��Q�R�B�U����������{��z�B�|�^�|
�}
��W(��\����U�:;=���Ƹ�ăD����DF����ټuvaNS���"~
��w\�+�QP̳*�xSѭ��=���IѰ�����6#2�Gؾ?ؾ%l��'տ*�JS?�9����,��T��{|��z�4ė�g��-�0Ho��)#�$�;vN���w���M{����~vD��* )����C\=bjz�M;p�!�9DII�zz�G��s�y� wt1u��Fp��@���*'�n)�ʾ��v��u#}��Z��80h�$�~� �����L�����I���2��j�>ଆ�#!A?h�
�K�=^��{�xv9�K�<�Y�9@d�n�s�
(3�>w�0q�� ��Z��J�qϱ��`�)��5����g��}���~��6?�D�'�7Ti��{��Q*���_�,�u�S>q�%���(���/{݈)h�ל;''�.U�%h�{2%�W��ߛ�m#��..h۹
&��ٜ�������ͥ�8��m-�7
hc��������P�EH(��������~����{Z E��+�]^�+�Y\�,a�\�?0Ӗ��+`�zz֎��%RA*��K��A9��>��XB�rK���e=���6�?m�˴)�(�93�}��}?́_�����;;��^0�`�8/LhKp
s��3�yN������2xHeͿVpPa�� ҄��mu+��_	,����v���� ��oE�1��䳦FH��><���ޱx5+��=��A/v���ٓ�e��0��(�x�UYw9���;��\[n��m�dm�����)!���������n{�L�k�Q��L����ܽPb>�d9�Iwiߣ`���L��g��J��=����]�ۆK�2��"�VV��S�\heu�md*��,� F�2U㘌��=Y��ߥdvJV�ZA���F��e4�/'�n	�zjcH\;g����P?��!�V�2c�b[oчƕ	���}�,$�����w�f�U���WI{���¸�%+�X�i�KFF�%*ߖ�p�D��y�W�KA7��ӑe��.v����<��+Jy�dM:��2�U��d�y�F��e'#)����$@�LV	���^NLz��#;���NUǲ�XM.���y�gP���-����I�Sfl��d@%;��i�o�i�w����m�|��s^㙮�[��Uam��� ?�Jk{%���J�K|���σp:w��w��o3BBL<�)�/���	bX�|ފ�NA��<'	܁R B�sh���bb��u��ޖ�`O��`���Y��W������b����a�.�p]�'/��B�.>�{��ޕ� �GS��K�D�(�)�ͪbԆ/# �����Q�fƢdMR|o�wv�Y:��q�ж�-?�5�>)���0��t0��?��������u�l�{�L��JP;� ,��RL/�<<D����1��޽��/���K��7([ox��!�pg��(W�J�e���kK�+ٌ�~��K�1�����=��F'�j&�'m�;ۂgg��b:џ�o돭~����X��_z����t��XS럥`!<l��Q�U��/��4
���{�C��Z�4y���J����2V
�{�y���T������ڳ�_�7(�'�$q�.�Z)X**�g��'��6;��+^�/!�8�/�@X����h��s�c9»H'�4ԡ�C#ӡ�����9­�Y�7.̩�D]'�Q}�j�)`P0���;�ib���4C�2��4m��e�^�wI�w1E9��^�������s�r�+��y��S���l�n�6�@�V<�ޖ�:P��U&��
��t{�]��{����h�gQ�vw�S��E�Xm3�DT�\�vA~(W9�:3P*F*45��!�6�I�(�S(ɓ�^��9r�
���t�~.s��Uu�ǵ'K�f^��"#R�Ș�(��S�m}e�=z��6�������p*�B}vz�b�+{ः�^��q�Ί�� ��G{�)�Q����I����^z�EP9x�le
g�<����<O�^���܅F�W�޶7ov��0
���~��']4�1��:;u��b?����*Vo߼n/�?k/h�ׯ_g 9�f@��Ba��Y���G����}�A2Os}���gO��J�_4����'���{���C珑�
ߤ��tq���>BᤢV}����O?�Ӿ �_b`�M��V!+T�eL�+l��/y�3��)�w��1�}[�]+���}��#��5�n4�Y��R��硪s	.N�d�Fɺ����C��	������W������+A�����(8 ��z%K�O �W�P�.�c��N!��5��V��Fu ��8/I��Ց�bB�i��������r��F?��9��H��G1���%r5��h���{%-%��Ζr�y�t+�� y )���L�|(8�h5�e�*o����h=Ƹ&\�l���JW�� �D�[	&��%l☪�Q@�Qi����VX��ȳ_�E�R$$��	�@�K���Lx�c\��*ֺ2��K/�����L�±�����I���� OOx�k�Ap������j�B��x�+���¦� H�a(oa"B!s9���{�:��J����F$�!*� �@��pl��}�h���ʍ�c��6������u��?a���%�k!̵o�<�&3����Q�ܖ���<�����lͯ������pĜ��s^��}	�����]�K0$�I�n�%�8[�xp#q���*Y�bɠ���`�d�}�}�U�R8UX�>
��p�c���V��+kmk��7s��eR��.��o`Z0��#��	@i�x��C����\�_*XCm"3Ycm%kJ�:�����R�����W��V{�m������;��t��FG��JK8��ܥ�eMIÑQa�r��$N�| 4��x��;�;��.B�~���a��N���4Ʃ���KK�#Xˁ���M��7/�]_�n�K�h�r�ĤGN˻XcA;�����I���
*�#X�f����/��M���n7#~�>>���XWG+l]�j����V��OS��oY�I�a�+�� ��pL�(t���g���*�ǽ�G������_��O~�<�B\��Y`"/Oޫd���P����i��,�h���qg�����Y�ߚ�N˾��G�G���qV��k޳�ŢQ��N���Y��^ H������d���^����E�8�r(�ySO ��kƮ�,�'����'�ȲW`l�@Eڨ-W�\��oA��S'�^��}~J:b� �{�s�3)��Px�<��N��ha�౳�A��Q������ꎮ�Sy��w���0z��7�/���|��z��4)�CK���;������K�]��^h�wW�w�%�+9la%m8Ш�YGW�(#~�=�����(QBͲ�*Y*�����m��,i�']/��e���,t�9SHX������������(��+���}��>��(��('�Lz�m7A`+���I�J�	��3DQ�T�����ur|����n_}�}��7훯pxK�*8��[��#��kevv(
�����q�.~�_�i�P|���)
��x����n_}�5��������4n�B>:q�J�+���k�E�O��ϩ��(i�����`dx<¾��/e/q���\���ի���<���x�W�v���IlSZ/����0:��j���j���t�>�{/eL�����5}C�g)�*
�����T?��Ի|%��$�D���u֒Pf����`"=1j�0fmz���Uܞ�G�_i�7۽͵ܑ֮NT�������ʙ�~�����3jA�"�%���\P%�����,K\�Əp@!���|��6
���R�M>�L�P�26���{��|2�Qh��/�dmR���e:�L�x؝�nT�Lֲ�x�<�}g�s�Q�U�(~�Z'L��Y.�ZQ����H^Z�g3T�����3l��d�H����׿��<d��!l� �ߓ�
�I`c��:�C{�2e4���F��s�#����"�H�n$k'*$��&�����&O	b���J���^�O?�K�(~��e]�%����i�I�k�M�m���M��m.\n���(���H���W�ê�pF�x� Az��N!���F�R��\��Xh��s���5t:�{�T�=�F<��0��|��`�y����f`�~�.J�t�+A Im������"}�6L!����a|���á�2���x�F��ǿ�J�{���W&n}�w\q�7��{uF���g�,WB�0����P�/�к�C%����\o4	��j�`E{�����U@���Y��;�e1���v����F��5�wp93�����.E�2�ů�V=nDv��ik�#(�T�3Y�ӣmaf<k���I���y�~Q�R(��8�*��:Y\F�I��[O�A��Q(��[��0i�0�׺ڧU�\�9L�,%�d8�*��Gםs9�)I�f^,���S㔝6�� Q��ff=-k�-�hy��\�s[C��D [A�D�������c#����R�pP��[o���&�y�ʣt��j?Ʋ�.&�:8ܕ���E�9K���T�gΏ�>�oЕf�_+=Ɍ�
S��*�< �~w0Ke(���oT���K��㶿�H���?��2��D�R_��V���>��;(�ĘJ�Wg�e�{��8�d�"�<�Q�����P�lI�c}�\�6:1�;��c��༳ԎN�����.�rf�W�cE�J�Q贏�
�P`n����(�WW�խG�K]T��?�n������B��A�Ύ��L��F'��g}��PP��2}����s&���!<�3��Pd)��aM�.�;1���I3�<y:	�B���HN���x�������5�"�S`���s`v�TA�^C*E(X.�B����V3�(;�[���ǹ{i�:�$ʧ]�vN��/Xg�(߆�_�^�J�(�
p�����g�8.l�����\:�!lK�mc}����!����$
�a��˧���e���:���=�z���}�����<I����� mC��PH�Q��vp�P������}P.�����^���E��/�l���~��/��_?��J�^޷���^;DY��n�@����=�U�}���ѓ��/�j_|�e��7o(�K��g�	ʗ��1
Y�3r���t��]f�^��y�b�������K��[Ξ�e;�cKq6f<q�MX�~�E�M;;9ρ?�!�p00<���:ϴVZ��hWM�>�k���o{�+f������D���q�V�u��_e�����6(�/�Y���ț�c�+�"(�����uZ*-��~i��ijb<w����h�Q��Kɂ�����_��3XO_�=Yu����Y��dn\j��y9��+YE� ���UɊ�E8��a�l��iXv,���HD��h��*cu�'�؁�9�� /^__ɽ�k(Y�i��B�!C�T��ɲx���A0��l�*Yg����24��E�Vp��D�L����:�!V&��9M���'C���IP�[��]:�p��U����H)5�$h5�Q�g�W��L&]��t� !e42�H|��'��+�҉�&?9�$e��'P�����~�~�d	���C, N�����I�M�_a31:�f��@Z��:��f��h��FY��wy����d�+�w
"��Bw!|^���H�ȅǱ�Lp	�j	b?�/ˁ�6i�dW�‶����B w���=��X�Qo5��A\�m��ꄴ/u}�x~���
�6��3qK��1�yN�	��Vz���:?�R����=�7��������㧠ЇI���]B�`��]%~nx�������BhxT{JɊ��Tu&��Y�(/�騰��_O-\��ޕ�,T ��*V客%��2�o��#�}E��2G�FP�L�E�g�~�i���d�UT����p�<���i	�B�JmM|���u�=���YD��+_�i�ٵ���L��p��S�k
��=���8F�G.$�Y�ѣ���7���j�F�rfؚ��cqy�������dI鷩pU��W�X>�ŝ�E��0��p+��}�������&}޶�98
�#@�F,ķ�I���/�G\K��Ǔ�t���^���%`x���4���஗����G���ܙ̽����z���/�^>��7���Eh��8������ʞ>J���y�QR��ֻ�\��B\�M�(f�g���s}�0]�o��Ik>�w���i;9s&��9He�sU�~��Xo�ܥ}��8� ���	R�+��y��bv�OΔ�v�����,�=X����>�{�r	?|�*g�J�)YGw�ƽ�ac���٦AE�� n�G�2�(XIg*��� &@ٿ���d*�����3Y�p�x�����e��Ņ[&��ߙ��@�p�i\Gj���(�]ў�/�z���~�=x����f���u �_"wA����/�	�"����"Z�>�Ҩҁ�v���T���{\���Q�� �����5��n����E����Qx~ٞ���ؼF�����M{��5��׳���)��k�%��7�y��y��o�W_~Ӿ��I����훧/H�E{Fz/_Vz/뷿������˟����s�+`�l���n��E�:@�}�Ӟ�4�$�w�vPjH��/�n��嗙�zA�v	�O�����!޻��w|��a�F�x�"J�W_|վ������-��y���e;(a�ڝ]���P��<��RWk̢h9�vA{�z�����Q�N�2��<-��6�hI���VF�?j«t��ٷ]~�4nϟ�m�G|y{���>O���N�e|�{��X�	E/�wЯ�g�~|�!���p󀼙%��>��;P�>����t4�8�L�V��`y:��=#7�W��?�d9���/ߢd!��d�Lx��;b�L�S����NX�������y����SIʚ]���h0BB�J�#��ųF�¸�jjf:�;���	��,����z�����P�� {%K C�T�FǊIџA��[%k��Nuڎݤ����5�Wx�����,�"w\(k+�%to�h�j�J�}?}�J�g��+bd�� I�Ũ�4	c�"`��s��d�%�Ѩ��>[_K��vɃi�h�Q�6V'�� ����2���Hp �aiSG����KG��a\�ܓ&�!-TLcr����"6�̔6J����E*�H���T	��N��.ڻ���V�@<�\�5M��P�a�󄟥a��?��1��Uf�p��- &BV��7xw�4�r������#���;�
V<Ò+iu�B�q,�Oio�M��'9��N��������)9Tz��w�L�oɣ{O�}�:땷z�p(=���_�7!�SW��g�'qm�=���xa:fn��<T�k�%�!��Ib~�	'5�U#�9Ō�Cs��ZF��]Y�>����@�e3���~,�e�d]ed�bP���!��� �t0�5t-�A`�b�47����%���5��������^P0V*<��opBJ�)�P��$KC�S�'e���Z���Y�;ဍ�0e�i�oG��Q=�$t$�̘g)@�c��%��+[��E�d)X�_ns+9d&!����.�/M%E�B��M���?�W�6H�K�����7��M��;��� O��
V����q�J��lqB��O�,K��I����.];�>*�K�U��o�Y�k��{��ɋ���(P���Ϋ�������/�\}��_#�~�v߽lg'���	x�����D�̌+xf)4�8�+�rKӳD��+@��t.p T��G"YZ��aj&��.nfF`E��P|����Ke �=G�{��U;7�$)�E�A>��)\��8{ws�373���z�'�3r�/��o7q;9��d��Oʳ<���`�#Ɂ���%肃�*0��K��ߑ1q���c.�dͥ�*����,/�7��M8��������[I�!*Y��߾~�<��=G���^��O��A����r����=m����(�����G�ǖ�s�.�����C�(z=D)Y�i��0��v�Y�����<KǤw�~e��=�����>y��_k�s��y/����/�b��2�~'�R�;;��i.�S��y�}H;;{mo����ӗ(;ߴ/Pz���7훯��oPJ�y�,��K��i_�A�z՞�|}�R�����Ȕ-G�#�"+����9�����x�7�g�*9��Lԛ7oQ�������Ǧ+�+��`6����8:<F��m��I�q���0�2p��(&�}�CO�MTn��8s�����(Y(������(�o^y�ӛvB����v8� e@����4�$&8�D_����w���Q�����t�0�w����_G���(@���ʲ��/���8�}�߄Z&~͂���8tp��e�I��r�� s�ə|�u��c��6��6vq~�������J���G059�MS��2N+���!A3p����� "`(�Ȃ�
��U���y�A�S��Lq]�`#i$6"��:��"��<�]�����6�=��ե����Uv(ˍ�r�2��!����d�흃�*Y�'K��g����)�m�G'�q&�=������k�W����N~4����O�<Q�^�2��T=�>��PywÊ4a��_˻#\O��5��q���J/��n{w_?��̀�M%�Q�N�'/�S�F�(ɬo���H{�ɪd�z:�
����$8��f�<GQ�&FU�&r�P�@�ȑ��E�$=h	G���:���0W#��m����d���LG7=�}�٫�aɱ��#�uC��+ <�?A��hm���v�{�G=+ؖ����Ŋ"N���%T�H0[�L�?����/i�jɰKO�x�G�:ǫ�u�0�"�o����Q��e�Y�r��>����񑷾������)�(��M�T��2�̻�[2	�H�:���+q8�dX�S�+���S���*Yκ�h�cX� ;����MY�}�4`�g'9���ힴwp�ŝfO�Eܷ�(���0{�,�yf�����ei%kZ�,� �T١���hKgUd
>�L�j��PIg�[Yaj�Fya�/JX�M!R2R�̓O<3��5��uy���v�ݴDk�(�T|���wi���B[Zބ����Q𛚋�55���r�L�΁g�7f@A����go�χ��cL���/~o��GF��^�{��s�P&mK�;�n�Kp���Նso�~�B�+����p�]x��^;@�:�y�w߶ݷ���WO���b���7(Y_��/��,֛�O���N�0��%��w�A�U��}.�MZ�]�ec���,�q)`'p��BPhCx��]�����*T��3d�#���3��si�o^)3��
���u�N&���;:173�Kl?z|�=|x/�ЎO��
���2�����d:��vI%��<nb������{�b�mm�ϒ?k�"��{��I�+��|��Yf���4����i>{��y�|��|��H��3�NbU�<>,%�M�,W�\E��4F����l�_�xǪd98b���N��
%ke�=�?˥V�#���1�5
�{7�v��'��*<J�.��	q���o&�B��N���.m$z�&R�(Y�}�}rx���Y@�K��e��S��nD	w���|/��<�gg�\���N{��x�*���ۃ��C�}��ew����{�^{�A.+<:.e>WH/�keVz�lq�^:�c��#��q����&
V�c��1+���o��uP�v�� ��z����c^-�ɷ�k�qݳ̣���ӏ=h�܏����������7_���]���(XY6/s0N�,�M��]�ݽ�P�����G��-;[�,P���d�.>o���m~-S��)�vI�/%?Y8�9��O�LVR��V���m�Q�x�b�Q��0r��%'����K�����-hXFqK%kya�M��o�/��L����R�����)@�.��
�J��0n>�9�YT�T��)����5�W����p�(���.���U~�+ŋ#�ٷ%�]��(��U�-�|N��L��a���4��������O��﮿�v��|'������O*�G��Q�X�#����T�FF=I���vV贫mr;�1]�&�66��3I�	���.	u�IB���ע�zX�K�� T��q�.��CS�8=j�'��Ü�tqr�f���,�Ť0��K��%��bx�^<��6���57��.�rHZ�l��;;`�������àIo����"t�,��9�T;R
V�+��lbH�������%��[m'm��������ۛ�s*��f������K�2��$X��z�c����NA�l܊��l_��N��O��P��?��x��\o�d߅�c�����
�=���G #�݉>Ȼ^ʯ��b�Oi�4F�(y(�]����r��
AJ���T�h��7�ԓ�5_
��'iFX�7:�ER&�2;����h��P]��H�LF�-�e����b>ab�}�Ͳk���)XM��{\�����W�̽�EPHG�)��I�F
������ɪ���T�C�i�C6�RAA!�Fb's�Y.����"�S�F��~�J��4�i���3�V�l����F�[��~�@���?�!m��k�/�+9H�"�uO���^��yٞ?��}���3#��?��������/��������������=���[����W�������ӿmo�>������:6
������,L��[|K�:��L	���h�AA�{�N��`��I�
���{p<E����ٹ��F�k��Ġ���wf����^���M(g�/y$}�|�+;�$-��@?~����?h���O�?���Y��?�����~�6Q,��"��Ea���M8���3N��T�G���_/��ŭ���I������?�Fg��/����W_����"�S���!��U�䛺d��:��rd�r�L��W�� ��+.#�JW��(pૢ�+=0�%�s�ee������L:%XZ	�{��i⏂�
�S����.��Odt�v퀶{�Qt�E��J_v�Kf�?�<�{C�B��)a��'�y���h�*Q�֦��Йi��M����e�V�؃U����c��z��5��k��w(*���x�Lq��G*����{(\�<�}U^�NYk��h�p�V�ZD���mCF	RyRq>�q��<�7<��JY�8�@�>���Q�rB!�y(t��;�VƑ�v�*Yh��kmmm-8�~fWh<��+d���`o��.'����%9����$?sʊ������R�z�i���}�m3@�s�+��6��E?�d�tq��?��W��db-�������I�:�,� ǡcWgm�⤍ ӎ�!玡p���cīi#i]G�,i�*ʀO��k���]0<X��9�t���
�}���ď���ȧȣ�i��1b�T���.����D'��t#�7���+XvL�1�.�T/�=noSB�,f>���j�V�W�9FV 5~a|��߭�g�<�Q�Vr����txN�>%J�;��qa:����P00��d�}���q�ã3�9���=�X6@, k��,�r:gK�J��;��4�
��mm�w���T������~�e�(Rg�����^:�)� ��������zm/���qC�J���������^��?�	G痈�K�R�� W��Ns�=0������(�W(gg�P�`p�tnh
�;��ng��O�=p�� ��<ǫ�40}�%Lg��ޖ!d߿���w͠�C�	+`�h�_W�D�S�;��������WfP���{ʂ��-�>X���fV�OU#��a��C�~YĹ"��
Ƞ�]D�k�摸��D�p22i��J������˚���ΐ����}Y
8
몱< ��"4~
��	����q����x ��ϻ���2��'�� (YV�|6��MK�0_���Q+�����F�����������LV�5�U��
��Z.谌޺	3�RA��Zi9V��m3I9U��[��%��{4�h;BO]�@ұ>i�V�-��4����t�LB�����,Rk����5���A�w㧯I�l�r]yp
m��s�������V�m���~�l?��?o�����o�������/P���=��o��'_6�F;�{�?��G��c��ٓl��ρұ���s�Qx�B�|�YLy�Qi�~
��y��� .����uO�m��,��ҷn�r��۔E��Qz��jpF㌘�F�.m��a�
/㯭���>�����?i�����O�񟶟��O��}ֶ�6�_�S�R>���/u�WW?]/���/�V障�C�Y��/Q���B�_��g����h��~�?oO�=�^P�+;㱻�v;<���S0P\������pGڣD�u]�� i�W˯Q��mY��o��F��~�� ��a��p����4{�+�oϋ�݃'�wO��\�}Z^z�^���7�]x�iL�;���v�(�B���ʒQ���e��:��4�:�
˝�>=�����A箍I��QX@��gҬ�㥑��D�sвQ�aN��D�X%%����#���mkƏ��ܾņz(=�LI��������>����2y�t�S��ѓ6�����W��*�D������tF���ţ�'P(��4�.Q������ÆF2��i�(����H�����#�����������W��10�����+��۾(ZE��}4�qg�tІ=�����:��a�w�֝8�0�I����}���*~�y+�,�ֳ�ʯҒ���h��aVa�������6}�:mC��!g�Q4G�/�̖*���R�,�m����Ң�o��?{��ߞ�|�^��;k��������!H"H4=��8	` ���D�9lÊ�;
�)�xZ�G�*�d���ҧ3�D8O�q�AD�v(��A~1?7�6����Ѷ�����|��� @'���R&Ҵ������t��~��h{����^�k�O#]�Ը`�0U��#4�6ǐ[W-a�6i2��]���Z�W�͐� )�9p�D0��,7�Fд3`klH� #sB)����T�X>�eG%ގ�ĚY��q|���� *A�Ӎ:�]k�% v�!�	� C0R�(%U5G��0}sμG��bG�|R�⎽zO�]�Χ|;�����Gą ��7oX'���8��2@0F'Q'�)�X� /6?��,�i�c��j��]�����B�]�w��m�Y2�G���e�4�)/p�_%���+:PN��=6��-���v�2p/��:�6��36���!%y�`�ix�!�[�C@^��ܑ��tDIk?�����Ć4L���ԫ�����}'R�,-Ԓ�u"x_L�H!��1�K�D��D���G"a;�}�ߋk��>�����X���Y�c�.�.������F�f��#�c�kl�=Y��ֱƎ�jd�:�"Ky.�_t��'0㌌Cj������_E������#ܽ��=����,?{�t�B�1�RH��VuB����PV�q 5��1\G�{����T[�������v��r�D)R%=�#�p���L�z�>Agr��������z��0x.=󰗣��r([�\Bܥ�2n�6�x)]uͽCxH�3�E�TQS��(iO0s��r��?���u�ba~���fg�k	����r�]��MS�
�_�`�OD(�>�sz#^���� �6�^��������&���p��Kg�_u��>�M��M��>��lL{��'e�/�i;>|�@�e��r�!��j��Sů��#�p!گ_��"Ot��
�ff�R\Jӵ]hV�(���_gK�Ք��Z����
�E?����M�c��^�8y���G�3:�)|%��s���/���wH�����O%e!�+?(|��Ӄ'�D��n������1J��x����}����w3C3����,!�����ޟC��}I멢��8;v����%
����?F�����=/��kGأ�f�z����{�R>�!S����J���a�D�r?Ե���I�N�޵�Ͽ&���8�U�,�����F���*}v�vF�>>�錞0���VeJ�q�qy��p�=xp�--{"�r��Q������/�|��A/o�s��t-
�B�#�Q>�˔C9�?0'���3�F��1;r��Q�����r��\jK����ty�d$@�x���z�zx�%s���'x%�8Uh�K�Pn%�g�,��{�X��wPfP�܂�����3b
�p2x��8��r*���*�.��P��*����8X9I"A���s����6kE�6�  �y�U�0��v�����gdO3<��d=r|{k��./�C��/޾��_g��%�'G���3+@��B�*u��{4&y�ߔ�(���uU�cu�F�
C�K&�'~���?r�.�v��+�
��� ��]�}lZ��D� 
�6r��W���O߿V�G��bW�9�Q��]'�a�4����x�,ε{�#6W���b��h�2��Jֻ���z����`o�HT��Z�(M6��?�[���)_��[a^zeK�	W ���N'TI�U,�JD.�J�h|���Ph�e:�!b5Ⲷ��0��6q�f"��ᴖ	R�C�L:��� ��=��U,�p�9�ĪPڦ�<.���(1�ՙx��-<��}|ԕ�$%#a���|0~�R��$���>����>t-k�`i�._1�S�yэ�l�8T�>�g	Eg��~�d^̇64A�~`���gQ�-+L�9�Ar��Ԟ,���oa� \�ꦸ�;hk��S��z��| ��?t��U����e�G��?@���'$yܪG�:�������fy �P1�35�����p��S�`A~���&y�_}/\	���G���$��gT���	<�G?J�r�5)�Xij�|O6=�a̪\�5ܭIY�����#��}�1��zw� ��{TX�?�Տ���A��~;
pY����L��ޝ���S�ro��0�
���G�;J%]�Byn��Kk��i�E[,�����C�AhXZZl�[mee5����P�|����}�-�;�����T��#��(��Бt��U�p_����jEd��*|l������ ,�ON�ПiGdQ��W(��$o��Ս��P4���&Qh<��A�v�U��Ȩ.0O���]{�4�� GtNp\ԅ0�R�9��,2}zL�5-�&. p/P�������N�x��lLjy`����p���[�0�������o���������|�=���Ë���C�~����wP��hX�Ӿ�X�8^�����P�����?�h���p)"	��m�
����G`�s4�>�l'�ӇhmlO?,k��A�����H5ًO���v��~ �r`�=B?�~�u��z8|�䘚����u���s�8}��f{�h�ml/�o����"�{��kޏ3�����)�Q࠲s��Kɑ�'�IC�f=.����l����b����I��J�L�e�G�G�/��g��{��{*b�u|t����Q����m�����s�o��������87gI�Q��3�e�c�ey�%�`_�K�v@-�BIvoڃ�[�G�/�%2�(Y�^<o_|�u{���EY�m����]q�5mm(���hN�����I�'`���^�)�������:eX%g�]�܀�E{��y��c�_�@n8	��RJ��O<W8�-��Lf�����ٳ,�vF�%���h�wݿȋ(|	��!u�"m蚶�͙@|��߉+�Ê�=��ř�~%��Vt�\��zՌ�ư)�/q���|��6K=� ���Q���o^�h^ ��\��)����t��%��d��x���n���wJ�+t^���:t���?�?I���b��Z��96Q�8X]�TJ�T����]�s@����";Pn�Q(릙��C�q�nΞ���������:9�bQx���������~����c��O�ʻ g��{�$	�G��, �@�s铈"Q����i�d4�S�Q�x6#���S%+��{Y��;AI�\$�:���l��򎬵Ŷ0����oe�"�,% m@�����d��up辠�t�T��A]��e �4%����!�UC�(Y��w�@�J������������ ��<�1�?"h��2�2�VL\¥-�e���o��Ю�D�qYO�Q�ud�� �H����#XG�*���9�܈�(]�Y¢�Dx�_[3H�z"�p�wx�B��wY�V�*
֡
���+����'+ʳm�if�d]�:b��j\�s6�2�kz���?� ��U[�ޙq����=���c�����$�[K�o,B�<�D��3�����'y.k^1&��T��6�R��t���^��C=u��$���_��a�G���'?�U�.dOC���A��:���x�U2&j���>�M��x|���+䉳���d>���?Җ����%���~�2UK$��!�]"dLovf�-.������2[� �7�{\�w��v�r'� ��z��v���A^������6?7A�c�g�k$��0�.�-���w�侜5���v۾w�ݿ��ݻ��=|�	���ֽ���ݖU������J��_���u9I��@�rӿR\iRhe3��Fc��Ŕ�F	^Ja�%�~�1N�ʙ�����^���P��&�D��b�/�^���I�CSa����|���?�_k�E�� ��K�m�m{��
��vt�K�8py�m�O�K��hhg9'���ҭ �e�Pl���5�VEƙ 	�
�r����CY;�Y�K�7C�RVs���O{���.3C��Z5��W�,)��ܢ��*Y�'�ӽDipf��6W�A+(/¨i���.���-L�gfsz���J[]�O=Dn���ѝ�^wp����Q�¡̤ ����	_��9Ь�L���5��ϳL��q�^{�R����k�S�D*`�(P���~g��{y����T�q�v����U����|��6}p|b�-,����{�;��/�
��J�J��]R�L�Օ��b}��>tm>��T�%뫯�Β�s�D�v�q]E"ŗ�k�Miq�\ז�KD�O����d����\{���ѣ����J[Z��|zy1�⺗���)��	M��q���p�й~v�2���A"���G�r��S�v�S>si|q'�ŀ�Y��4����50���G�e���/^�͂�X}L�_6)��W���s)@ʹ�:�˳2�M��S?]���p�4Y���x�M{������s�q7[;�UH�`���� �2H���gJ�	m
C|��2�%<J�!n�w�/Sy<�3L��3=l�I�տ�3N��\m'���}FI3�g~��'<����r�mn[�CC�,��:!䄁����|��������Q��0;%˙��9]p��f��>��
 Y����3:lxZ�9rz,b�ĥ��"l�(5��@�".{Ґ�ϻ��	Ai1�� V���:J���
�mnv*3Y��žb:*[��k�$Cg�i��ɺ��,o�w�V��B��EҘ�*���v ,� �yDKJc�0�-"�TJ<$ZRK� l����s�5y�4{3��+�fL�_�&�:!�Ncq�R�	r�\AX$�Y� ��PF(��R�\
pQ~^�rF�,�Oe�r�R����QY�(&��/��X�I�3�O��3��ӳk�νWg(R0̓+��R�Q�h�c���3G(=�e�j4�	��#�{t/i]�h���;�%Q�ٖ�ԣ`%\��r�`���]U4�<u�~@�4�紋8����,J@��Ã�K�@������}*�y����g�>�v�j�v��q%\�wg����{�c*+l�c�~���!L����g�I�g�z2X}Uft�����2��	o�wy�#p��+@9ڔӷN���I�#��Bk���Rz��2���)c�n9��W!k�M�x̲3Y�n����PN ]vb���KuI���Ͳ?j���s����L����(:U]�T8	���i��u�6�\mn�o�(V�P���=l[��\��Q�K�ŕu�F[���I�cVX�~su1��'���p(����0�d�F�
*��� ���,�ZXt)�bf�T�z%k�r8�UW�t}JZ�s���mc�����|���?�_kP�k�R	rP�,z��Y���|}A?�����r�r*�j���٫�pO�´K�T�@؁K��ӫ�^Kϵ����4�����Q�F~"='y�z�萅��(�x��%� ��X�ڧE���7�pk9���(Y�$쀛�e]^9�k�@������QP��T7r�K�6�����0�������^{��%��[�K�j)�{�3�'���չ˶�d{Y�}�(Y�H`i�Ch�I��m/�N	t�^><)���٭���n�J
��xt��	�Ωd��p��B���rWf���*N��Km�����w�O?^ ��Q���q�Sx<aB��.�o�v������,�\D�Q���N���+�6��<qOz=y���s���t��ј�؆qh�H��LY�#���ڧ?h=�h���E�
-=���>y�~���l���i"S�f�h�l"|:��>I��I��0�z�3}���r��Nz�*�Q����X���I�ف�^ȷ]�
^�7k���fѼ�?�M�X�k�S�
����p˩ݔ+{�cӊ�Uʝ<I����x�F�}��]ZHoߵ�ƗgG_ 6�E���R��!�n�ۂV�zk����j�[c;�K�$��_iu�y��X��ESi&ݮN��`ߗ/yw6�iCy�4��T�7JA$��`�<�,�ʕ��Q�Q��G�9鳺�����/T��jOV7���BI|n���d�W#��tk��o�Q1$ ��i�4
qtk��G�|<"R�O��Ī���D������� ����Ņ�6;�"@��N���¨d�?��LV�d9�� b-T�$b���?��cT���.���6��,GWq���_�����`�K����j���ĭ��HBo�eL����7�|7	[g�D�~r�(���q����c0]5��At���2�!�S%,K�HC¬���l���12��.krM~��ʾ0�������*g�h7�c)X��:�=8�i^$�Г�!�wR�D�T]_���'�yf�$�./�dG� ��.�����Y���`�c���Tm�Q*O�I��oL��	S��$ʿ���P�^�LV�$V���~�#`�(m�wm
]����|��{�u;#������!ytf�o�7?�"Q��k�nT�g���!��ݗz��z�0BŸ{8]�1K�	/�J�#Ď�[Vg�=��E�}����^���#���D!̐x��Ɉ�.Oa,��Σ4�)؋�v�loo7�ΏU�H/3�(s�Jk��0�3Y�.�"{J��h[���R��i�?"MQC�D�3��U���Խv���(X��[mYe
�i&Ǡ/��)=�1����L�.���e���(^+�KK�N�����uי����)Zo:mV/�l�L?2��l�f6�05�ቈY*���Q�S��d�R>O.u�$�)�}��>U8���]Sa����|���?�_k��Є/����o���˃��=G�C�= a2�X^<WO�p��&
ܞ��B���K=5=]��n�k[(�+��z[ �\���������=ti&�C�[]�Mh��ۣ���AA��J�(��tz��/��4������R�.��ė/ ����]9Ga�Dt��e������fy����ʌJ�Q��7o_ei���̮af���Y�=�do
Bҥl�aw�J�+�)t[+�����f�O��`�U:����^�~�"�*3b.���]���,�K���!��13��8e)XX]�l�����_�Ӷ���p�ేmwo{XpL��.7(��So����L�I��^o�3��8�曷o2����d�_��Jd��� ����7?۳_���?e�Jr��fۣ��w?��=~�޶6�
����s���~���ŗ_��(�U�C:$����e����8H�aA�d9����S��g.iƺ��Rf���/iC����\(_(��ԓ8����F4�.�q���Zf[�e^����oB1�<�>�7��bU;%K�My��r`R�8=���
��W�P�Z�Q��n���+>t
����D=B'�:�q�cy��m߬~L��U�g�)�z.kHٻ��e"���0z��I�~ӯ���������ƙHfb��cd/�$�Ak�cz�)�^j~=���D鿷��6V��-Ҹ��R�z����� x��LJ�*Y|�I����e�B�VԺP۵�"��aX�O%��d^�E��,��B�x�07���P����|�
� �L;=�1���9ђV��c�u:�{�ԝwTdA�pyM]�v��!16���*`�9��/����Cb�!�D�\+j�z�9�__㙠I�6.�q���|�����B3KW G��li-�%Q�q�!U���B��2$�Q��t��D7�3��0�1���q��{el*�\*�r�1�yW�#���6�5O5�����x�,x��S �KuL�x���G�c������,�8��v�Q�l3N�Ǿ��z�6�?
m��7�֩������-�4��*l�϶
�� �tp�3&R^����|�������'m���Y��;��3�4NGXͫڴ�S��'����ߚV���J�m,_��s�K���^����@�/�Yc�o��*E-��A��ds;J��xrJz�	����
r��>�½�����1�Q�::#�'�]9��d���\?0Q�H�s�u��������Df��"4�}��yyI���/��.��M�*��o5|٦Q��m������>�:==��������r�vc{��!�N�L���mأ�Q� ���!6�.}v�>G3���|[[]�m��Y�IaS�y;k[�o���3��� b��GE�D�'Z�G��۶ɨ�#
�� �d�8�E�c(XC��o2�hxh��!�����m�aG�n��w��~���u��&�m;�G@3��F� �{��9�P�`��m�hi3&x����
����
 �
nn?l�}�<��=x�Yۼ��ݻ�|�X��������,k�l�J8�q*uѭ��8�*��^P��H�Gܯ�~q$�����O���t�=Y�L���3g.uD�.�D�~���>JEk�2����f��`�g"q�~ģ�U�^�~�N�T�;J��w�s&��w�!p@c
!�e��T���D��e,�{��A��U_X�)y�8˷\ʷ������;�TҔyh�([
�*[�WU.�tC������\۾�����?m�_���ㅶo޹�J

�V
->x����{�t��ۧ�1�mӋ�yv`L�Q>|��]`���i��{ld�B;f���K�93L��P���O/W9�'���J�����>F�Z#��6;-�0~�ճ�{��Y�S�!�^w�^e���2�\��{G��\8ئ�%~:��	�'�N�p���+e6-OXߐ�
?;���c�]~�pOٗ��֊%����n);F���e�V��C	|�P�W���C�LE���+�<�����cڣ��VE��߲���|�������g��.i�,?�#��ҩt�͋�J�䪚ݪ�Y4]^}����{���L��}���x}�P���E�P�F��G�S9r
%˺K7��G2ذ��6�c��r����56�v�S���1�>����0��ڬ��+�8�"���i�C��Z��� �t@*��V*��u�+����p� �@�ՠ]��+��O��ֵ���|��ԮKDW�[jq�~��bWļ�92� |ѯBr�5R����Yު_��g��=gƐ:�H�:��ȈDۑb�d8�|�<Th�}O�a7!O#�!ԍ͠��g��z���R��YiSskmz�Q��6��]�js��mv�^���j3s[|Ǎ�;���ʳvnްX���]�x��&�������vz9�OZ�=�n;(ƻ��a�C��|;C��^D���`���w.g�.�T�Br�e�۰8A Rx�J(=������B�o��]$��I+���wk��H�%�^��U�`�5�7�{��,IGB�bq�O�p)���7.��c�*	f��p���l����t!�-0�����㧟�W���|�Ť���z��@�S��ݸ5��C�RJ���0���^Q��{ �{�B��=f������<mO?�����rU�5�U)Y�y2O�<k�P=Fwsk;{��<��n��:	Յ���(Y#���1�.ɚ��$w��5�{�`�;�5��ٶ~�>��������?j�>����
�{�
4U� ��	�>Ҍ��K�I����4X��V����eY�uEHB8A8��.��c�I�fN��h����0��L�MC�:�9���T����Y����.o&��V˄��C�
�(��O��~�'����?�o���?i��'��������{�u��X�m=l��ڊ
vy�~[��n����ܾ�=p��'�o������j�@Q�n ���jH�5_��.����##P�*��Q�Ը��P,QR�3���LA�c�V`r��=��Ƹ|� @�e���$�BW�'�E��|PP&�i�N��YZ0n�UЂ��g�OA�K_r��r��������G���㌔Ku=|&�A�<��=WO�<i�^��저�x��eG��XS�.g\YYF8�h��k��#��	�����8r+�z�3�Cj���9�̣�3K&}�z�K����ia�s��x:�=qQ@mE�,������Х�J	y�
�.�vyy?�i�¡R��R0��(i8�G;K���+l�����g��`���9e��U2�2�tS�P����>����4�3��^=�I9,[�?�.�kT�\*��hc�ZEL\(<'*�[�J����K�%Ζ"\�v*xI�������ڦ��*�R%�g{<�/���6�v�=��;��������ִ	���>�@n�˭o�_�F�n��*�Efx�F^�y'� �����m`o����l-���(�ao����נ�tŸ%��KS-A�
�Z8�L�~��;f����80�Q@.e�N����Z"�%,񺆰\��@ά8"�2����m�t������6�t��YӵN�#B��ֹ����3I�6�a�a�V�%ԯ����ۗ���<e	������Nw-�
���r���/.����2gT��2.�X�WVњDQ�C���5�kd|��E�Zl�Kmrf�M͢t�x��n����6=�q��}��E�B��C�ªh��e�o���֮���E�#�X�d�Ӌ�\.|r6�NqU�T�.ޏ�Xi�Q�bG����}X������ՙ*�´L�b���s2^��V�(I<Ӊj����3�A�1n����+	
?�Jnu�����ט�Q��U�A ���}��o6�j�i�[8�on�߼�����V���GJ�1@���y��g[Q���op��|�v"	G�aN�f ��wgxL:�+���KBڂmO����$���!�3@�L�Ѻ��t,o��ٶ��k:i*\�0Q�Vf��j���W�G��wߙ��y^Z�/��g��#�t@��ʂ�O�RW�+ff(�$}vf�%�`ml�Ixg�gV�����;��q���i����(K���$/�T�ʀ��bf��'Է`���[��锑�=
�w�(����R����,xw����Hmz�¿�8;�e�(X�Khzڋ�<���TQKџ�/
hkk[���B����������)
֏ۃG��<=l������?��g�(���B��_n�Kkm���P��h}��ڧ���}�����gmk�q[]����(�Bf�_�|��BExTiP�)�P|ͧ>�=gX\j���� ���]�Ժ��VNE@���Rgg���A:LJ��/N�����{�+9֞B)�؇���.��>�i���z����bF̭���9W��4
�;uui�C4R;9<n�;{��˙��s��(LEg��}�� ���ն���V�����aK	� tK������*G��ϴ����A��Z��`�c�Ɠ�D��`&V v �CGt��i�r��9�,�r���a;<:Ȁ��I3GV����<:����T��J�r�d�,�䪄�/Pf����+�
�y��Qrp�˥;I��SJɷ�X�`��yu�"u�H��)t.uWѪYaqQ:_����2D�`!�K�U��'/*^�ۢ�5��}Q��L�<��8Kꅌ0� �;4?��ʩ�����S ���[�ϲ�1��VL�ڶ>�V�3D�+��%����G���g|�怈˖��Y]�րF��P���+ʞ<5U���A?���}�k|��&��c��ĭ�Y�.��g��+�U����+�^qfb���m Zn��J��\c�����[g,?i�~,&#0ߺ��v��C�DK�B
�^1���H��npwc����-D��1U��r�w�����;J��}�5=�L'��Q̌��Y#�������4�ɾ�#a��+$੃O�<���Ql�٢�'�HH\;0I�U�we�l�G�*!M���U
W�.�u]�kx�=XS!E�
�Dxs)��$J��
.LU;Q���ױ|ӝ�NM���>5U���ƖH{�η ܧa��
��ߐk��)�k�]
�bU����p,t��X�g�%JX�|@�� �Q:��g*Q���+Te��h�@(���F$�ó~�;�D<@+�4}���H4�H�2���=�K����nӿu?�7]�fx����_�A|���w��D+����M�����+o֡�K8 �G�f�*C��oU�rS#x
����:����.������Щ�eX,g�L�8���@�z5Y��)��@�ZL��pi�B���@�|���I{��1B�6B�J����r�٢�+��̜>
��,.�����k�Ƚ�I�����@@�a��69��ֶ�O>�N��{?@����om�h����>=�FG�;xG���KP�D�)�WX� tq>��B�@,�&�X�0��&p�_ᾏ�8�@_\(��Vұ�)
}�Bɡ�����f�������N��ࣶ�q��-�Tͯ�T-���9h9<c�k�!�jB>㳼dbj�M�̷���6�R6���V�dYჇ���}N���y�f�ye��l�h�V�e葸�~��	p�&�ǳ�X�6�^�i*Z-Z�	�Y�Ї��1�����[���{mED8e�!��efo<U0p5=��,@��?Ҕ	e��C�+�6����-���<J��B�CX\��3�px��BE�AU�P=��I��~��H~�����Sn.�ז�v/Z�n���ŔM8N #�����[?C'LUU��Q	��e��+ZT������Iϧ�QЄ�)�l*�Q�H7·������K�*9��rɝ��2cO��������T.�*����RH�q�s�l���=oz�S�X���&�2ρ�Rp#�-U�U�-u��+��%��%�**X�U<?��/�NZ�_\�>:���#�5p�;�`�k�~��U���2]�D1����YG��5@mG�o�,��Zi�L����`������5��4�K>i]���T�#�Y;՝�������TfU Z/����s�A\�(<��n`�H�WY�{���Z/��3�?�S'l��8!��I�s93JV.$�eEʠiX�D���-I��f�=��~��灏���DM;㷤QĮ�S�cQ�x�?e"����I$"�mCU�7S��h�2cG
��1+��y`�JI��X ˯�Ʋ�XK���<�XFC�L����5����_!���`�~$!��3O��;bV�7&~<K@|�M��"|���h�%z�g�+Z
X��΂:�H�]��0�:�B942A��qv�KǼ���ɢ���y$l١(O��`<���D�B�������t�:��߻�.�b��K)���!�g�6� ^��¶��8t8lx�@�N���:T���l_�oq=��{�6{p�҅����$=��,��r�[��j��$M����&(���>H����nl�M��:���ѩ�h��d��!��o�NUC�<R��>���*�'���ʔt�l�r`�M~�����Q��;_K+L%aT8�+�I[�f��!�Q3	�E�e
�W�`��Kz$m�
�p���A79wi����p��{���R��XG�|�>�����G#�=l���mr�}���W 0_�7	�|a�}+/�ӺY'i�ʐ�)���3�O�Q�xA����Ʌ?��}��wrז�#��@W����c5�jy�բA�#�]�j@*����kϧ-S&�R��C�����'1��v��L�:�wF�>!�p��%hu)��G������[��:����}����>n�Kk��D��x�\�a)i��Sy�RR/���E��<?�5��'�~rv	ek�~�1���([��{��ou�̀���A�f� h7 p������(�;���_xH)��#�02^Y�ME�t��J��-,�'�J�˺j��i�:����viT�㌍�F�%��s����977ۖW<%y=V�@eGE�7��=*rQ�p��,�5����A�p_�
��?�KY >(�a7W(EO�l(��,.-d�N#�����{�$�P��7�F�p@}0�������=��l+2V �0ox���
���l����⩶W5]|yʫ~��gf�j�����9��f���5�@t��!I����+.uF.�M�o�T
%�k�=���-x&-�>�l��_����, G<����"�-�A9VEL|Մ���jW��OTYY�� qR�۠�EY�,�H��ȏL,u�]�(�y����W�8��Q�q�_g��lL0�ct�/�QF��,�\�r�<I�vA<��9��\��/����������I���}o+}dqi1ʚ|�`H�����><[6뒲��W�Ѥ����cR���oeKy��_J�k��I<����5snBa��F�Qos��b�Y�����Dk��p U�1�vLzTC{�&��iP��-X�!���b���Hĸ#QS t�i����IFM�/>���<xE%ɹ'�OH[���rr	���s���ݜ�.qb�2z$�D��'�ySN	��x���c�z]3��*a$a�)�!ғ�xL��b�G8wٌ���o��a:b,�o�)�^3�F���JOR4��@��i�.<qqM���WD�|��V�x�@�(8�}��D�Bi�������=��eZ��u��a��w3I�Y\��\ ���~d�]�q�m�0���q��	�*lCѺ�!�L���G�\jmb��]&�"��)
�8J��K߷n
VEO5�%M�9;G<Uц؞S^�]��Y�$�2s�
Xd$���.!�?a�jvJ�`$��C��M�����%��l�!���u;; 2�:��=�i+/]�9�(�j� >m��3�}���W�#��5]�3ܭ��X�"��7Km;��5�!��d��#��	7�#�8��Hbt˔O<,%S{�����G�I�Qʪ�}�WJS���J�(�]FI�O��p�Ha6�"�X"���/� p�#��>�;92(���$����\b!�U����f)脞�}g��c�D�f_��0�G-�]�t�I\G����+h������
�,�nȖ���]��1�?N_>��Д#�%��l{��~�����}�����O���7��=�R��ҷ���I��>a���&#�2�Kq^00\��Z�G?h�RUK{
�;��̂���ѹնL>���>�Ώ���i���3����ơ%F2�径Kp�Z�M�8c�"���I�c�sT�:�M��&���J�|�_����5����`����ρ�ӈ0����{7��k�[G�Oѷ����{yt�.OQ ������ӯ&hS�V=����g?l�����r�ڐ'��o
�-�҇B+n���(�\�d<��=��t���z�����Ǣi����6����=��=�����'�kK��A/x�<;�pϫ> (�q�x� �4al<��߃�c�*iˈ������-J1�=�;>9�|��Ig��Yi���z�8?>n7�!�e�*5]�ݠ 9KC��kmu�}�����|�}�?l�G?i�'?m�~�i[�XoK(rk�Ѕ{m��6��3���=Fڵ'� G����3h���D�r��B��R��uO���]���C˨�(e� �c�]��#�/ ^ًI_���}+A���9�4�ڧ�rt>K.��ې�.����A�GhX�=��4���+�FN�:�U�3�Z��2��e<�i'�oIkBG:��Ix���u��#�gq���|ߺ"�hi�^�	�HQ��B|���!i(��4�Jm$��*�a���$���R�ZXj���{��UdiW�-��	����V��x݋��S�s9*������"	��CH ����ʳ'3�Jγ-�9tֱ�Wj����u�YZL����� b,���ax�@�J�KNQ^T���TB��"�iNx&��v9�)O(��X_�m'c(i�%��ن��3�C�2�b��|;{<���Kmkۻ������ͭ�����Y���iᄻ�K�﷏?����'?h?�����G�?�n{��;W���|�����ɣ�b|��@} `_�1v��z��r�(}\7'�c���T��ocȠ^j.�r��dC�Vi��a	v�k�W�O�Z���6B�?�˫�k�k��)�K��re�O��xԌ�3Y"K4l�n\z�I
��խ�I��"d����	�I]A���ru.���-�4�]��G��r��9��(�:kIM�M9�pR��s_f_�u�;{WN�2��I[6�;��無�k�۹2��W���&B�6�r�B���#�>�W��3��{��L�d�:]f��B�{��K�I
sh����X�X�&���m}��9���U�d
�fvʻ̴uK��)��ն�/����>w�3�o����t�wR�c�Kg1��N���'~WlS1�i�X������~�Я7�����q�~�/�}�>$
�χ�yvi�W�N�����%N�ߚۼn�f�� n!�~�-/I�����)���RQ.%�]��������^���1�c��G��%Ͻ[0Z?(�8�숴��0i�4����{��Oד6�T�k��w��Ç0��msk���/BgƉO�oT�K�>���&�)�-��ˁG�^����O	��~��������K�mck&x�-���A;3�p��4	�4�q�7K��!�e��Hp�� �%s3�}���׿W�[s����`�۬��^��}�٪��\��Q���}Y[G@z����~�W�[h�<����d�f?�	��M��
�����4|��J{��b��zb�b��_I�˙��L��E�A�X��ѹ����n+V�O��򚝴��T�.�=`�m	���K�(p6�!gP��$����w�z����?~��{���������m�������G�=}q;ta:�h�Ԍ305 �}9YbU�:-C�0�ʒ�j��1e�*:$����^
� �iy�OauD�^�yӞ=ٱ�n�,��B��Ni�4׺9��2"�e��⌶�
�]0�ty����;��~�au��図>(ig�Ǥy������hGi0X\��IW=e��Zr�#��V�	��|�AFi�t�	��+qk�CM���ڜ�Rѯ%�X\�8|F�B�ŕPd��Q'3:���K�TS�FHwR8 ��\��HZ"���APʤJd�����x'�|%K��1�mC>u~�-��$���ƕT��|��Ň+�2w;������n���`�x�I�,�|`�����ֺvss�ݿ���ۃ�Cl�ߋ�����ѣ�駟��~��������?�A�����>�������h9�᭡�/�з�a�Q��;E�F�E���9r�a�<��a�����ZiW�dIw�c����ѧK��x�lUػ1°�{�6^�t� �N�"ZIl��P`�y@c�E`�)t�8"��i�mL7�f���K�\z��:M�Η2Z>lF��4�֝�F�rV��s��[�X�Լ�A0�ʿ�z�B�sv�yF� J;���a�)I��m[�
�h��_x�vL�,��.S+{�h9åruk��b�ܧ��ޟ[�=e��В��0�4���y֒o�0ଫ�%�@]S�~�׵6eu?�u�(�#�*Z��9�q�`*^����q���u�NqǦ}:��x�U�|���ڴL��mR�m�t�_j9W��̝8���t��΍��2� �;��&��M��b���>�{~�1�*�����B����t�~�T޷e�t��f{�+WN��M�o�O���]�"vQx���Ǫ��pw����0�M��K�.lN:�c�p �ש'F���e<~���� �Q� a�2��c��-y�-I_I����D-��{�m��g�]�b��=�o��.F/�X�T4ץTu
���v�m!D{��_f	�F�u6���`���o*z�^W���<�e\ۅ���t�����myۉv�	çy��T�Tr<��y��
������{��| =yN�f���n���f;|����;�A�g,�=��r���3�K��/
��t��[j�ݝ[�@���i��'��)G٠p޴L��c	�r�z��=����M?��y�[�&`�-7H��>�w;z�Ӡ�_i���]aqq�}��G�G?r����?�Q���?���1B����ʲD�)g/"8�L�
����J��-t�^*��-3P��!��N�Rʹ��*j������|����/ri�G�{,��9xa�������|��F��?��lI���({��{h���4����@8v6+<P�<(��篮�I%+�_���el���r�:K�%���@�5��Ҷ�)����4�4�Y;gpU�C�T��<-�"��n��
gt� _��JĳlR�� 3(}�[�{�����G�o=��,����e��U�Omg��f��g��*��Y�b�(ȿ�O��I�Hk���Q��SDЯ�፸�r��gk��Mx'���:���}(����(���S�_�3.C3VW<8f-|�A��͍���ݏ\�C�z��G30����G�O�U�������C3���lR%����*bBܱ�zglqY�X_l�cCğ;m �kif)�E��ȳ��ｩ,Vʖ���؃Px�ူ��B�5{u�`iEx��b�+�i0=��n��lN}�,	��I!L"�M�H��J)�I��Y��!��Ͳ*\�/`�Se�Jܰ�%n����K]
>e����Y��S����Q�]�|�	��X߉չ��QUj>��{�\�&�� e�q��{����^����i�R�����Ehk����*X.Y���u	B��;�\B�٧�X�k3+F��@����	�^?�df�Fr��K]��~`��L�g�F�Kb>������g�e�� R�?0g�+�����?~ɛ���G�U�,���`�I<�͟np���L��Eۻ�T�K7Ow���S�B���wO��6�_M�3]����;��bsk�Y�
��I~�gO��X'�2��pT?=��z�Wi�n<�i���c�M�Y�nt�������>�׋>U����C@!��VyЎ���y���D�4kT��j��25�8\/U��G�;ף;C-��⎂�Ǧ�
��K�@�҂�J�����?!([m��|�2��O�ґᡱ\�� 댁��E�"/s �
#5`�x.w�)p�`�������*����,Z����E�|����Vi.�_��}�=z�Q��3��(J���2f-��IQ<����x�8�Y���τ��s�cP���ĳ��[f��3�s���C0ּ�����ɧ�Q�+
�q� �)X��ػ{��C����*P����\M���-S��p��wp�h�{�gD�������[47&����a�|yy�MM�	�(�I!�N���*Dk����*�J�}q�����sY���'���-��n�O�\	���߾����W�W�/��˿m�^��~'��%�Ԭ�H_.٭��r��
���8g�<@cB:!<�<?/e��~k�G̿w%�ʕJT)5�;����]d��	�gi�hW�*��Y`�j���*,�o�%����U*�Z�t��� �m�=���M��xa�S��LG�p+#g��#�U.����r������?������������m{s��P`��;	/2]�nʚʗ�K}�g*W����;-@���Q�����|�d�
�z���T��xc�ս�?ϑ��?�4��ا������x���-�}u����5��Y��Ԭ���j�.��B���(\��R�Ƴ�o�_���(c^x��&=(P����2h5�1�l�c�����>�c�W�W:Ƴ��B[����Z����%'h��>�&������&<h�dY��a�Vq��V��a���#B����&���ق�,*N�c���F�" �p	�k�ʼ;@P�[�����:Y~B��D,,�H���pu���:�1M��G�1����f�����!������Փ����+����w���{b�V�����~�o�v`vI'�U�j&�6R���^)+�QFWFX�|��(e�T�la/��#W���:�e�.#t�k;	g _�,#a�c}ע`�������X]M�-<#<|��-�5�;ﺱ��w�A�ō ��L��;�)n������� �v%�ӆ�5]�|�p	4x.�t+�_1��w�h��r�^x���k��Rr�M>&������_�mE��҄�x���iCo�����* ��h6�>��I���~�_͈Y��n~�+��p�O^��q�>::i�߼mo^�E 9�޶��q(�w�P�]�߯3��cQ�R��N,q7=vp"�w�o+Z{�����]X�̬�]�[��Q��FM�G%@�����L[Z�l��e�ݦм�X�ꆺ{ߕ6˓�h. ,��#�
-.YQ��L�>e9c�nK�%�e����7}�	o�ip�6J_�kd<������=x�>��Ǫ��7��(�,	���D�%3$��mւ����p�8����E��Zv(~�д�?��Pd��(��F[Zv��88MYƨ�dE�e�������uÇ�5}�5"_�0��d�`GG����0��~��a��a+�tE����d�tjff��"p.ʹ�Yp f�sSAs��@]\Bl�H�����~���,�k5�g���]SIU��RaObt	��L�,���� �6�=L_�����f�]�����o�������o?��ߴW�_eF�ڨ9��,�V9L�Ijiq��!8{i�G�;���)�CQ��H8]��JJ�5�W	н�[ʕʖ
�������{v�.N��B�	o.9T&3[A6���L�S��*/�a��>���6����9Ț*(�[p"�F�S4��W1,H���]2	<R���e�6����O�������(Y�]��?�	J��j�����~��}N�OPHX�@�ԕ��_
\͢:8hI��2h�V)e���.z������D�%�#�ۂ����CL���Й>Ϛ�1�m|�j�#(x���˸=B�-<���'=�Be��x$�J�kcC�j�����΄��ݻwo�"�g��S1�LNR4�h��S�X�K�u?�Û�n�Ao��w�ԇ���W�)Y�>�)�(X��u��.����_�HR�[S�;��]�`&�|��N���OONC�\�-��ְv�C���~eaE�>�ȣ�l�f�zA,�5"z�*�t����ܖ�L��VF������Pl�̨u����f��{��_n��Y7�u6�Zr����p���ގ�6U��q���/�	�ō��d������z�����)��w��Nr���{
�Z���:�����u��t~y����?�R��8g�<z=���0g+qI�-*~H<kA!�%��aӲ�^g�ӭՏ�I�2TK�t���3�e+
��5+p�\�޵�����}��&�r|������~�P���b��L���ꕤ��p�t����(1����ܝIYI3���A��� Z�W�.O�Vr`FҨ|�W*�Ў�F�k����6D3�d�bD��M��=ES�Y�[���Z�z�Pj��{�'�S��!��S��M[\�k��ˈ��駪�	Nd�ʃZď��O�km��:ʊ��6wM�C���[�����$�X	X2�k�c(ZK�mu�~[D���8c�0�ؑ�	G��ݪYjk�LV�gQq�#�&����iS��V���0�І�[ԯ�Sp@~f�~��9\XZl���٣��������=X(?
�If:N�X�iOåy�w��̅�߶��*G������)g�)Sּ�?ze%�aiEk�M�R	��e ��i�w�o��es
�"����R���@X=>i{{{mgg�e�����i��Ǟ��������)�7�+��2d��)�'y#�^!�S��L�J��w�B�'x�{�T������ laE���y��������ܶ��>�ޏۏ~�'�'��O?o�[��w��|������ߵ�%����?��{��eY��i�p��ZG����,��%�fM��g�^�L�����)��͛���õV�}?����+��X�M766�0̠�7_ݶ67�@x��
����O���"��~��K?|�֖���*��ˮr�fA�l���V�c��cx�篢p�f��܋4P���O��R��(`�Jܖw�U��((f�#Y�^�RiJ9��$\��6���<�ի(W��$#A3�ʃ��8v��-�rX�'#�tD�*P*X?�����G�������������O���j��(u�!�����	����Y[Qɖt��3nY\`,F��u	��gp�8F�-�Y�rVc����p��KY�b�KZ�Ų�� �igg�F�a^�����J�״{N��	����J���^۾����@w�x�{��������^̕��k~K�pwP8�#�U�!��S�ɛrNl͕�'b
��T=�N]��'��:/5'�9��h+k���J0��$��tąސ#|���X1�CcA�cÓ�Te�U�:� AU���?���/�v����a�]����,n���)�0�9~Ñ��#x�H��4No;� �Y}Iƺ({��WJ���M��P��f�~P�{v���vA��恅��+�6��'��	�g�P�&�)�&̜�W��{��v+\����S~l�NQ��f�ݛ����k��bU(Ƒ�������;���{�ȐK�*���ꄿ���!��7��_l�k�a@�oe����0jxC7��mY8��mp�˿�T'���տ��@K�0,f��0�����ř��_���CR�?4Ҹ������[��i���,�`��Y��.K\��?�Wy�~�����*i��
�̸�l9cW�/�K��o9,�t��p���N2Hy&"
���q�(n��g�T�g�aϊ0�,�u%���ɓ�MM�OI���?zx�}�����w����Hn���:�&�"��]xi
S!��8�Rv�Iww�fhk�Q����ߙ�̒K�^#��v��㶸�'<+	~�WT*-ǂ��6]�&]I� ����qن�����?�I��|'}�\a<���-�g@�fv�Y�{wۭ;w�<�Q�XzT��~N�@I���J���u��Y�ڳ�<�γ��,��Fqh���@�%�|�K?�1���2.ĸW��b]�ڦ�����aW��㒓�����4�~��U�+H����v'y��s�:��p���oY��G�7��M���b*��;\�:F��7Ȃ�G"���������oLH^��g���㼸fޛ�����k�P���g�|ޞ�?kw�?l�?������g���?����į߾n�~�M��o�epow��sVQxNȒ�Pvo�{p�^�w�N&��^;V|<��-�~Ēx��N����v��(cK;g�|���]������bf8�8��m��:�I�Z��-ziQ}h�Z�Ү�-�>����ͳㅓ��M������L*����U��'���=kO�>D�:��X��;�y©�KGʀƽ���.Ǭ��A�F�3�Ez%����M�g���e�xu,'c0��N���|���3q�gF�����ʄ���*��R�T�J����4�J���Zu���
ai/�ϕ��
��ظ���5��>�v���"�2kU��Ï����>D�T�,g�aj�z�A�E/ҍzN�%4�:2��+�ſ�i�'VxV��	21U ��� 3��B�� F�!5���g�Ux?�8n���m�j��hG�Y�(Y��hGm�߼3���2>�d��=�%<D�Oc>���ɇ6�E�)�JK��6����aN��J�Wf^ݞ���9e�9c�py�������Y�FAܸ����+ L E���:*�U-��S�rx�oN�`���2C�ʚ
O���T�a�tLڇ��zV����V'#�@���N�a*?��(qӖ
�]Ƚ:��v���s�l���|�=6�_���	$��r���_�%t����1�3��2�ŉ�z4o=����*U���a:��w(9��7����rϣ���?3w_���,��|����+p�q/���L����@$?j ��,�x�冔��d�g����fA�F�Q��O	=�u�t0��_2�\kw��l�<{ܾ��||���2߃.���>�fJpU�,�ǢV�T���_��7�\������*Lzӛ�ϻBp���|Ck��OU�Ey�v�*�3�#��p�W���D��K�	D W�*�j0�G����=o�-k�������e+�+Y*[�����杁M��$~�����k���o�J_EiE�����]�['�L(Q��ǭ��h��"׍��6J֭�w���ګ���\v� �4�G6�Zgt���Bj$�j0|pR�~~�<b߭s'?�������w{���MM���ecE�.�+��8W���J����'�� %k�`EL~b\>��x���R�q��D|�vN'B���g�}�~��_�Ͽ��ݻ���PW���{��'(\_|ў}�)J�=��zV>v�wQ�vs[�[�"�[n�.�eSu���N¤ �mx/��tow��Q����2�&ar�J� ��B]�ȓ|�j�
��a|{J���#o/��Є�x�V��(�^��呆��Rl����^���b��ब:!͒��n�(+n~2��<ݺ��� ~I�z���r�T��۠?��T�\�R�T�NUN�'�KR6r�A��	�ɘ}�bU+W�j���5&��c�L�b�3��1����[;K��t��3T��W B������&�9����1��Ī�	�0 ����Jښ�<�կi%+H�#����?�9)��$pA�U�-Y������F׶�]R�QI�9����LV�B�ᦡ�H C�v���s��8��kv�<7�@6�D5��p���,4�Zb��T�� ۇ��_�%`QRV��V
ئ5���Ì���\e*��Oj=�@�n-u� 3�`�$��@W����|L��� Ć!�� 4��vy#��pk�ľ���G�� �L������C�����%�<����|�Gei@c)Z�I^��̰�b={��fpd02��4A�c�~j-4��3i��+�,�4�h8ۥ��7`:��d��e���w0�����ٍ�p����5 ��6n7I߲tg�w�/�,�X^�E7��GLp�����;����ҫ�W��L�5�\a�{aG�^)#�iLg�%�{��b�v?��s1�1�V�M=?�3�r��G���*���5g��r���3�0Q��#ظ��m�*}
=���%]gKߌ K���;9��٧��p�N�b�򆪿�0���X%k�(ci����P��_l<&�Z�z��ϵ�X㷮�~u�����v#+W�����ݨp�`��.@!���wœv��˴/9[?��.|����y���bS���J�d�M�������!V��s�nf�gc� ���P`Hs��T~�r��,;JV�����I�(�+�_ƨ�n:�gBB�š�q�x���/Ws<���  ��IDATt��l��Aiz�V�*�o�Ӓ\����'E��5C�IH�O@���sʣ�ð,�|!��<-���,N��k�N(�w��Sס�dt^K*���`����R����G�������>�sI(*(��7J�Vp�/[��9
�]�����{�)�u*C���4]���$hvwv�>J��r~p���NV�wM�Z*U��*���;��fL�n1����~D�2Nx�[Z5'Oy�gb�/���! +���峾5�}���,Zu2V�,3�.܌I����*S�n����C�󂎛kk(���%���\��+�=��h��N���n�yYPff��v��_n��g�>���`����g��m��j��)(�*�����>U� 'TP� @c>ֵ}��>2ƪ�Q�X�C N����-���ʭ��&f�^�^=�Ŭ��π	\6����is�6u$�Q�E[?�g;1meU)��~��J�(ibF�?bDb
|�4��a�]Ă�P�i�0˨��3��B��E��K-Iτ��Ҫi��_Y g3�I�� �8�7��*L��J%��P�h;ރ�S�~L�Vn�Jx��������[�N�(%.].>%]�6�py	�>"������]pP�������l����>~�7@�k6�TW�b�b��8��7x�"�#�L@E�-��ˇ !@޿������ϼ�U0���+\}GÁEz�m�bd�r����P�-=����r��E��4�x_�YM�ÄV�]��t:�v�0���	H�8�G��\�awz�ψ؝/Č<t���*H=Nlʹ���(?�&�'=��lO��&ܓG��ʿч�7�{��T�=ωM��/�o����l5�Q�Y��:X��bԴN��.�*�0)C~ݘ�9ڟ�1v> T_wp-0}�o�ZZ�@��ik����\]���������G��W�V���Oc�$ 2r���o7����� S�ZmF}�<�� ocK�n���W6�f#~~3�����2� E�
y���H���u��?�f��������z����̨��U������oΗVVr)�[��B�so/¾ۏj{��BC��?0��Ǡ�wC��'M��θ�N�C���_�)�l#�F�Z�!?��[��#�&������jK�����O	�����1xC ���ا3�K�>_
����HY�Ȏģ¥Ʊ�t�R�c��Ii��F�dL�]W� @�Y����67i�3ș�[�g��Ӻ��4�G��"k���\e.<I�L3�,�dk�T�
��c/�k~������)����ʜr?�\^ޠ ��%�\fd���&�n^��&��Y/�ݭd+��
vq7�31�ʎ�� ��N��V"����M0���T�7�몓g���.�R�U�틤I��B�b��w�*�����%��ݻw'�:ܾ{;�����)Yǳx~kѳn��W�N�R�-�#Z� ��z�I�lC�K��d������ƪK+,?�6�в@��#�0����X���e��o�U[:%�ׄ��깶߂M��ʈ�;\\=�~NĚNd��=��d%�3�F:���mVQ���S�-�BhEq��KqJ^P�u��z5ސi3#���@U��^���0�A�
	NW/b	 l�=�f~vqbnmq�Z[]BXqv���y�f(��\�|{�#���������z6(�<����R{.��bW��]$9����8��s���p��Ն�r�g%dg�p��8��!8����vt|֎�;;����o������o��j�J�5�9{zH��EŁy�rs��Z`�͜n�v�}8�h�����F�8^G�pG��v��������N�✞�ig�����vqB� i��%] ���-
�:�g������D/�_���wg�t�	���7i � i�w;���m3'�)�W�����H�������URf���^�8�%]��f�<B9<�o3gm%q�q�b�6ic�g�T������A�vvخS����m�p�����a�����8�<����ͣP^s��V�\�AΪ��G�����qv�R�o�3ma��f��sܮ��q�;O��%�k��5h����E�]��S�������R�A��,	�a�>#���]B��������7�d�8�5�:�U�|��2�!J�,��S�M���!�b?#%�q�M����2:��)�gm��7���K���`Z��z�.�k��L[�W,/�\�|�AK>�p}!}��������kfs!�ٙ��f�]����2Re�^]8��LyH���|i�����9���.'q����k���Q�_�{(V�~�U{��(+w�(1}Bϗ|@@�[p9�N�&�0�d�n]I����H���ԣ��n�m��)��_�r���&���u��n�|��V�_��<@�0� ;���tU�-�s��x�,�fH���S+oMj< �荏���U�x[gB�3`�����Ԁ^����QS�?u,���<�-�ɇ �B�m%k��J�j�x���kیy�tx%	��;�a�r��w��t�=��-�>��G��V�J��|h��,�W�V�?�����7���fx����5�#,����@{��Nc�r���ɫ#�"�[��	�||v�N�5��4x:]��8J�Sx�홓����l�R�F ����k��v�sӝQ&B�'���ݶ��ٶ����<�>�<�-�.�����*�<�򇀇��S�N�#����݃���z��o�m�|��m����Q{��N��ԧ��v|>û�m��SW����m�~�$�o���~��,|��D9�����8�m[��	���k��L=�,��ԇ�v(�g�SV���.�;���~��%tH��6%�<�v�5?�΁BY�墽�Ņ��|z���gɓ��'������\��9h�{�iK�1�z;��3��"H�Ƨ������1�[3�{¶S�TFp��d�:��h�9v��0&-Ck���������v��KrlA���lyk�'�r���[m�zP1=w2��lk@��}sV���o��ݥ�֭��}�e؆֕�)2��9D,m�Ȭ��`��Ӗn��,���5r��<߱<J�uI��z���D=�P�ζ��kre��Td����w�*s�|���J��G�'�,�H�WYH�U��%I��xd��<�G\��pBȉ�����D�_�|$c�,r�g7�iw����6�*RN_��O���[J���n'e�/��w�8{���=�<���2�/�g8��M���'F~�	�P�J��������Z^�BPg>�$��Z�gè�Gk]ZL��#L�a�4Gyb깿I^��q*�?qT��,Vf��娙g�2���4��^.a�i*��l����O�g~��(�9��	x5)0���'�<�>C�9G�p�t�����N;��v�t
N��w*=�Z`�(��v��g��Mx��Ļzw� FDZq���3�p��,�}/��!�����dE.���}��aH'��
�r�����	��U���/�x?�e��=����3 glל��-���0V+�J	-L��mr,�&6�:����y��I�n�]a�ք�?
>m�4�?A��]ӻʵ�y7SΉ鈤	Kzѷ�?�I�2%�T�(r�s���ղϻU@�n����x]������a�+�<$��Kw���j2�F�♺£�M����0i�g���a�����v<�-��q޽u�J�i�H9�128�D��)�B�+S8��Gn/�� �h>�7E�#�����+�a��.���X�#��1�b�[c���ɛn�v������3��0�_���:��Bc�hs�"��"�"<9�9B����5�z5�'ɑU�����h}�H��[��ʏ��(��V�u�m;W,�g_O��ת���L�d�?�B_}S��;�q\睫}��L��o���O�#�{���
�u�d�,�1����w~~�����
�ֻ���P^|��"W��k"*�F�u�!����~��Hxp�b���^�y�~�w�����߶�o������/����ߴ��w�ŋ��M�l�Ɋ<u�`�*�Z���"�h�Y��Y���l~��ܕ�ms����9�վ���9m�T>�	h�	��}�I,��v�}/~���֒߄��M�m�1F�:���a��ۧN��N�����u��c�N�[���S�爛
MAx?
�%p��W�{�Ql��[7n�r?�{���!V�`��*������
4�2nP�\o7r<�Ye���<���a�2�<l)���5c�{���E�g�9�`}+3���U����i�gz�btO�J7�M���J��?��@{:���yd<���C�ů�T�aFL�z�NnX��U�ZA�����f�fb@�*٘Q�
;JX�/�M�`�_ppc�n���E7�=�R��4	0���ͺ��KK������2�o��2R-�i��qE�
�n|'�Jg]�8>�%v��S�ĭF)? �]=�e��:����DFB'�>�I��z=YH��^�ƀ{CM8ߓ8=F���u N�}��t�"r���b!��EA��Ob�v@:�p�[p�=���ӣM�]��>o����Te+�2��K{(bS~�Gݭ������o��C�v�}���v� �9x�	��;~�y�}���wqZp������ �^��2���^�<�M�K�q��@a�����{�aw��ፃ[��U���ϭ�*o��:�-r��,�QFv��$�Ц65�ۡLޤ'�6&Aď�c��K�#_�9�2����s9?2�O���1��U�0�#�'}*�ÍbL3Nk͊�bu������}Ӳ���C�V�!y�8Ka���̣7"93-�R`�M�*Z�y5(Z�Q�J�A��7Q��aӿ��&�6=,�'f��_I�桍w�CMҘ0���g�}^[g<Y6��Bwxn�Z�m���,�s/�PacRV�����j3h:�d;���}�(��mMf�?��~�س>�sо)(D8֨ D��8[�i�������^��#/i���2<#T�W��IF���8�o�� �0�z�q���c>��:���)�7&�+}'x�]�%�����W|!g~F�c+#��ho^>^��ׯ��c�a��QThZ�͸�pN^n�D&�>w���*�Ӭ:��m\]Z_�����_��_��]%�/�m���վ�����wߵ���v
?���юn����,���:��Y�Q��__x"U��{��n߹���y*��O=�Ÿ>f.P���vF�Ð�*���V�� W\�ۭ���*
*�����u�E�m�*U�;�8^�fƋО�_w2�������|�旗QFyW��#��<yâ��
�I��IG։7���G�;�u��<����A�~X�6&}[��Ҧ����@nƷ��ߧˌG֥�J ~��n�G�;�f�W
 Ҽ� 
&#�d2�ӑiF�0�A�3�{�G:�+(�"�I��V`~=�eL�x*VN���.�G��uQ�q�T������U2��Y�ζPyH��z3���N볩D+!7�*��i�siv���� YM�����T��l�f��%H�6�H���c
Y��3}�4i����4���4��Õw�����s��լ�d�
��e��􄸂s�����f���w�2u�"u�:("�(NJә
�
����W�*���dU
���P���Pbʯ�/	s�CWf��P[Ŧ��jek�c��1y>���@�OH��h��0oc��o��v���ΰ�֧��Nߴ��5� �xwv$���p���6?@��+�)���r~����&�	`_���M�{���/�c����F�;���wJ��D���[V���嶸(XCْ�;���t,B���d�Ğ9�1��5�:��dd^�z�~w�>?Ô��Ǧ�0�!�A���g�����L�GA����^wg����?����	Ye��T���PZc����GZ������L�����X�3o~d�׽r���@�J^���z��\C�ZBɢ�HDq�vGW��W�ˠ�@h�*���X��
��?�^)��Z_����Oܭ/ߧ�(g�o�U���wNj��=��v��|���߷����g6���1�+����޺���߀�2䂘�o�i!f�6�v�O�a��MѨ�]M�����\�ZXXwԔ��4��3άX.�w�Ne�~�ė��C'w��;w�׫���&��x��������w���O�{����N���V{��E{�����Ջ�����0���D���v��*�����<�V� l���S��㶿��R����µ���p��z��}�ݯ�wϿio�_�|��������I�C�U_^���P�����.�̠���@>�tE�����{�Px�
���{w�M?T���p3N�aW��E��AeJ�*�y�� ����^~����> |r�-����~Ol��`���dyK"mO�"�Q�M�t�c����s�l(���V�e�$kW���i��"�{�{v@X�Y�X��骼���O�Uł�W~(/�S��v
���e]m#bO��_'��W��;�Ɔ��X�O�+��k���w|�= c]�z��5���!�Y�,\V?Q�8�d�j��_m��g�d�#�id�q�>U�Nh+wӮ�O��I��cR��X�}t�7��L� 2��W�lfV��h+,��U[M#��mm�T��W��Z,33�Ǧ*�CԳ,<��"�mEv*+�FW�Q�����F�#�lc �`���a-S�Gi�I")
����ʤ�V��Z���zD&qM����N��A�Am� ��%�d]x=�[��־l��-}移�c���sJ���}��w�g�խv\�l]����Ļ<�}�*OW"��P �KP�:A���j��8��.e@a��)~'�J�	ʏ�(Q��H]�D��4����W(`(V�/�d�� ����#��{>>�Rf�
���8;|8M�;���u8?A�;~C=��KϮ�g�S�e;����p��Ͻ�{���m9�&�]���և����:���Z0�b���V+mBI�E���+h2P!���7է���0�*��m|�0DH����s��@E���s�p�q���Q��T�����'�U-��Q]=)%����I��H �����)W|E��g�T��%.�פJVȒ>��|��y��������0Y�w庠�f/0��{˫m��E�P�D0�:�t�1ևѵ����6!y����+<�K�@��ق�RG�W�H�y��j=uE��1�'��g"�8���
�4�fR�ғ�O? mlG�F�XA2���Q ��l�l�t���t����џ<��C�
��(|M�4~h�[��72�#|eA�=�r�L�K��Q�vU�ӯ2�]H�.ʣ
�A��`nߺ�Bo�\C�I�|4���P!���O���+��E	�|c�Yaw�m�}�޾|�6޼�6���ҟf�jFĝ�Pր]�3��N��2SϮ��d��a;9���gԔB���~c� pǌ8>k�G�m{�lg�4u�Oe �Y��FG=�Հ� {�R��eU�|�k�����V�T�Qd�C�Q [X^�w�T�n�h�����*��?�^PL���67x�<t~� J�j��>��o�<�<*UY�-��o�y��7-���K{�(�I���*Wچ��x�U�U:�.*� N,�9!g�;?�-�(qԭ�D$�z��7�.����fI;Q�}�W��샅J'��ȸ��
�9g��#��6�I�M��(�U��:A�t�jTQ�-w��h��~����
e*rs��A�B����F�
W����Lj�W�/T�o�:������'�
��(��	Nɧ�x��vU/�����1�}�-�g�����KEZ%��L?&^�_o+����¬�L��&�'�U�W�5UIU��0"��J�r�7k5q+Pa��BU�KT"6��k�~'~#\n/�c��*���r��3�������w>ޓO��U�"�Gݖ�%�#|�����W��@т��,օ篎a�����_3��V�u��V=�'��	v������9��ClW�	�9�Jw�@��ֶ��:Ômr(tn��]�T�P�P��P��\�>?.��-�n�l��i���Z5Si)��(4G�('�(9�(<����������T�@܄E�:?^�4	*P/�P�P�����d%��2
��6ʖ�M\H_씼���D�
�s��)�#^��ݼ?�|*d�n��mӞ�Ќ��\*Y3*Yϴr%�qc�~����͛
Z�e�Q����3�����V3��1C�I��1�q��<���w�$R6�@���<S758�?�7}ۉ����ɧ�)c�AƸ�;�.�whx38_��}�0�Ŕ�t~�H�K5��7W)���Ǹ���-�zо�k�A@e�³n]g�%�!�C�E�p-���������4i7�!�����X�U���W=�vM��c��D+��81�u@�1شA���-�?���:�j�j��N���-㭊	t=;c,M����7�C��+�>O���8[�g����5I�t�11������P:RȮ�}��s}0\�3�t��hO+�a?�W9��ǤJ�#M��b�*�Z�V�sŋ��T)Y�^'�/�)���+�+�q�w�=o�����w�>o������~�P'K�Ve6��G
��8�y�Z�0�r�����N]���s58�g���w�޵7份�ӎ�~y�96�T(W����~�A}GY]�A�w�j���ԟ�)�����2��v�������B���r���*l�ŕ5�ڛĹٖ��P���9���3t8w]�l9J���Sw�
��͉���/���{3���E�iW�|�PZ��*5J��R�dy�&�eM�b(�y	���.�G{xE��[��!?��D�W�5�ll���0��S�����S7g��L�g2_�ٱ�6�Z���O��r���=V{j�,���)-�P�K��z�w�z��3l�%r;v�_��YFy��Cv�a�qrj���72v�F��w��T������C���~L���g
��B�d@*Sc`��wU��j�tBx�42���!OD�����
���BiItR��8Zd��Fo����Q1���G�-�����4�h�N�n��$����j�ئbC�� �G�`�Г ;n���������� z�V+�t���g��8U�\Ͳ�B�Y�
a�X%|��aC!ę���*G*>(NB]�pu�B�Q���@�-]u��7�xU:��n9�S�FN��n�<w �~A��?���{FA��E��v?�]
ڕ¦��0nH�+@���
��)�p���	�\��>x�an2�>��|8}Kqޔ}�&��3�������{�ҕ���T%���a=_A���U�3�� a��(�c[b�VՊU)ZQ'+a��x�����ug}b�z�++Y�I��b�ݴ�5��Pg���B�� "@T�@����Lh���W�tz>WfʝN���Q��&�)I\�̢�$Wi�����d`y �I���He�/�r�o�w�#������<G~���+Ԓ���A�+��O�!�Yg��r�|>B�-s �w��Td�浰��*�<H�,??�G~��+4�����h��˔�8�b]X�v�����:˖��<�U�������v.�H�.���!F�m�c�*��IF��`��_�4�f���_˷ }Q�w�����ɹE�ڛ23a��j���.���#��ϧ�Z5qr��~7L����}���u�P\��wҘ4���.@F��.�@�e4Y��v̺G�DP��
�cAVe_89����f�VX�"�i��D���1=�X���B�َ���p�E�������5�0�\t��8'�*g���էs� ��.!��f��U�ʭ��<;�� ?[jK��m����B�{wo����j�([��{��i�Q%TUm�S�*�QvW��	W�t��q;C�����oa��J�x\V�\1#�	πW ��`ρ�|-G��}�'���U �-�PVl? �U��{؇(��n�'�p�a��_^I]���9i�s;6$���v�SW�T��M��q+���s����f���|K{!{��v'e*�[��n+e�Kd���'㊞���R���m�ʶ�o�3J�8yֿ+d�z	�n_��u`^�Y��h��x�Xm�U,iS�ֶ�P/8�0��0�t�	��1N@�
��1�"�GnF�T,�[񙬬Ev��9�SVF�ů�/�@�ΠSW���AV��]tl�5&��t";��{�3�=܁�(�AF�d+A�|��%��ۯ��Z��9�qv%k�i 52��t���ww��Pd��T� j+˥�,�)�P1Ư��*���E0"e��#5Vl�M7ۈ
�t����?�$� �0��."�?e ��~�u��QY��k��2b:ʎW�P��w�����8�U�K�w�l�	Բt�<�f�R'�2U�t���y@��D1�(=~P��04���������r�$[PqD���!�Qn��.��v���m�������}PA;�½���V6��0��*��?�sU9[���9*��u�7��Mάen�I��snMw�ܾs��Lﲭ����̳�H#� �]�U�z�ޝ1���0!V�4�r�ӿ����Zɂ.�a�T��j����a�����s Q�+�ŀJ7<"aG2%�t*ĄYiʮxq�K�EG�������飕o�f1�b��껤#���0�)�OIZ�-�������nQg m�L��IQ�@��!�o����k���ic�+H�G3x�O�j#�$�M��j7�s�N���8�;�>n��-�3���v�f1x�v�~�"�f�=ߏ��:�1e�G�}Sm�CStT�+̠-`�/��ޗT
��_x�Ԣ����:=�d��*(��{���.��13흠ڝ�ƖT��������Bӆ)���A��y�_�K�0��Q�)<�ϞE���DpJ}���Q.�@KI�~�r%?�E]8<:���M)����B�� -.�����K,� ̴c�<<>N�NE����e���붍µ+&�@xʚ
�
�+Bˤ�����䷲���$�Xo޼m�_�A��D�r�R��6DW���-�^����h+(�n�hk7V���\�����>\�:��6�Q&�ޡ��?r����P�AmQ�>@_*[*U^񎌎2��b}�m)+J���Ҳg����0���aß��#�poH�q�&8ތLi[��a���e-��K�C!`\l_����O?}־������||�>������>��O�~��~l�|T�&K�C�N�Lz��A����ӧOR���pe�ݹ{�ݻ�ݽ{�����&-A�����&i�V�)Gq��N�X���(���ca���1�z�>l_ʞ~���U�߈G*$�*S������t2Rp�{�+�WAe�>l����N��.�+bԗ�{��8#��Iz�G.q����^��+[�e<M���n���,�6ka��W�]X�����d��q�q2O�V�U�dHȑ�@��+d�D�8޸]d@Čp[�^���T����ސ@�'�QP7�ǥA?h׉f7%�dMWR���2��U������h���|ǊC#�y�	G�� � RJL���Lc�)gu�Ą�rE6�
Zۜu�.9�� ����VX��*�F ��7J�[ژo?�7����!8��#~�Qlù�&��Zqs%nfF�ū�t	���1̠�ͼ? �!�v�-�;����r��$���v�3l���F�vy������Z�X7
�E�so�����sp��L������{�v#-���0��)?�Q�\�7i��5>wg�Y�z��4h�����C�4;����^Oc�]�*\��O=�ob���7�z���)�v�H�	�sh;�k�#���è�%$X~��ɖbnu��DM˨�	�%�HC�j~%D���@Si�2���ۑ��ళ����߶�w�mwo�Ӽˊ=a����"n�q ��[�*����a�L߇����������qcY֑��U�\!pPBi�-��2�E҆�]��:П�3��&�{8L��߫}F{���&ѯ�𷽥7�\�IQ/|pf=��y����ل^{��g��/x=�7��`�0�(�ڕ/�_�A�Ͼ+��g��+!M����1�2�	4�����u��c��p8�/FY
��2�w�W����}s��q�heai�mq^
������o���	n�s�HE�sr�h9�8��Q��P�VVn�`�n7oz]������2x�Jv1�2����l]T��GY�>\ɷ���bLd��o/xP1P���@W�6�P��'���7�o�˗/ڻ͍L�ge�2��a����(��JZ},�>$�Y*�W�Jw���U.��>
�{ԫ���q�7Sx�\��g4�_ϛY6�#��&��i�Kz�ta�٦7���3��?���������/��?o��_������?k���W������?�3�O۟��������C9r�N��U���c�(��Q�~�G�h�����O����}��t�x}����/U�>��s���e�OI���2����<(�yK�ҝeJ�Γ/�Ըd��^�V��
j�~1�O�+<�H#�L*��j����$G�W�}�/��)P�T��������R���>m;v��_!��(Z�b���˕����$>٭��mFi��o��Ҽ~���C�;�����M%jT�v�~�go� 1�L��gz1&/!���v��T��>"B!�m��ԉo�02�qЭ�?=,�@Tq>������e��B��mS���N8��u��B��E>�s�w��.���|�.�I)7c��4JG�����#��Z�����S�j!���1��
��!V>pJ�9"�2Pi�bW�n����m��-��B�Im��S�r�J��9��f�1�+@�g�g���=�r�%�a+L����
\m�<��
�ͫl��� �T�FI����;�)�i�ô���!���Q�-�u�;����2��h#��ؖX��B����.S���64�#����)�wy��=��O%�/���T��+J�6Sa�j��C�|x���è���^��]g��+\��?~���
T	;N�$~����HǺ/�-��M��e����%4�&���[������LW�\N�O���c ���W�[��5n�>��L?���פ����2������I�Lꢔ�RH�-�������^���Q�~6É������o:���0��߇���j��ض��o��q�e�T m��|�`y�V?h�Ԁ�A�/������J�~������J�'3��C��B�����1Ɵ�		Gȕ~�u/|�ޥ<�燹'�u��#̒�B�+Yn	t�²��=g�D���"�j���:�M�
ԹL�4�¶������^���w�=G��(~J"@�l'�G(e�'�KT<��gp� e������}�!P%j���]�GO����<n�n�AH_���EW���`��7�i_������S�� ҏ�����UM�{�o���n�;���ݠ�Їx!lZW��+)����Wٖ(�t�D�Rh&�9P�Ǻ�&x�|�W.W��W�-�k�ܹb����2�n�*X�\ri؛]�P�R�·�������	�����6J�'�>m�'�D��������_�������������K��O���W���F�RY��OJ�?"ϕt/��\��ٶ���>��(f��_���/��?o���G(]���_�?�s������O�/���ӟ��}������G��K�Tjݞf9�1-CA)�
�~�XeF%DMze�,	A$-�~e*l���]�>R���x�c�V��7q(Hy݉	W���V(��@�}l�d�.�x����P��o�1�)��16@9G���8N�G��Ǻ	?*���+����|�C��q�i��(�╱�W�)�G��������������fc�mmYH��*� �6����b\J��U���2Pq^�k��� �d���y���S�8���[ƵbFA���N(r0+�ٛs:[:��
�8{��=WW��oB��ۓ�ڃ��J��@�l���B�];�h��[��m��m���ݽ,k�R��&5?+\�¶���as���:8������.ʽm�%g/��r�[�e@�
�#�Y��l�v��E�u�陹 O~�y�<*J���
l'�]��r�s�1�v-[�+�%Pp@雥����_;hIȸX�(4*�G|��e�eV��L����~��f`��qK��ZeqP��e>!������to2������ؒg�I�-۾�����|�.(�yg=���u��?��$t���y�jO�66^:囟��7������o�ڙ��C�ֲ� (o��jG�K��)�\VA��� �������ܼ�6Q��2V�H��3�8�L�EQ!�RX*Ӽ�bU|�\'��\�H}�M�_@N�E0���g��2����Ҁ�IG])Jܼ� ��V�Z��(��KQx�����q��J�Y��>�yL���pU����\}�rƠe��/����B[������|�[���ʫ׮dm1`8p\�S���mA�a�'�у��'��gO��Ϟ=C[��}� ~0��eJ��ؼ��=���&��Sg"�*���ʲ~�@?�oi�Oh�:�����Pe?�ͥ���ö��m�{Վ�w`c�r��3-�.[��zmAƃ�����5��O��)Ϡ9�����-��),Uc�z�I'�U�[�6?�i����nc�q�8�îv�F�㷚1�>Ȗ�)���=�]3"����ҏ>d����0}�[�fs	�B���}��v�~����{�|Pޕɍ�%��<Q ��6c�:�mۖ��(m���é�أ4�7}\39?����� Wul��Y�����2����v���+�ٶ�����6wQp�.橣;��%��+&Ҭ;O�5s��u(j����ZnwnηG�o k o<��Ak"��x�춭W�m�[���
�*
��ʻ���e�p�޾�m�_m���������y���­��x����㶍vp��A���axwr��߇9/�Xn3�m��^����{������]���vc�>9�Ґs�)mrL��?:���m�oI�zD1�_����.���tD�gʃs�p��~l��@�!_��%��b�k5�U�N�˷��o~�M{�қ��<��:q��nbó�]�x�xS��m/��Y�����xf߈�ğ�q�f.��Kp�'W�V���Ezsm}��}�z��Y�5'�#�HZ�lǃs�ZhI��X;s�nޞo?��S�(W�~���O>i���������n绉Һ�n����Ɖ�<ߺ��퓋K�����xA}�ƽ�Xp��]Һ�V�^2����v������|پ������������c,���QV�/�O���V;<�oeeJ>��u�2e�b��!���9��P��D�En�E�UιF�9ҙ��g����3����F�[+'�SZ6��R#hܺ����9+����E'nS��U|�*e_��J�zAX	���<'{�!L>�M�Gf�S;�[m{s��}�ʝ1L����+ɦ,��-�7HS<r��b(��d�3��'���2F�{\����Z[X����niu�0��?�o�m�h�e����VƩm�i�'ã#gaS����a�_4j���	8���I Pڧ(�[1�
F.Rq����= S5�0���z&I�K��~��X0~��B��0W��Z�Q�e]L��nI���) �U� ��	�b��aF:Bt(���3�#�yW������>���)?�a<K�jR�@ZCa��>�4k���i�RP�ś�-%�[�&�nW���3a��	�<���)0]�)p&���"B'"��PeP2Z����{��z.��*~�ɘF���uw���U�k����=0ލ� Bv��FL��ߏ�%(o{���/^�����ȥ�Ǟ����TB���I���iw/����EJ9���}f�U��K���`l�)��ضc�3��Ui��:3� ���*�}@�H�?3�������Jǁ�v<�i��[��&���w�A��;������B3ң|&��4�+i�p�G�Rt�=�u߀q8H8p�3'|9����DJR�����DP�/v#����B[g��_D�u2��s�ى0�ejf3��
��)&o��8��#���1��k~&���MOf�^�N�:��t�!L�#l�d?ȹ����~j5�(,-�h��nA��Z�0G9*S�L)�}�����*�Gf�'ܧy�t�+�c��!�8�C�j�׆Ogр����4�mR��V;�4A��Q>`�cۏi�2�n��A��"�z^�s4������bGxg؝�q�X!�sX^2��w�ۿ��n��/�}���U���o�w�_�/ߴ��^o��7m��6����|���k�Oځ����9*�:/�W��@Q����PL�,���i;pUl��nEoE�m{�݋����������*���Q���m��[�����'�}8	2O���"�v��>�����?S�����kmE��+^�P�P��������M�#���{��-�ax�<I���� 휶O���R=|t����z}y���o߮�w��~�$�;��_g�O3�;���1����VI����(;�'Ϟ�g�ﴇ����;�n��7��m�r������w��{w��ڭ(N��gIo.��X��N�����-/"�{������������s^�d��_~�~����?��_�?��?j_}�E{��~�J����W�PfvQ�q���������9�C;X��@������*L7��COLT_r��m]��߸:e����@�^��mllDYz��m�
�m7�m���l������ݬ|y��-��w�5Oth,�w �%T�q�$����� '@ؿ+{�աw�N�zw����# �w��s��@8Q�z�?f���� �'�i�l���0r��n��GD��	��y/J��as�ݎ�Y�������cA��&9�S���x=b�J��(�(�NBF���p��'�0�L�ſ*���`Yi�ExO�D�I�K@E𽃈����=�A��31�&�KeXO�S�?�U�m��u��f�K��a�5��`ԟ���b��6�+;f����u��Ý�_���j�Cg>W���IsV��r��LwI��R��V�j�3J�[���(X?j[�X��:��tuM%�!��դo�~�V}��g�k��\��gEV
� ?4���Fu�=}�r�k wB`����-�J�L^M�����E����	3qkWԬn��k勾0�e*�.�p��q�LVf��jғ��4y�s�x:��}�����d-/�0.1X*8��*�g�r&�$��HϾ�L�)I�;�o�C�qƔ�5���^�XRP�=�^A��ꇏ������aJ���2�}>��`?�O�Jn�:=�ʜ���۷kpG(W	sP���Y�m_#�H�zTQ�4��S|��0W��;��=�i���nc�#�i<~����L��ְ,�I�Lj�0 ���X�u��}n��bn�s��<B�7ҍ��(YЦ4i������$��i��f�������p������t�y��+=���D���q׌ʕ�X�x�Fa��G���1�#�0#��U���gZ�����VV]����n�Ȭ����{�lx���^���DxT�\�٬}�N/�p7��7�([��h�]G��A�<v��=������(��5�G%x�|�
��V�g�n��آX�8ѳ�v�}�c��;��M$��v~�BC}кmA���C;��w�mk���Y��<��2��DQ��wQ�Y�ԇ�����
��<�K(��o�jO=EAx�V\!�~h6���[��6���:sp����\C��N�ύ�C�}I����׮ʹG��_���<���ݹ{�--^o'�������W����F;C�ۛ)?ʕyT>�IW%�eԞ�/Q���Eʰ�3m�XG.��B;�[`h0� ��a)B��,��
��"��B��5/O���)��6����гW�z�ʝkk�������v_��ΝvE��<e��=�����{i�q̱J�����u�n��w�z_�W�y�7;���1o�e��(X']��w2.��o�0mnnve����P���ׯ�+���W(`o�-⸣D�-��\�I��W�#�aj\���h�K�*�*P7?(gG��A�&w+��W�͟w���ъ��cT#Fh����B:#�E������#s�@���}6^f8�����w�4@���a
���ԋ����#�2�\~�d�E���� ;`gt`(� [E˯���Q��,s	0@a_ϔ��c��d>��2)�̤�S0����Y*��]�)���7層�r��RPaI������?��Ca/;�'�.�Sǽ���&�S&yO��i�?ӝ�F�sfn�t[�J�NY�We�26;��,�R�{0�n2�c�r��'`<qx�0L�����Ai�>�7����c��b��+%��$�O�7黕�~�̻鄇��q���F�2�+S���J_�ys�w�i8��%y�%�B�0㆟�xNŧ>�@I�hs���_/���s�Z���;�I��IeA���������j�ժ���lx��v�:V �E u����Nf�,O�9�"��U�� /_���a��gﷀ=s:d�T�F��J�1��Ӽ�M���$���v�D�	�G�B��t�>]Q��vns�&n[�ʞ?
��4�#^(�a�6u2�`�?��>�pe>~��3U]U�����<P�dl��@)/P1�솂��%w�{m�oY!Q��ѿ"FNR���#2��d�)��Lݝw����1�Hxp����SZ�vG��a�L91��%�QɲO'4��u�U�~B9S[ҡDȟ4e����/����B�+T*;����v�����ɣ��矵O>�4�gn���	?t�G~�o�m�����w���������(h�qtr���0��\��u�ޢ�8/YF���n޾����<zFne��=~�	�7��#�
<�J��%|��������0�<��}J�O}Ҟ>|���}J:O<nw�PRh�k��muke�=�w�}��?yܾ|��}��q{��~{�J��Ay��

��ʄۦP(֖���;ڧO�Ek%��>R�l1^A������9�t�mq��K�*j(��D*Z���D�u�mr^���'�۟��/�O�J��v��-��"m}� ��m�}��Qn�n��b��*s(a�н�q*P���|��t�������
��|�*��3�e�m�g���~��4�����MO�*������*��)e��2�y��@V��/')w�
�|2���o�I����i�xp�q�핎�Ҷ��[�Y�2���C�z����1v��8f\��]��~/��C)��ގR��⾵��I��i���*^���^�BQ~�^�K��&�}�sB(e%��g�.�>�x^:E/z!ڍ�0|�aJN�7#���C3&d��c��l۬����������[�����O'w���bNFn�Y AW��:w)9�)a�����~Fu�W�r�ك�.��JM�k��
!,��Si�������
�V5d�dݻw�=}�=}��ݻs�)S$��V{�R<�����{��y��;A+�B���re�ؤ�,G�C��4keD kHAC�JX�ؽl��i�`�ӟX�
Vfu� �a�~3bZ�� ���|�Gi�2�6��[p�͂��[�^0(�h�Ξ�3���x>kʿ���1�Jh�Q+z�'�Fw>��_���pO����C���{o�L��P��.�7��.;��(��I�4�"�ǆ姎gF�ڵ��vma��-���O^����Γh�W٧��P9�]�[�#9i�-�n����\����,�02�2=>Ʒ���Z"#�����/+f8�[W��6��a�z�'� ���T�����R�y�x��C��M��1��3�E��.�!�;��"gk���\���9{-_��:���:���p��
�c��>Ͼx� vF��n]pzwg;���)�K�7�Ҳxө��Y���c
?I!��[�GH %̴�U��{՗�yQ6 7�M&fd����
+��v�0�GB2ގ���9���}�������mo���1��w�x������C�ٗ�����mye-8\�S�c�s\�0U�x��O���L9?rO�ދ�������S���BK�;L������6Kzy�M?�[�*�n���B�=b�u�[]���x!��uM�qD$x
.�s�Ϻ��#����|m ��G��B�R�%t�D<3� q���L�Kl��pm��-�3����a{��߶��ϯ�~\�aa�o��\����wo`�Q����ٳ�����(I���&,�=} ~�����s��w��ju��2r�v{��a���O�����Y��/~޾��+��G�e�e�'CW�}�y�J�Ͷ����+A��?D1{�r�4�x�O�!����e�'�x.���{�IOQB���>�"��3W~��g�������[w����\�n���O��~־���ӯ�l?��O�O���=A9�����޼�߿�[��<y����1��W�e�{��J���AۥNQT�PE\U�l��4���r�3D��/�P1U�C���U��������Ϟ�o����i�W������7Q�PJ�Jl�������߶�/^g������5x��E�@��eu��AY���m7o,�G�����n���s5����/�"����m�� *K����Ev]��L�z�������vQ���ܗ����FG	K'ɑa��||����M����(�c@Ҏ�e�1�@�BzK++y��\��ToW"B�M�9��>�yW[�<]�?S���1�&#��0�2����%x��um���8V��
��v�]���`��v����{h�L��ynd;u&J�a�u�]{<�U;^���?���U����9d˹��D��� �U:Ztbam�ݧ�ݡϫ�g+���o�߹��՛���uyI�2Vu a�J���u���G�B[�(YR���4x�4��X����u�'`��g9��P�(�[��1� �td�U[�1��4�}�Q��<���E?��@�VH��!��s�o��;m�g��(Z��A:;��2�P����d�rA,
�V�`.��;�����Dq�w�l@������`@���u�΃���˾�N���B}O�6� ��E�s�'�!�<�~��?J��n�(@��n��!�\��z��{�����M#�K���O椌w����}0�<���@�7���Vx�?mOs�~!��+U
���������VY�UȲ#d4�c��\_js�k��R��Wh�nPϼ8U}�� ���1_D��ܕ�~EP �=ϵ�!e�b���x�i�_O#�I��`�|ޙf��LM��<����ʿ��5�_��{`�K��lz�ecq�Z0O>�8�C�t��g�H��\JG��?d�n�7��	�J�L�_x#��/��}��d� n����Ǐ�OT����\����Vf�6Jw`�de���T'�F]�sb��<xD:��z�]�nʲ��X�O9GQh���
�2�gm���<��z�&㢛�p������	��f�ټC�:��f�v��z��>x<<�����w�?j�������C���*������5������nH����Ol�u:�����׌�q��p0|�$�'�po��l����mm~ȫ��	�(@U|�Ǧ�h?4;�E���M�44��q�Ş7�����1���,~�D�Ӌe��8n�>;�k�[��_�}�!������?���,�x��c��' eR���6izˏ�/�l�p/JĳO������q�#yE�r�
�]䒻�/-x��Q&Y��җ_~�~�󟶟��'��3쟷�>��=x�0J���7oނo�J׭�^&㙣�����������y{�	�JГ���G(K�	s���n.�����}��O��_|���b���?o��s��g�����ͻ�U�����G�����'?%�Os���(Z_�O��t�yܿ{�=��w)��ݔѨL	�33׳���w���`�Q�oS���iZ�M��h�:��۷SE�:J{�o�{Wx�>����?���g�E[r�l1�q��G����mB�{9��֮sƉ\��r���$�m{W���-��������P8;}O?9o��nG\o���;�y�"�w@��c�dU�pl�+D� �S��#�^����Wm��f�R��D ��c��8Q&N��s����_�_���Y��#���vtEG:$2e��n]�-�x;�y)����HƗ(T��BW��焩�?e���8���G���T~f>d�1�Y�~M��������e�l�U�::��5�n�c׎�~�;��Qw>k�?���e��(
K��3�FW���ek��ƿ
sŻ�-"�ܼ��nݦƌg�G~������u� H��?����/^�E�6���Cv*L�`�!e����de%�6�,E%�0X�-b޲b<`_kE�Y�,)���ڬc�"Z�I�N��&�YMAj	%����0�G��v�J�|)Y2^�&<x�*e��K5��
A%kgW%�T�����Q:�l;B{/Oc	@�h�|�$yذ Un�A���|�P ��E���[l�f�L�\~�PpP�0�%��9�-5�'�+����*3��
�b�;+.��s�#��z73�k;�qc�<��`<w���I�C�1���J�JW)K�	T���چ�Q-Ϧ!�>�$�4HK�{��J$��<J�Q���]��H�a;�O�3\	���D��@!
���g]^[�*o��o�dݠ���g����LZR�y�HZE?y�,Yn
����ٲ����u~���o�H�����/���ۼ��7��S;r7yN.�/H�i����I���(�(w�u�f��G�Q�E��//�'�2�������:��Y)"�����V[f+/�����𨉒e���8�DX���SDVu���OO3�;P9p�R幊���|����kr�����_ԟ3��<3rVtmM����]�N���mHQ�����R�V��^W��^ �)NC�*<v�&�{Y!�:Q�p�,�w�oڛW߶���vz̀���d �����c$�(���Ö�n�vA�Zf���q�"8I�R*����t���� &e�*{x���0)۔}��i�s��[�z���:���� ��[�5[�h���ڎ>rz��ʶ77��m��YV^Vo�eB ���ȴer�?)8Υ}�?m�	���g�݌�Ӧ�ƄX;]&� 6<`�~��V&�{�c�m��˶��M���O�ϻB��N�7w����A�>�7\�m',�s'>��3�V�Z@ɚ_���A}���e���mem��ɂ�gW ��
������xО�l=}R�~+�m�7nx��M���+�,�����Eq���ժ'�>�R�����Bu��]�C~�v5J������̪�E�=���*��o�k7�Õ��'Wo�[�+in��A\����)y�����E��}��(?�c^8!_��P��;I��w���x�D�c���o�u/�@�qUKL>����CU��� F$^k(���7Ic�>���
b�,��Ǐ�?����_��iƎ�?'r�ۻw�ȴ;(*��9#�2�¾�����=K&�;e*���qF�	}[ן�y�ow�ml�|����ߵ_�����՛�J����p�:�!�s�������mm��Q���o�E�ʥ��Q�� ή���?��6a=���w/����ū�m��@h5���` /��,�M]u��[u?���ny8ϳc֕�?y��ӳ��[�"k���_��1�;�zE���+A\��$���Q ��\H���n*KN`�ݵ\8��Sw��8�8�*�n�(Y*p�JVp1w�M�O�U9&�����Y�Ū��=L�g��z��H���I��e��]���~�����5���?���x��JV_�:�XɪUR�T�P���u4R0[�(X8N*�έ0(V䕒���KI�JRr+�LNc��p;��Y��m�6��t�=zp�}�ɓ��	��6v��Ԧ��Q�@ޕ,�,�;��I�p��T��f_�����H�4Z����j��1��Y�ʲy�܇|m 
�W�^[��UW���)��@���wuU��V���_E�+a���i/љQȮ-*f�����V	��PiS�+[h��A�}��
?�5�-%�tM[?�gP���=a(&��x 3�=��<W�I�a�Dv%����rD���2ZJ�ϓ���խ�p�:G�Җ��Ce�Ҭ�Q�=�U,��+��e%�&EX�5�O�p�)2ԃ��;�O%K�;2���Q�B�Ҳ�:�Z���Tz�ˊɻ0��ބM[?��O�}���8��G̴]�kD�����5[$TX�R��$�����3 \\��� ��:�W�#D�3<>$?�?88֖���^�R�,�9�1��<�zt%���W�@ȼs�a��(L��Ԟ]�#�{��i3M�s��D�r��s!`��,�8ބ?�*�̬.�tV�b�ܭp�)i��NU��3ֹl���EB��0��0�Ơ� {v��b����/����U��
7�	��L�>�z�-,�e��v�.E� �hd�(@Ѿ|���[�!`���ģ��c��1���� cK�~���m���C��+W)Yp���X''Y���zǸ�G;\F8�1��A~g*V�")u~�{�;����/���X/��+j.(�jAn�Ռ��+x�Q�����
��].P��:�ʫ��;�m}k��d��d��(Y�/)S��9��-��[W��޿���=~���v[ZqR��c��n�T��H�J��	*[
^�
�����B��PT��귶�Bs�.J�]^1��P��d;�|	�lAo�vr�ƫ��I��,�8y�Ǜ�T��XR��N�Ƕ��:~ ���J��{��=4W��Pv��z�UN��b�\�	%��
/�r�\yG�^zNݺz���Ro�E�r%���Y��N��N� hn<ݲ�čc�+H�y���l"�l���j?���՗��kC���~]l�w���9щ�|7�R�ֶ��T�\�������s
��u��������|���:��/��"�bdxA�W��G�J1Cڊ'(jo�m�_�������ߴ��ߴ���v����B����|^��L��N�!�����qM~i9�k{�y�	P�6y��=���'��Oऌ�B%O�g`�V��:�'�ʧơn73���w|,y�W��?�����k#=�f�q�t�����;����?c���t�m���Օ,u��D���8�O��)W�<@٤t����������ϛ�[��m�nq}��!}�v[v�1�����dmA�~�A�����P������xj�]��.��Y���s���DtiɯV;���K�<$��\����U,�v�D� CS��bU�V�2#�ɳǵ]�=��*hUv�,����Q�]�����i���(Yh�S�]�r&K�DIˆ#%����!Ȭ�^D��<�x�S����)�%@%+@����`��U��<2��SJ�D!n���k*.���)�/ʚ� �坊 ��-����F�IP���XU������L�����PY�V�J�*b�3�����s�x�/�k(]�nCiK�R�\��?�gW�h��Y�eu�v���>3s�����	({=l�w��;�v�-8��u�V�X�$��wCɊr-	��
�ȉ2Pk������ĖQE �a�����'�����({��c-�W��V偻^T��e<����z��b��z���_y�2V9�>a�;��Y����PJ��U���MS9�'������'՟���:�e�.dx@�����yؙ��vA�)F���V_��<��ay�3�n�O�����>
���f��ߍr�q	���g�GW����W ��Z�c��9��ʡ�^w��������iB
 d��Wb�M����
H�R��v6�X��Wc#\��woۛW���f�Ï�_�]��3|�]����;�=p#J�+��g�Pa�Z�}�h�� )���jĹJ>e~��C���A�4��)���C0$�m�{�$�8�E�L��ZŲ��o�ǥdI�ҵ]�Y�%@�w�6][��'b�ln�u� �S�X��ҧ?�T�	���v/�U�Ye�t�/P�0�J�=���z��n#�n�i��ȏ~���G��F�	
�NVT�d].@��f��N� ��+LI3�X�ƾ��?��ʚ㭇�)�,��ʺ�l�F^��E��u���$u�Ƭ�D�W���:>�G�K�QH��d�(	�3���W���o��j2��v��ȕ���#/>��Aǅ�3�R�E�ZM0w�P�z�V��S�����&��3o�Ca��
_]�E�ŝ:9D�z����7�՛��|WȪ�N"p�C��� O��lp�?�R�I0"Y��v�o�k�?��I���O)+e�8#n���_�m�Y�ڷ[�]1[�]@��@@���ye���n�SU�t\��2���o�}�~��sܯۛ7��&J���.��A���\�z�YޅE�s�O��p{C�ۍw�o�u��_�]�{���`�([ ]�z�R�y�^����׽b�2�I��s�J!p�@k�����h[�B��Ң�Ndx92���*�
ִ���I�>k+̳CM.t������jy��s��.�;��GY�n�����W��\�R�m���{ߝ�?�f� �a>Ҹ&�?4�aR���I٨O�Y�b��VL���5�:���3�,���U�G����Fɲ>Q����dm�4�r?��\�N�2	㩕�R�l��/�0"�Ҵ�!�j�
a֔6W�F`��У�e
7�x���y�c͒�=ѭ���
���5?D�����Zm�*YԆ](�P�͖y���N��d�\M�d����|<d>t��k�#=ύ\X	�~���j��uP�@W[�uTT������U�\JW��vU��a0�R�T����@¡��O���y���h]G!B��?ʎ��G�m����~Q�H+�Ӎ���j���g�6��(M��I��]���<�E��9�qC�R�
�Lz*q��ʕ�/�Z`>��-�v�ճJ����b��Q�I�?gp�О(yY9�})Y�Q��H%�4��9dU�Ѹ3�HAV<CJ�-�����&Qʐb�7#S��{m���
Lc�&z�qC��7�n*e_��q��*@���_����>�1����
���u�y	��u�P����.{ =[�0�Gw��3��%<_0H:8:�U&�O�Zq�:s�#���#
Q��}'�\[�A'��noF�P�s��Ύ���k��Г�F�=x��U��3p���DP���Ǻ��?(����[��gU��U?�����tO��������kے�����9��7;��no_���M�S��3t�/����*�y��9u��=?��u�f�=�!�Ƒ"�*��t�R�Λأ�e&�i��a�N9�4�? C*����{FbH�Wi����&Al?g��
��h?J���ΎC��#\̍x�nW�1�m��*J(�f[*���Sm�Sȿ<����F*WiR:P��O(o�Th���gG�peq�m��y�0�V��x>��+"^w���^�=B��\Dɠ,�(Y����c�s�H�y��]�rwI>�J�=�V�&tzN�Տ��My�F�������r��O#ȗ�����+Xzݵ��}6�H�͋"v�� �b���k{��UQ�b��=#�~��+1�🀗J�Q��f�7�D�� �Ə����k�Ĩ�mn�{���z����.�s|zDwF��W2�eK�t�%c�PB^�zӾ}�FYأ<*�*�Ɵ<��S�uHs�l��+�$ø��+�����}�飶pݝ	�dM���]p��|�Qʌ�fPTI�]+�<s(Y��Oo��,4���#1^������W(�oS&�Ky����``�pk��Ǐ�2�WX:٨R;��d������_�~��7��~;�=iGȢ�A>���mn���Q��'����� _cv����W��0�B�ʰ��v�h���F�F%Zo=̇��<z0�de"��l���Yc^�����&��%L���vW_���U}�����М��|�s�2�V�,�|�r����.��-�U��O���U,y�����Q�nٲ�xv��؀1�b�Ņ�m���\Ls"��;'b�<~�o�-!_�A�d����M)Y�[������W��H�d��3κ�R`9�G�A���ْCWo�C�i��&�ӽ�
DU)
��D>΀�C4�ʖ���v��:4��3O h�c=~�H��]BEf���w��o�>���������s�vv��<2��"`�8����,Yd��k#T!)!Ė��OVC��g�!j�Q�/eC&���KV�n�J�s~%���{&��Ul�{ۄ��-jmN�������@޿��;yy���Θ�ƞ�o���n��7 �B�`v�w�(Kkmf	�b�.�3��,�;ps
n�k|�7�̈03���FG�E�j�\����[4-�'�O�$m��&�,��rcڕ��$�5�s�w�:ω�O���k�ױ��p�nk��n ���v��R�^.�G��!����e[���t�5h�3gC8�إ�*����YY�=�Ϟ��*���F����G �Tf[0q�vr��Mg����0#.�x�Nƨ�d$��M����e��1f��J�JZ:���8��,�Z>PA�6/�})3�Q�\a�?~@�DM!��c%��0�L�!`8�;�Ʉ��R0�,�o	*���,��e�X��J�z��������J�'o��Fy��U[_G�p����D�H��0|��AD0庾��5`�-Ȩ�ۦ� R%
B^)�$���������!l����{(SR�n'���Rw�ڑo� �W�?k(����`�e{���m�շ��h�]�"��J�ߑi���~�������'��N��ѓ�+x3�6�������9ك���6B?mQw]�dᩡ����4�m�! R� �i@��o"D`��-WAƒ? �V�п>8�B{�XųmU7�x��ش�?���)���B�F;=�#�9��_^nK(X
bٚ��˚�rf�3����>N��+��9��B�Ez�8��V+�i�ǸܔAޖ�Ck���� ®T�W�N�h���qk���`�U�\޶߽�?����
�N�]o���R���J�I;<���\"8�~qyB&�G�=n��[aN^��
��e��X/��Y�e/��AQ�m�"Wx6�s��r�����޵�w�m!��Н;(
��d�C/7@Y��6��zw�io77����~C�U����ZIosk'���O%��:~ �o��]�w�6�C� 
?��R@x/8ϓ~���l��;��>���A3.]Ϟ��ݬ��?_G�XG!@i���@�>wpr�v��u��/��׿qE�u����a��0����@��
��h�S:�*�|�%S�����q�!�xW!pB`Ekqq�-�_�F�2E���Q�P�^��Ψ��}���Q�5/����mU��YŒ����Eִ?2+�qyj�*j�a��O���5EZs����v��/CNv�H���C�x�:g����zWў%?t2r�ՙc�c)��行�^X����bBQ�w��k����9�d�cPpc\d��ͮz!�<8����l��~���,�$�㊳f"/c5}O�6�{�R����q���c����3Z1ny�q���c�mz�����T�J��tU.3�j��W��P�vr�	'7�Y�����΋�v�<��f��G��*���Ud�*F����%�Yۥ��m��ö��uJ�N�z����\������������?���x������0G/� A��J*�ke	-Y�K�j��d�y�����W���"dnVn	7Pqm@g���CgP���4}��J���r�oS<R�z%��͕Z�"F��i�de%�����.�ș,��q��W8�!ϯCДpX�qZ�j*]Ҕ�Ky,[w�3t�Mf�?M���B���g��v��L�ρ�O��R��LB�����)�d>��N�r��$ݓU0��%W�&��2�TԲbUg��f��aeP��թ@���+�������B���9W��;q���=an/�v����J�n���t���L��?���#m��v��l�p�e؋.JYE���*\�b���L�+���E��Cک�A����/Ɉ��`j����鏭;�U�b����~R^��yb��$�h\t��ӻ��X���A�#|�2|�;wِ:HZ�QN���Tn̙$��ζ9�ጬ
�u�l$�<�m5�{w���/�/�ʖ+/rV��������+x����)��G off��p?+X�o_�-������=9o�Rs����mN
�U�𵶄ұ᭮���
���st�,Dq�3ᢴ&�T��:���;��N=i�np�*e�ܔ1{��P��3������y�x���l��ҺC�P�94_@��A�C�~3��?�v��|�}��ޏ�C�u|�UA�:�'� �)2���=�x�����i�C�Q�2��-�bFZ�#��T��_)&�	��Y���Ezo�sw��r�0n�S���+�56�qF^V�iz��ƶd(���r�1#r����ܓ'"҄^���7B�!���_P���ٞ�w�m[[o�j$}ғ	���{�o7�sW�ی�� �+@���J����n�c��IaA�}x�J�[��8y{���n�K
6�;�vmn5���Dz�w~��lo^��lng%����Pp�����a�۸5�ի�:�3�_�h�m߽xپ����g��6Q�6�vI׳<��߈���Ώ����u�~�����6�����a�� _qKz��m�a����r��U�ö�����M)M�<�^�̩�m�Ҷ{@:����V{��|����o����w�\^o���c��l�
�3����T&ry��������ww����5��϶7���Z=WAbXȢ�[=3���;�7��4-�U�%<D�F*}
�N�R�	9dRwY��2#��k��A�N�z����������oue�)���"i���7߶_��7��5���\�o���9���I��<"#�G�Yʐ�	�euø���rs�uO ��Ord�z|��T��I2)�#�dɣ�Y�����q���i��_qd����A�g��)[i8���	��Pz�q�E���H8һ���a�_��[\
Y�W���|�-x�Ne\�`q�V[�y7���];��奕v��<{�ܻ��T�Ϲ���� J�,g�  ��D�YP0SW� 4��D�:>�J��[�h��fb�DR�05+2�,�6N�O!�ސ���0�G�w��C�֏����d���G�[7��dU����Ra�dh:�K�*Ynt��I�,W�./<�^a�H�:�.�s�*%��Y� �F��F"��O|�UC�Hv���/E*
Yl �SP��,�~v�^Q�F���g��l��R����i�e�?�C��\y�:7U
Hm�n���W�G�EI��'�=��;�i��/~�p��l�ZV�K����ԕ�(@*B���=���X�4�����(wV���uW���j�X1$l޻RX+�^��_\��v����h���"�	1Lѐ\�~5 o��I���N��/ ���?㛾��?-��]v��	Ի��I�o�p�V\=��_�FO;&�埾���}ݭr*P(Z�.j��1}��g�?n�(!�:R�:=>�����~n����_�Qˣ,��R>U���5�,߹�`y�A�w�r�Vpt���7�ڛ7/���Ag��7���Ҙ<�ۼbf������V�\�R��eI� q,�P�)9x�J�H�5m|����(��i8m*m�H�[�'
QYo��:[���SW��(���#J���{��k�K%+[~���0����>���n�0v[z�qCH�x�/E��e&t��x�t��M��/�|\�j��/c�T�U��U�=�������|qr��\Y�h�;8ǴCK��=,m'=��ۏvN��vM�:f�|b�<�3�9&֛��I'�����;mk�97B�;�Ga�\����m�#1�%c�;h��Q�v��7�Q��ѩ}J%�˷ȡ�*e���c��Q�rU�I���:�0ٖ��,�����&J�����북b��0�T�^~���|�E��B!��?������( *P�P�޼�@���(m�Q��rC�[�X'��Lc?����D�AY�@Yr[�
��'�&�o�SAR�z��w��|�Q�T�^�(�����uD>�k��~���
��\Y{��m{��u��Q��Fy� ����[��o֣�y�C��8�d�҆�쀂q[�8`��61\�x�"i!Ag\PQp%�����.<�-{�!e�흓��*����/]�Py+K�Dِq�HЀ O+j�����Q�pү�8�ǕSx��P9u!7^�o~gq��o>���]y�;<L}���߶��yNl��3�l�>7�w�(��92}mʀ�UרD��ȿ-�23c�<[>1��*��J���(X��K�����C����i�P��$�TX���i]3N���j�m�(���};�Ue����ȳ�?l}�-�Bg"aF����mk!Cr�ʃ��o��;��|&Bz^���A}O�����tc%��-,n+Y}8�,��gn�Q�R�'Y���(Y�=�iH!H�]U�e*�Պ-(�12L+��)<���*�����g��[~�����z��n���nD��⪳Z�,��=�%�����}W�P��_�Sn;�yG!�7��L/��	�U�@y�njM�0��]��U,/�H �q�x��8D���˕m;�֍
�.g��ȭ�]�ʌ��x��f�}�vc��>@�|-ϕ�յ�ٳRu!�6��'�[���LCO��Z�i��G���sY�|���R�r��P�PtbO�����զ�(FY�T��^Z1\C���+���2�R��O�܂������UF��2�!q�QI�Y��
�I?��a�7	4�M;��?�1��a��y�)ZN��O����IB�bDƨe&a�I4�)����]��Ņ/�]�IEʫ������8��6b'b�}�P�d��ȋ.�l���\d�2�*�m��<��*>ޮ��!|��c���v%�A}��1/�Cpx����wv�Y.g��;j�B�Sc�>./O�s�I9�si~�-/��N������͈&�;� #@ܿ���;vB�W�Sy2�ȃRA�U�A�p�(O*X��P#Hm"8�~�u���Avۣ�¹Ӏ:�M��O�2d=��V` ��[�y;�k�8�A��w����R��n�8�Sޏ-���>c�?,�.�qyR�r�N3�����r\��)���3-�`
�{���B�^o��V\��r�4���F�Su��J����ڲz��wCvվ�����T�?���'�a~#�Ɨ����� ���n=���ڠ���)8��:� �ͽc���c���]�r�ۯ��I�x�N]%��b�u�؝�T��/�q5��bs�[�6�(�x�\�ۻ���N�z���
��<��R���<�}R/P�@���J�Gv��H�J�[O����8:��vCߏ-o��%g��r�M~N@�t�m�*Yo޺�����������u��w�;ȅ����F{I�^��
J�g�<Kt�-����״�������u6�E59m,�6�ŝ�& |f��㧘?�#W+��e�!��IHu��n�ZB��{d���-һ��8�S�w��:��d��4�W�U��I�}�(��8���t��UW�Y~Wx�/�F����b{�L��S�So�Dց�z>xkg�}���o���Љ�UJ��ig����Bc�*K��9���yZ��Qa���!��);cjL*Z�Y,ϵ�l�*��t��8#A9�յ�_z�����c�i3�&��'�7�S/�U�z�!^�ֿ�}]��������2TOs������8]>��*~c�L?#^_Zk�+7���E��Ih�������v�6��c}�,�w_�dmnA&���Z%�
$�:�UJ��z��/�K�-��(X}��ڲàlP�B�U ;���܏����.�+�B��3
�n{���(Y��i7V����EX	˴�Y�T���f�]pk���0#W�<�a^KQ\:X`��NӠIc����È�?�(k��!U�å��ݯHu,;?q�����a��'��2ʖ��������t)ZC��������V!+Н0Q�<G�2&���*a�3G��͸���"�
Ӂw��Oe̸?�n
�&���70W�J�ܓ�s��w�[��
S�b�xU��U����gy����hf�?�?Ӝ�X��G�z�63gi^۾wf�EklɪN_�`
�Sy����r����o_�3�q�h�D\�Lּ2\��
3m��,L�q|��s����/�1��/,�T�T��Έ��>��'x)���۲j%��֕+V޺T��lͪ�Cj�qeK��J�&¢��A\���>kO�<��<]�r����7��ߴׯQ��w)���<�C<P<~T2R'��30�]��)2�J��`Eɲ��)|͉��:K\i�r���/��bol�k�sE�rY�*p���:�	^��s��c������m�Ջ�����E����Ca����֣v�E�j�<��*U�L=x�E=ﰼ���W@Tĉm����jpӟg�:��&�*��4������X��_�j�Q����܅du��?��J�-!��g��In�{��wߡp��3�xٌ��؞���e��LN�U��ItC��c��r���� M܉\��T�~x«�� U�@O/�&�����e���(Y�{[�Ó��&�s^A��
ɻ�c����w֎��apnw�r�]s���?�nm���{��JH)]�(nA��"���(6[[<{V
%DEf��A�?�
XV��J�J�+Y�0�L�u�9��X��KI�Y�����[�U���ϣ�l�����ʊ��z���^7䩄�������Э�v]�>P�p�x{*�������@�z�������|��k���3)��j���)�
i��Q�N��~��U�D�����e�����Ƭ��� ���Yzv��u{�}�����>mO�>n�+(���%�(Y(���1��_�!��簆�O�%��P��RE�W�]�����br��L��'O�g��=�[(�Z[C������ZP�cyMS�+On�v�
^z�zq�3�������]U�萑A�F8�*W�(���s۰�0ӷf�rUJ��1aB��},�x�;M�+<�^t'n���M���+�<�������iX'�K��"auG�����L��<�T����q�����-GB�/<����W�<��7�:��
��H{������V1�֥O�A�.Ĥ��3�7����1�짔$�N"o�F���s����D�
�N��<
�c�&���<O�Hð��\�� �9��U���G�Z^	���g!�B�ts->�E9"�R�Tt�R7 �������0@+��M�^�35i��;0!�X�����!`�Q�TZT8����jh�<����p������37�ek��܍�u�ׯ��î�7ꂌ�3��T�����%!
x�Ґ�5�w��݀yb�����I���g�ke��8�I��n���v;�qf����pK���v����!�������J��-d7LB'�Zv"�����7��0�������]�/1�����_�I�2�/A�YJ�xO���9��:�&�ԫ�`ݎ��d���,�Q�4���[ �����&�+2����9��MH�O�-������:uNq�g;���6w�뗯�w�~�^|�M{�������Az���x�}@n��#U�7�Qk7�K�ן2ܖ���0�����o�"����a;=@��|�6N_?��u{��;�ݤK攡[����-����_���7E��A�"[(i{����.J��������}{(x3��2��������4?06���
�c�)4)��C>G(�
����＝y���V�*��6<��4���~|{��;��^�fs{L	i3�\%�.�9�I�X2�)�讦�_�����ġ)�b��h���~���%}�p�m�{�B�m���J���כH���^]�����l'��q�B��B�gZ2a 1+\�����sX���|)�ʍ�j��tt�A�2�7�y�+��]���NO��?��8��-�~�ju�F[Y^k^�Q7#����佀P��D:I��nپia��-��˫IG��ǅ�M+ϖy���BQ#�#_9�}i[���wʺh��7Z�::�&�0���:������y��=؏�*pz�Ջ���������V�<���PTpҼT�>.<���}�=�mbXe\@q~ia�={����g?�G��(��[�i̸��(�x8Qg��G�4�S�H/�P����&@Xi�=t~��Թ�����x�G.*�\�#�&}�
|떿\��8�jm�#��퐝�;2����X��})@�x����H�%�#>vMlYNね兦�7�0���/��L��:�O7�}J����|�����&��N#L��p@��L�@����/c?�v&�s��e6}�����F~�L�C�F��+Jd�t�hٸ�[;<����8\��+�u��"�Z'��W֨0뢐��*�w1y_�e�����F���&+�yx��˽@C��\FE����Ue'7��<�cDJ�z��Os�%��'��%���Cf	�T�
1��?�*(�����B����̂@���P�sV�b$$`<[
E'W�b���m�ݗ�W�r�n7i�o+��Mo=DS��)P7^���;�t@+�z�{��dpȅ Q�p; 9�x��g*̏������qs���9�6=W��z�⨂؟UU��JU)��w�歍����V��}r��U�)�
݇)e�,�z��^���tژNC�������rt�ܿˌp��v���6�˕n3�����G�i�c��݄!S�0�g�J&�#N�3)�ߔ�I�!#�` )>P�[�
1a�0t�Y� ���yx�JR���	�`�1�����|�po�+q҃g���k~h�K��f�������֡��a?�v=��U�~�d������w�����io_�l��hG{���a�☄~b,��}�������6�Wތ�5�A�?�]#޼���KZ�G�mo��ͷ(v�&�_�W�~�6߽h��9���s
���!$[W�պ�g���+e��H��~ciP�9><h�{;��`)�����@QPn���(��O;�o��W��Oh����Z���K}��i+GA%�-�^o������pw��p���f;����R��� ��W�����kg���4�
�gK�wչ@z�n�55ʈ���T�X�mށ��WKǏ|f���ԭ�o���h������~�O:�9�������qث���LA���	��Cв�x���Z��b��,���G^����!o�S��;?��vp���=��`��������g�!��T�9�P�#��TL�����(;�ܪK$�/ޥ[%�|�ϬB��s��Ga9����{���\�藧����Y�����?�H�I��=���S�\���'�f��ϲ�R|M��A,C)P��	��P{��|�='�?xDIųPԋ�?9e���I7֖��?k����Ǐ��E�"mu������v�9?9LzN��J[�	y���:/V������<�_�k�	
�*~��{'��GwN��¶�#���P��1o/���-�ŭ,��[7��7��H�7��(��\�� M����J�J���4(�*��^���1Ѯ�¥q�r'��uH�c|+9U���(g�q#���!�+f��+c�,���O���c��1t謄��)��z��g��֌?��Z�G�M�b:vI3���S����B�4��5�^i]<�K��C΁�Ӟ�����uK��#�$���W v��������&��ƻJC������%��@A�.�N��Yb1��S�Fc����R(<`&~8�r���$����0�g/�UV�6G+�g:N���Hj*Ib���t�3��3t��Х]CS������O�	�[;`́�B�P�0�+�d��ɿߍ0 �R����
a���ݞ��L��p�o��=�Ę@�;ǔ§����]a��+�ʢ���{�j�b)qW��*i��_ޭ�iĿ���(��F�Ӗ��|�FښzU�Mƴ>J��gl mL�z푖�E�~z�I>WL��¬�e��&�j��1^�5f\���55h�����9�!��_x�C���M*\*X�g��_��(�A*p��j߅:OT�U��7�*^���f��K�;�(:�?W��f̠9u��0lo���o��/���iϿ����׿B�Bp�|�����m4$F)2����s(`s*U��(X���q������O�N����V;|���{�M{�ͯ��oۋ�~�^����{���n���C���]��()�՞~^�������I#�M]�:q���b[E�RX�½ݝ�����2�ǔ����mmEt�0�SF>�y��W����1Ew0t>�qe�ϖ�?+�z�.�M`+����'�#���+	��������_}��m��~��ݜ��M��6�Z��6���z)J�Zl�v���Y�J�4k
�nA�o;[o�:��������a'�\�fQ���5��Ь�Ź��sC^��N��Htr���*,=#0C�WJ���jL�o6��턯�����6A	��	g����c�G��9޺
�G��Z�.Eu�D+��Px��m�7�|W
#�+����Y�.P	�2���B����iWN
*������!ЫЧ��s��z �((��u1K��R?�������;�#�����v���F�J*�RR���PO
�Ե��(+�r[���ԯxͣ]��2O��\Yl�?h_|��ݽ�
��MC�������v ��"{	?��fm����8~*_*pk++��ڍ��"�%+��~����[_��������%M�5O�,P���eQ�#	��e�2�ۭ����;�7��,˸A�Е<���2y�����`22�d5�um��c��1,�FΖ7K�%�U��iw��w�l[?�9�'�w|�xL������?2>w�J���}�����6�
����B�L�
Saÿ�M��K?��M�I4��7��yZv�Pm=�5b���	m��6W�h3�G�:��-4�D��ax;I���ׄ�x�Q�� Ai�K���E�^c��E���tCZ�ZYG�p$qՒ�(��ҹqWX���ѻ�,I�#3B$�@R4c��i���qJ!�Q���k�g����ui;��0���_��j�	2�%��jl��P�yC�W3�5�Ս1�b�e���W��|Z�HM�T�욎A*��� ĉ��0eO���t��}0߄�g�m<�5�p�0�����c*�~(m�\�^qS-ڄu����<ήe;`V�%R�r��J_
V�QM�����Գn��t�6�G�Ƅ�S�`�{�9_&�	h�Ug�0	3Ic����t?�Grw��J��=ekE�˓���Ϙ!�"�� �<�x&;Pe�(m��)n�x�'c�ʳD�}�Mf
�I�Z�v&��Wb�4�`	Y�c��/g1�M��]�i���޼~ٞ�������������|�^�h�����;�Y<��Е�
t+�)4��3���k�(j�o_�7�}ݾ��_����_����P��"�nm�A��ng(X����2��,Av�@��,����M��UI���V/D�rˠ(��,J����7��cUpO' �Jw�:���ȫSL��w���q�t�� �2��W�㪿�s���U��w��!߷�d��vs�ö�;����n�0o�{���0x�vwݦ�K"�*��*P(�W��*hJe*J���#l�����v���!���+�7�_���/P�_gU����uoF�r��LV�,P)Y^��K���aU�ꛣ~2�a"O@�$BH��
��o8����VVpP�Ԓ�JEMa����#����۷o�v�W�}��*B�2�b[]vbe�K~,�}���2�V�/�A���h��)����q�*J�+���6?һ����޹�ܿ�n� ��s��Z�)����e�-��k<����n�m��e���;z�/W�Pȩ�Ў���X]m�o�@P/�`���lGQ�w��+wȥd�"�Y�t ���r�Je�|Qb!�K��3(4��o�ݹ���F
�V�l+��ɑ+p;9k�6D�����(s��e�YQ)AZ��~�CI2Jd��'g��h��[]Zh���8��67q��$�tݺ��<O{/��n�ĝ�eU".,7�'O�1��'(|c��	 DBp���䣦��_���������򈐱:�=�?����m��X��.���y���te�|~e*o��Mj:�a�>��������?	\%8�%Y��i}����+G��Ȓ���p=�����ք�Pzm;�x�n�Q����i|���\�4A�&�7��WHu?��V��%-���H�����r�M��?t ��ƣ�I�B��)[������(b�UA"֛����f��5@����:����m�����r���TN��0(\e��?<�-&D�m���'P
�pO��3�1$r���,��v�C��C�d���5�ix�Gs�{;H�U��γ�I�'~�\�>��4��$���ɐbS}Y�EM�_	��v�2��y.��%�����?>g Զ@�>+ӱ��mc�)L,�;��3mc)ˮ��I��w�+���������y,>�^[StW�W8]%_>���PO݌��3�&�b��T���cd�V�h[�T��_)��W:��C�"���<C%�6N򅎅b�����y��Rm�]=�l|��5<ٺ����o9R��7�K��*Yĳ��x��r������}���/�m�w�����տ��گ��/�7����Ei���p����a�nG��8����My�b���oڷ���������-i������޾���&�������Jԇ+
���3| l�m�.e(
-��_Uo��L֗t��B�\�pz��&W�W(��9
���yt:�~��Y�� ~I<Ϙ^���[��z�`&t�{�t�����}T��)���
Q�N�2�v�]���uF�V?m{<C�����F���wvN�ہ"lmD�Z�"g	w�GW��V��Α��GI��Ӿ(�N'�n3�q ��e�,P�?=+k������YI�E�::��j�[�eiּTTǸ�n�S����	�G}��If_���a����r>7ϡh�Ť���*ߐWX񾓷8!�r��̣Ǐ�'�}Ҟ}��=y��=y�=��i��S�>�����0׎�ȶ7��DyBA@��V4��[7WQ������[����*�*�>�˂��mP�uk�=}�����/��y?����^C���y������<��Z�ϭ"��X]nwn�l�n���q!�>ޫ���UVT&n�ӧO�W_~ޞQ�U������!M�!u�MJ�N�V�ma�p�cxF:�6��QHTXB��S?�k-�.�)t����-ӆ���'����*U�i�ڦ�d�+�\#�q1D>�CZ%� H��t����U-(/arK�+q���Ey�<�xH~n�t��l^\��t�KK~}�2_Cw��2����1�)o8ƨX�`Yw��(w�)G�U��Pò[�p�D3�}�gӊ�60���Ҷ_Qt�5	���3���iL���m�#�~5W,+��)���g<�#3�:�S �r\��jb��i#��'L�<�˫!���y�u�.W���R��r�c��l:>�������~��՛�|����P��B)@6F�8�C!҉��Ƹ��f<k@�_!d@v|����n�aW�Pk;<����ܨ�L�`� ��|T�<<��#"�X��l�>~��ˬ����#�[PF�� ��r�71��斷�1�l�og^(AH���s5�=��@��L@f`Yk��a*r�?����,�럖$ZO=zk�6ސ}>v�t��vf�{�@��9�ξ�C��3� b`ۉ�� ��P[EE����t\@��Y�f���$P�
���۟��в�����<�J^��oA`�@[�ި�ː'.B��ZyƳ>z�T]QOV�6�*�F׼��?8��*�4��a��=� yAiZ���K¼G(��?��%8D�5{� .�A}�@��tF��
Z�6����j����g}Y�(��;N���椓4��X�Β�W)9Ph���Y#����؞��A0F�h}SW�X����$����>�$eK5�ee��b���C|����2')�����=B��1wٮ1h�!�\3�;� N�� ��Q���� ��<��ϒO9��@�:���PJ�ipX[[mk7V��{�͛7ڲxy=��ֻ�n�-|�]���� p�~��� FڮZ�:5 ���50�K9@[a�q��Ү3 ���������`o!XnF�{Fޢ�r���p���N\U��h;��^�U��mw�-J�˶� ���_�_�����o�w���(V�$���n{qB��7e��g�o ]�hZ��q��~i;���+��}2M�K�FD��v��6/wG0K��9
����K��| ��M=ԡ�m�/d�a�'}*�?����cS��z�����1�64m;�3���7�%z��^G�0Ǹ1��:tbm֭{3'����V��|}��� �lѝS��%mǴ��������u��c�[�<�s��p~�M�n�\Y���4X/ƀ�}�5ݎ�m�8�2F�͒׌�y9K#44�2x�{m{ە��-4����[϶A�D�i+�3�
ڎY�;}R��Gg��w���ˍ�v|�F�e��vz���T}k�Z]N�*�j��#/�;Y*Q*�k7����n��O��$�����,r�\�{o�=@!z��a�L��g����(Z��d}���9���_>k�}��4����o�P|Tzn�X�^i���l��i�~N��?#������O+��k�oyu�ݻ���;wWx7����q�߃�Y��O>o?��<��="<q���i���g_�����O�~�?|��߾O9����]Ҫk�>�K��Y�qE������ڟ��'��~�����,�S��pw��%l�Fnmsץ2�I/YEY���?���������~���ϵ���J����N�)�+ˬ.Ϣ��k?����W_<"g�9h�1�|�~�������D�<�]~������VV��5����|J�\�v��(�@��"���� �������n��lwn�ὗ����L;<n��˝���<o���E{�z:���,���P2� ��:^�q��"/;h��:=>;	��9z�P�v>Q:�G���bo�m����9�6�~l�n'ڮɃT8�DJ��Z9E9��@9E���M>;=HH�
�(��� c2OdL?�	Cc��ñ�6�O��Y�/_2�a|O��6j�#&��ؕ� �f@�4c� �:�C�7�Q�(��%˄M�&�������ʝ��v�^n�);4y�f{��Q{����NM����(Y0�u��Cg���l���H�h��,���z�3dC#���2>Ҵ�s��3B�G�00��Nf,ng)*n�\^��/.p��fJ���	�y2�,���2J�3A����K��\�q���溵}���ǈ��)�����9�u`)�3�\�-�pm�`�_�[Ϥ�!{�Qķ�?�|;��o�E�Ō�:I�Ǽz?m:>v���;F	H���CA��$0�;�Eۆ��H	�7&��Ch)S�����R����]%v���$������%V�p=�$��D�<-C�l�B�cz�I��R�-�nv�j����� � D<��R���	�Nˆ#V�t�I���������{��;*x�m�(��S���_�K(Y�t�������U��S�`�3���z7ꤼz��z:�tz��P���B�-cҮ1�+�+w����whF�!d�?�R�>�ٙCB�̾������ʔ�V}5�\ɪ+����5�2[ppݙH�V�`$V��m���2h�q�=@	���j[�(@�����@�]��,�o(Ȃ*n�ǻ��؋��P<X��5�ʩ
��W��zz��>���]j��=��6Q�T��!֍7(�Uy�޼z�޼|�P����}�3	*��0���ÞM+>+�/x9�3�U�����ĆV3a�pU>J[Y=������2�7s0�z����*�9��Ϝ�H��Rvi��!Y�I�n���#f��|�I���d��~d�,�=)S��NdWCuG��+G�8�QW��4hLe�å�b�m�}�67޶���\p`��D���6���S+pd�������;�줤�5
�[��(�ߩl����5�-�s�T�#§�W=+s�U�;��~��e{�z�6T�A�oz�-��
?X�O��JA��}`��݃�����~��f�?��Ys���1߉����?�"(<_�
���L��S��B�Wt�m_�����W_}՞={��q�=���vV��I>A�2�g�|EJ%�U��?�4��?��}����<Ϗ=D0����b�i��?��O����)
����uk-[�n�v���y}��v�=zp[��	���x�D}A���)��ۧ^1����'�|ھ ��>�O)��Ǐ�ي���Jգ���'�P!<��� o!��E1|��I�ɗ_�_����?�)
�ì�ȃ�����N��2����T��8�e�B���}?�*JF]���0���3�����~��Oڗ_<�F�1=hso���x�ٿ������`�xN��l*Z3�P�>@������/�����GWV�aʱ(�)�����7]yBA�?;��잷7ow�7(W�=���6��;��Ud(ަ��al˝sX�e�A<�����my쬝'+�A��Y������l��/���>��Og���3��4Mـ�CC�[
M��I$�a��*�Q���`>�?��X#�ob/�?�w�u��G��w����!��I�pI���b��L*X���(o�e��%�+dM�����r�-�T9�rB��/x��c����{wn3�S���������%J��7�4~)Y�F<��2V*Q�I�*L.�f�\���gK�y�𷠵G_�X����"D|���ט��<��f�l�qe�ٶ��`���$��d2O����r���qQ�;͓�,�ە9�n=>�@���6����Y>V��d���WJ���['����L>YXb;���-<�{�,_�/�������F�R�� ,G�� �t��(4�nD�g�(M_���%ֵ�Q���6�m��e�`=�W���-S��8U����od��`�ָyk�Zi��S���u���Ĵ) �/|_�&��G��T���h#����_/Q 8v�ʾ�Y(l*�*;��~y6~�����a�����Qu��7I�h̭k�nb��֏)Y�x������)��:��R&�I���Ԉ����L��|�vϧ�J��qL��UYlH�>�L|��:�,��>@\7o�Ҡ����On�"��S�]�ʭ?��̴u�Kٰ�^�����7���WP��ge�L���P?,��,����d�U��4W���} g�� '��˳�J�Y6����YuE���;�:����ì"l����}�{;9��!�=��]����y�>�*�;3�}V�S��19�9�͂���l&/(�e�]�Y�ԳJU�p˖ ܡ?h~�1@���sճu�ӎB51��;y��̓��_������/�L���_�<�����ʌhS�suȉ��\�M�Ϊx�R��u���߹�tw�����.�[9��L�їz�V��c���PGڣp�Y~o����L!O��N�F0���v~z�.:���#����la<����(W�6� �`}%k��[�<��>�.Z��x���'(D�=��K�r���|��0οz�׶v���3���}:u��<ܱ�>B��P�n�WVQ �D����$�����|�m|����
҃��ڃ{w�I�]�?L�J�}�ݒ�K��C�G�p���F(�u�f�C8����h=y�$ʔ����mmu�ݼ���̟��}�9�����O�O��b��t\�������Vp�{��<h�<Ȋ�-��;�����h8��j��$̭[�6��%�3��j�'�=CI{���w�o���w(��!�<@k���V��ܒ��Y���	�zx�L�Cg�� ��⣒}�����OPt��&j�m����_����۫���}��:'#mCH�F<�C�[�.�O�����<�GHi]�TV�6�����~�n�<s�A�:y�ۈҼ�Jnm�@����o^��������붾����|������0'��6A&�XUu<P�sBDy<��.?��>��Rj��/Zo��c����\9�I��×E��;�:vy�	CV�du���o��|�3�)���3�pLE�r��.qM��#�c��3y_aR&뎺��`�]P&w'��h�I}��R�n�v�kT%�I	�����"s[j���P�^�dm2hA��Gik�gl��dA6�GJV�A*�8*3d�p�~���(��(F=!�nY��Cf�F+Ć5�D�[�,3��l��r�"�ER�RpQV����T���ʔ�@�(Yﶏ����{ҕ,��%+�F�fOf:B��}к}��H>6j	`�ﳅú�y��h]-�8WDĭ��$��}��WI�>ejí�#!�M�Tgx6��d8���fT �ZP�N�L�m��uR���V��.������o��>I1��`r(iA�$�y��I�"֖6d,���*���R�^J\՝��8(���;Ä��.m����=��>r$�*g«dQ���i�P%�=mm;�B"�0���;��Rg����d�ˉ�h>�ی[eű�N�I��Wă���W���e��w�&_
���Mn��%�,��x���CN��-�QJN����_�@З�]�d���H����9P�~�tueƹ�-�ޞg1M�w܇��`�щ>/��^�28R��0d�����Ҟ�XByJ��O��?!>�i�O4߁�}*+E��s���CQ����+�Ͻ�^�dP�/���U֟ʢuXJP�8���a�<L͜{U�O_�䇡Qz.�����0'(}Oc����j�����+�t�5	a�Vޡ[L�3|�qä����_��/�����I�t��u�g�����M  %K^l�Jsn�����ν�q��mof���(�����M��^�^�C�\e�vbT}�����&+ˊ%�\Mjx�J�
JJ�с�u��?���ͳW�oo�m[�������������*�����(]no��L++^|�� � ����Ѿ�OR�������7��K����SW�T��܅Cx���'���o�-,���u��};������|������O�/����'���ɧ��c��;��Eouy~19�K-��\���FM{��ʪM̵�e��ʵ��{y��=�-�x�?��qeg�s��a>��{Pwnߌ��%��#���(sQ|P�T�n� �F�_�����8�I�H9����[dZ��	��^�`�rs(n�Vٻ���������v%Э�˫R�������mnmJ��R!�o��`�mP�5��v['�l���ZIE�gu���u/���*���g�X�|ʝ痳�u��͛����z{�v���N�S��O�xVIZ7���\;A������%n�9��A	q�SK�@������2�0�dy�JjǏ7���P��}վ��e{����V�=]~I���
�*�]\��m��fy��s\��� �M>�y; װ,59W���G�ǭ��*Ya�v�p�}��/�1M�J�w��	��qbm(Y"����G�yc�X�a�4c"g�󴷦��;�ǎ���0�p�D1��/�e�J�;��j<S��0��wr�>�B�T�ZZ���&���Z����?W�h=����J�:���ma�WJ����:��3Xc��Y�:�e8�W%�!�O��iӃH�0O��x�ʀ�d���O!A�'�s�`�� ��+Yj�����-9WJy[}�K�I�zt�>�\�R��ݻR�ꃽ5�d99��*T�����Үx a:��?�#d�8����0�3�X���=�ԯ^�]��A���t��)g��'�^�.�UB�5f's����J�/
��{�Qq��PW���?p��%��u����j^�]���@%2��$p�
?�*xvH=��c��i��UQR������Nޏ��Tg@��+�n���vw�,���'����.���/^��Tl3�JCa:�O�# ������{i:�*/?6?�5�&��g�Q=���`�c�_����8cSV葇��fm���H)X���;��A/?�/uBU�Ϸi2��7iN2��6�S����D�PW{I�>�6��Un!�<P��we�F�LS����m{{�t�C���7ᗴa�f^���/�W�(Y�k�+��J�UB����0�r�־|�kj%�"�k�O�?��Y�u��ɸ�!S��1���VQ���3s�c�Mю�Q8�̤i��<X�
<�m5��ڶ&q�������Tcm����I7~��A	Vi M�Q�_���^��z3y�_��\�q��}`m]�r俯G;�����gQ�h�I2%�8�?�H�ms�UW@�;��h#g��d��lC�E_SХ�2�i�Uo��ue~Ӿҩ�G^�֣|��	T���<���w�d^���-���9\o[�޴�܄��m�`m���h���Ǹ}D���nŉT�_��Ms.D{�w���+�*��yr1�6w�������K���Ej����8���@3\,��A#�4,�,�x�Fr1t�9�N��J�u&�����3��tcf�`�?#?�����=$z�^{�C�����z�]^:ձ�i�iZ(�SS��PWqʨ8iO���k���^ad}�~������rI��(��Η�*�] ߃vL���l��w��iD��,�^���e�r��g�e�E�+����q�M.w2����Z֧)P���:�6q=XY�a�O����xj4E�B̓�j�a���є���g��8?���@JN
���Ӷ���޾{���Y��ݸo�W��������(�܀���`ǒ�1
xw���gSa�Ζ�tP���͓���F�����#�ӰI> "��p��0�Ω�lُ�$m�,�rԔ��������5�/�]�.5���.�������wԶ6������{�h?�0�FV�Q:�";�3�b�j��:Rv�v��eh���wA�����˽>�N�%���Ҙo�Y��ozҬu.�� B��a��6��QtJ|�p0��kJ���� @򿯜��^��0�ݹ�[�v�u��2[�����5|�+�A���|��*�����g������4٦����2�?�1���l�V_XZ�oc�T#� }�E����7r
�������UL��M�_�$5���ځ�^��`�ܘ�� APqZ�*��8�� �H��B�}G��{���� ��B��0C!�J߹��?���\��8Q�Ew��ɿz�'��;�f������\������	F�(FMH�Z��]��Rb�^������=�td�6��o=��aKc}u�n.��)S;4�V�v��t�:s�)���]��f���4�=��s�9�q>B�#��L Vu�� �q�0��q1��Qw1f46bw(�{������ѫ�w���5�KQz(1��z�UGJ�T�$��:��	ׇ'Lw��.��?����Bk����J��z��ݷ|���%t��^>�����	'���TK��L���ko��w�u||y�����s�UՈJx�Pk,�|��J�T��N�0��DER��668G�3������[�I#S����F�F�`ɢf���E�W7NaƓN�4�h���m�U����i��EK�|��H����O�5*u���JF�ʁ�� �+�l4_� �Jf�*c�R����~�E �
�
xf-�'wYs�O�5g6��B�z�}���h���mEٵh�u�{�\9��z��%�������:�G��k�\_���h����ٽ���QgZ��v��٭!N�e,IgЅ��Fu�(�F�z�V�� �x�Q����YɣtON�Bgx�n%w�V��U�_D���H�cDm�o{\��?�Ý�v������pgG�W�s�� �C��Smrj��?�A�t����W��
���{��_�'Wm��*��*�vͻ~z�^z��K[��1ޗ���3gg82��t��(R�<��-����E���l�)��V6��(��K���w}�1��Pyu�lP&ax � >=q��v�W��#�����D�CF�`X�Vg���F���9t�ī�#;"g�@�ӱl!%�·ֽk&=�B�����c�k���H�;�kڙ����^���"��ȩ������~�À>:rj*���'�I�M�3��}����
a��g�I9n�c7{�Έ���}^������7o����߷�O���#����t����|F�m��i�<�dM�Y�Ѡ�~<L6�2 L<��G�}aaw��Q�Ao乆���$ƘF���(i!�/Ѣ0�\'��t�����U{`�Xv7�� Ӷ��owGt��|�Y1ډe{�(�+�3�Lx���8�;h��{�V�ma���	����UG�N�\I��<iFw1�
J�A�ƺ�z�v�{��K�^W����*�r�2���� ��a*�z����e��'K�<�:vJI@�8�\r�F�)�[7�:�fΑ߉���N�Ј4q	�jg�p��N���>����c�H0�X��@E�%HL�)�UF@����VeŦ�����޹���U	B#�����|�g6�mŢ��Єu���fϬ����x�cU��*�Qg�zU��;��@<�i;�g���&�hG���v0�a9��;��NJE��;T�����w�����?[��������{���iZ*󊲈��S��>ކ�<�u���Vy{<s�B(�֍4H��H��O��9�����:<�iOx>힏�ug ]�u������sY�g:�ex�^K�Uù|�I�<*)�X�P���
OqRǙ�F9�g�{�����_���
���Y�̧� �����`?�"_|�$�X���o�5��ٰ<�e�|*�ذ��rCs�>�G�����/o�}�	�3��:0��ɻ�P�u_�E����J����|��{�G|�����9�l����1��}(#Xv
dd��{�G��l��Oc�����#�^_��29z*�:XŇ�V��"=v8y� �/<�8����=z��A��9<8h��h?��)�ÃCxh�ce~<��FP։sJ�[�]�c���g�hyNNF����'� �v�Tv�9��$����ä���*�P�Q&X΢O�V�3��5�j�;��s�<�|I�i���a�x����K��4��oG���I<�p
FѸ�QƷ��3���Oœ�)0s�ydD�g���Ǚ=����/������]��C-����/�[���P�u+o����F�F�
����~�v�ؑD�?uOD��T�_�
>�Ϣ��R\j��$�����#�!;�-S�]w���<ϕ�A� r�L$r��7��4Wd@��M�5֥��v�-y���>�/w�C���Fwo;���x���i;�(���1�z���K`��'?M74��t';�!�;�Ɲ�����x�dw7����G����s���n���]{�槶�Qk��mq6@ %7�Ѐ:�Pd�����Cɏۧ������������>��mm�=
��{��Da'�wxx�s��vض0�6>m���o?�בK#�671n�WvB)#����3�S�=>��?�:��t��H: ������͛�o�p2�yu�RM�{;�M����Pp����-F�.F3�jc�D�Ps�3q�d�"��Y�+�2b�{!��ec��rO���/�<�Y��/7$Y}�@]����v�Ά���&����Ae-%�yx#�to0��>�$|O�鼕ߠSeWߩV�P�2��'��W�Q�>��tK�WU
$���O�:�D� '�9��f����f$�-�:˨!��ĳm���)�k
�A�����g��-�p+���v���ueC����s���^2�E^���`�]/���;|=��3�\;�(���ߥS����{��R/{�J�����H��ŷ����I^Qa4�Q:���]\isK�1�΢g�67�s���1=
a¶�������nu����U{&�)�8��=$�r��;0��u
�Ø�T�*�a,�E����1�K(C�?�U�$Da��U��S�2�B�����O�eA��BX�	�@_Q�9U�^�C;��uE91��.���(�ɫ�bWl���d-\ޘV�#0���UV*M�7A.#K����t����OoP��=�H�0P�%(	|`\�m�m��5�����kz�m� �L�˔?��y� �'��^]��b�������'����^��p~��"^����t��*�4z�,�s���|-����m��ct)�$��J�72%�'�Y7�-�.�_��/L����J�C��� �)'H���-��͜�/n��Ƣ�5����BV�2�=�g߅1W#�<S<��V�Bx�P	�ũ���@D��m��w���~���u�輪�� ���w���r�ן�뢧����2ʪ���y/xșr ����t@�A�s�`��y��t�s'=UC��03��t�O�)�<�.m��uN7m|b"���>{�����2U��ӧM�7(Co�&�'�4��p;o���ӴL_�����R�N� �#5�)��d�rk��LK��e����\ْ�����ʗ�"�^�ԛ���?iM9�#��A{�U��4�#����|�̇���i��]3ܚv��]BUF��x�5c(������i��K&\�/q$�g����W�=���=ԃ��˷���7<|�y'�5ڲ������)k�<H�6˝z�1��q���=�8Ne�|Rf�3Eb�[�|�}�/���o95����]C>W'JW��?'�i���+r�5|�N ���#u�>2�p9OQp!�ލ�[��{7>Xߺho>�{���2N�s,���Ki�J0,��q#k�Q�3�l�m��͚��Zw�{��-fѐ�)020xv7wۛB.����ɬ;���qup�y_��Fב#E�m}}k����������0��n�����E���G�fv�q唷�O;��ϻ���{��i�`�aX�{�>S�޾��c&ܶ\Տ���C�4p���^o�yX3e&�B��`G��~��c��k����0�t���C҆��G�,V���E�Rob|�WF�BZ�-#Ԉ��� ��1hs�Ra5�#r��ͺ�&'xGg.�O�c�����Z���'�ᣥL]԰�\�n�:x�����T���C�ʢ�C�R䥥�^���,�p�K��[�K�Y�kYx�Σs�m��0��#'����_ka���|�^8�K��u&�>��Qw����9#�k�A��k<B�ѱy�����V��������1��eO���b(#|*�X�au%Gʥ��5��"Ϗ�U:ǧ`�o���4�����"��?��8w�����Dv��$�T>
�eK���x�#����mj~�M�η��Q�z.�r7��w��&Yʌ�,�/��S[�C��;G�r7>�7H� �5.2�/'�]�	� @�U��0��GrU�����X��P��x��h���T� �U+n�y5h�1�:��Y5��,��{FVA��,�F�N��Y����&��:uʋ`TV-+Cf|)���:GNTVKUb0�\�.L�@]�{���g�����	V��F�J^͍w
���T�x 	V5�NF����=���R�����&�s���cm��G�C���2�4�4�0�h�5��1�r�Bg<)��� C�f�z�Ψr�֛�n$�e�j��+��4�:V4��N�Z�^������;�G��*,�{k�P�-���U*�=c��{M�7���m�`$f�qyM��%,�
̝���`��t F �?=u«�C�$��;|x_���ʣ�.�]�Sa������H�O�3c�Y�)�W�g��G��9���^3�U�hV�,���ƙ�� 9�8���r�=
&��˭̹��B7y���@�:���s3������ׯ0��fa������c���(2��j�9z#�uU��Ai8��?�ql�Ijdʬl��YnQ��<�(�4�1$;8�OЪF����Jy����}T麫�w)'�M`��҆��хA�G���Gx���%y�L�˿�w������LZ�c_��T�(�}z��l����}8Ն�ń;�2}�h��;N�3_.��|����B�	��\��C���e�|���	�rJZ�����n��n�������I{wY��e�PP��+#�{�'}�m����uｗ��g�V��	X��\c*����Jg�Xʫ��6F�J�8m�8a�69#k�C�Р�.�+8�{c\�<3"�]�,���] �1F�����#ksC��i<�(�nѭ�Q8�.��a��idM�Qv�S����(�	�H[^Fyz�֞>]n���{k��?��mC�?x ������Ƅ#%�0�is��8�&�`��M7Ex����G�>b$m��6c`mo�~?kz���:�ȕF�O?��(�;�cl�庱�a�i��S�Ar�;��#�TN#������-g0�ݝݬ�������Ț鯓V�5��ã#��h�Ȧ���P���ɢ׬��OƑ;G�45�ΐ�J�Z�"�[��r��<�8�A��Qwփ�7S;S�I;==���oڷ�>o���8�B�Y��5Y��?x��vF�3�,��M�	�U����,G��Aԏ�%�J9H�~���`�Q��i\gm�����*q��SH|��j����fUg����ŕt]cgG@�U�y؞e=l�~�0r�	��	x*2�|�8鄄o�0N�<�1�^>��gv�(���3:IEZ&�N`6=`����1Ȓw����w%������$[i�� ���}���?��0ʩ��W�EZU��٫�j����2G�(gg<R픣�C㓄k�`�z�5Y�����m�q��ȿ��������(c�:���,#K��&?p��.�.hC�N[�(��W�Q�TdG9�H��qG�l�{!ja�,+U��s>�r���h��g�����F��]�v`(g幃K?��tAG����H���BH#KA�p |od�<��Pa
� g�+q��	@��}��s���C�u;�����۸�x���?`��bH��{����U5bUu���*nY�.�����n��P��eJ�#WeP��n�,G�4��j�^�e��ǰ�팥L	��r*�`TJ�@�5��=��]�|�,��� ��EGD\A`piK��сb�^�q�B���
�.����0uil�z�rUY�����
�q��5͔�Y��$�7/�gl�M�??�e��zj9C4u-��s
�g�)����ۺ�}�͗?��[p���+��b�}��w5�U��@ɢ��&��D�P�»�"����1���u}�!�8P#�z�xۆe1�Jz6P�Q���^/��%�n���I<;������?{��i?zܖ�g������7�Pb>E�s)���V;i�$�e6P*���W�dū��=\����M������)���L��)v�:{"�`�_4]�� XԦ<�(d��~:����ŵe��S�$C��H��)�ː+�,^����+)������
K6F ��W;���g�QT����l���^~I)���B�hK�xseW��Xχj�{��\b��\��_�^}G_���Z�7�۽x����5��YG�����⼎��U�]�+ҵ|�v�n��,u)���?�F�Ϋ�Z�����΋L[��"��ʥޓW�K������b��	�r G���Lo)#�LC�3��)��(������	�\���u�q��S݆�����ؿ�8ή���yy�:+��3t�R�h��x�xl|l�&\Y��:��ĸ���<����1G��O�1��*��~���o?|�=��^F��¬b�����xG��c��ۜ��5o�%o1�4���0�0����G�������������>ai\��r�F��E[Jw�Ȥ���~?�R��u���61��?��o����۷����g���{G�0�Lw�2����r��hx������`�AvB����%��]d����S�NN�-G�5�]��SN�g���3g��H��Wֽ�1��LeU�['g���%�.�_�����[��Gmqi&m�[�������S0�L]�C����)`�J��85�B�үtꨫJ����|�h2ȵ{�����P������W�|�\��Zɑ�t:ȏ�eҴ�UlQ!�vq:/����-�3R( W��2�J?�S P�<w�:��%��T�+�M�{,�/�������i���w���P��]A���rur<zU�랹M;����O.���i�A�������U/�̫��9+���{�5������0`�^�^�^����@�B�!n�u��l����rTԎϩ{���r���C��m�����Y0�s����D17��n��tPB@�4���t���==?CYw��n�?�!2͈B:���F\���ɂD�FB���/�7�I�!�#S��9�8�!x�+�)��HX�Km���� ��P�� ���P�ٿl{GWm#�茆�@C�r��j(�+�	���kXv��w�c�s�E�z��ĳʭLC�շ6#�D�l��h�u��`^�) �Ƿ�3�+(�� �9FIs{�!����!\�W��k}U���Hb����K.�4�0�4�N��Q���l�]���vu�M��|���m,�`�@@'m�FJ�����S��Q��~�S�����X�o��L�k�9M1an�TC��v�bxD�� ���ǘא����І��x�Yq(e�!��\���4Z ^�VW��oy��tL*�V#S���F����I����ОV��\ˠ�VaH��t�P6�ݹbt�Qq�>�JR�B
�Ѝ�a<h1dE����Ȗ���@�`p��Jۯ}�ɍp����w�~�]�-�]���������:� �5�M�⅔���9�6��
1���7=Q����@I�p@^DIt+�K��|lĸj`]�3J�ZS�̖G-�F�{�i���Lg���/��>i�8负s��-�O��Uyq㌡q��ʚ���o��.�.�`o]�Iكc�f�4e�;O�iG�4x(�Se�C;r�&Q6�ɰ���V����+dhC:�����1��ihTFo�Y��r���#�qw��ʽ�P�C�d�"v;�0t\�o��zCyI��L��IE_�M �G��]�t��0�k�%�o�Lդm�.����+|BJV�ԗ� �o���
���Q�4�Xr��"�M�w�������x'_)Á?��O�;׻������uW����핋�[w߻j����i$OeU�Ǥ_�Zg���!h���F�r��E~#�ON����Ƕ��E{�g�6r��0p YBW���+q)�O�Z����PY�m� [[~/c+g ��[���2��g��h�|z��ֈ��{�i�F�з�h��1���SxU/Oem�#����ݙ�ClG&y�L&/��G�A�k�#�����������]t��v|8�Ngh�&�ՙ*Ҥm&�C9<[��
���晩^xG�l3=`vaz�=\�oϟ��'W�5�����~�������z�en:p���wD������o���ƒ#S~��O�b�xr~_�7�=����4��S<�roDa8y��9xu�ᤦ�i��D%�^�!�{��EwvaD}X_'�Om}�)�o�G��m} �=Oԇ�40��9�����	�aFȤ!����kt�Wmqq�K�h`��~/�V͵kȤt?uEDm�v=rK#�m�o�74��#�٩ɶ07ۦ��8�G�DGy�|�����_����U{�2���Mڸ��m��7����}����޿���o���	h��4��?���I��Nq��Yn�,C�P�.��9k�D:=g�9f�\CЊ��0��ܫ׸��hy]�:M�fhc�W ۷�-wf�\yh��필M�'�gr0�,ظ��k� |�L�WV�v8&G0z��6���в��'�{�0�`���/�_���~���6�c�g+�y���p��#ˇ5���щ|"��T��v�Ns)Ŗ�:`ȓ_dZ(Q�T�)�}�կ9�M�#b��e���X��W����Y�^�'I�
�X����'�	 �D�q��"���X�˨���x/2<���(uw3:��4?����ǅ��:��ٓ�`y�_�'S��Jfb.��܌���	��"+��k���[QX{��x�~���$�X���� �y;5`zz6g�LC�1������:s�u/��_:7���Q�Q૨|�����h���.��}��}�׽�ԃ�A��?�cRR�$B�beS���U�v�NzELt���/>���WWV{����`�|�����6�����B�^��
/�ܨ�n4C� Ì�s�D>��0��a�^eC�b@ѐe4�2|�����v9��*^8�vv�y	ׄ��0���HL�S��2E<�� ����u}����_��9�p��V�`%R���E�P�{w���zJ ������	W�*è�����{�.y��?s�k~���s������Ƌ�<��{��Z��쮜��9s�U�C�ڧ�^3��@�XD���Pמ7t
~:]d�
AzU�'���3+�>pf����>E9��M��sF�OZi4�����yNX�����T9��Gw�H�������+/�3�'��x�2�^X3�!��q�U�иCp:��"��,���}���`�!��T�ܜ �I�A8��r�2e��,�|}r~�k��#{�m�������Ƿ�����a�Cz�%O�+9Ű()�Kg�t0@5��=��:����M������=站�{���S.���Xx"���
j��~b�`��}h��%r3�Fvh4�p��ý��pw�B}v���X/Zs]��������R9��R���=i���lO�ݞ���=�m{��[�m��}���h�����(|���3�9��6�������/۫/W�tT�^
�_�+����A�)%�/�^��+�?�1��\��q�Ai�U�2�������#��6����u�
'��Qc I�4�)̟D���:H�|(,u�xWsJl�Ά��ӹs�F�k6�?�g
���!�r��y+Ǝ#A��?%�leN�,�4|�L��D��mU�qų߲;�����A������U�r;4�ww
�cc������C�h�u�i�wp��������^��D�T�I~��1pS0�'e��z�����~Ѡ�T��~�,���Ô�	ߔ���53�.8�+P7�v��Ӱ�Ѧ�
�M;b�_�sw��S/��κ:s�$8w䦇I�M�|!1��o��ʮ}vT!�r^#��٫r�fU�w�?6q���6l
���
ݦ��_S�D�LG�x��ep�NYD��m�Oy-���h�y�B��	��,�]"S;,��X��c�7�&������)�HE����<�a�-�<h�����յ6���5��C�����Vo�	����D��|��@��$�]����;ǃ��e�>�x�*޻{7��q!mi�b������3��<���=��k\��v����.}�G]�g����$R�Y�$i���QWE����"*�QJ� ��PT1��/�#D�.����Ȳ�Uh�H�빔�Q?33�u:�Y���@=�tև��L�:�󾴄����K���J����>��oƹ�\n�9�q�+��&��D��� D����w�������рı���O�	'B��-쉻�?���O������t�[۩�l���O�M�k4�|�x(87�0�{އ���x[��,�0�`���p?�f�"��E���;f�V���D�UB��kt�s�A������1��8����|�]b ����J�\�|sn����'��4 ��Έ�`FE:�RV��7u�=O)K�l��/���\_�\��1�:W����1i�pPX��������.�]�Iu�s������D���o�����}��]�q��Pw��S�R^��ܫ9��>�N������PY�W����H�xjaG�-�:"_��*Ҽ�=ST`�!�m��dc��o���n�%�1
��#o��Ļ�"q,����`F�C[Ri"{�,#u�<R�<�V���ė��>-��F^M!w]��ۊ�����LCe�Gj�0�}5@K�+Һ����'�m�J�U����*wÀ���)��H�s���w�u���h?�%���)F����v���u����q{��S١B���
l�����|�������:�Y�|���p�H�>S�``��I�W�微_�JC�QqV��S?��	�3��%oL/�^���!�>>�k�;��>�pwy~֮ϑ�Wԣ����i�3Kmvq�-��D�=m�P��jO0���������_�՞<���w�g�l�|�V�^���g��M`p�a�����f$J�S�s�S�]($�>e:����>�����n�T܆Ε	�{��C��OǊ���^��[^�z�S������I?u���A[�O����Oi!F�4!� �N�+c�~���)őG��ȰW�3s��!kf(�
��C]��c]�O�w7�5�u=�12�.���V�4�5)��CȚ�<���gD٠�XvdO?�w��!G|�u�$��'���W�	{@�t���<�0���9��3G���fi�͟
�2��7���);��Y*�҉�(K�e�ޣ�a����gӀ�~e��d����N^j`�rTĊ��A�hȦk��Z���Q��)H�!�zՑ*�����Uޜ�;P��L�~���3!�'B�R#J#���l�l#4d�Y��5k��Z������N;���]K�vL����FYf(�s�a�a������A�Ț��;��FV��8�)3��Z
������<�:s�|Vm��<���
D���gG̖���ö��I[\}Ԧ斨i���z����m�|APa����ˇ�뒍]�Ȉ�{�
n� O-ܻ��!���G|_`���k^��q��O6Ɋ�-1���[�nhb���ϓ��B�]�g�X��P�մk��!���|�*�@�B:��/��� *�"��{N��-��ڽ5m�Yz�!�	{��]���IyWʹ��y�
2+��Z�ϝy
�Ť�u�o
܂1��?y������x��g�֊�\A��S~��u��
���0	�k�K^6���t�=0�K��'tnd��!����ʋV��`��iXiHma�|jW\/�1��X7W�ꐶ��~O���63y��gF���d桯=�kkk�.������å���� ��Y&n\=�@�dN�ϼd���Sz� U�igN�e��Q�E���]{�օ��^�4^�Q�sw��{��ݹ[n���
,����<���UF߬,kSaWBH'�{C:S;CQ��� ׄ�8���W]U6%����V��o:�wt6�O�|6x�S�t�����z?�.�𩒖�vAC�=�UB�p�]]"��#��t(�̠�c,�G8�UP�w��m�&h�7���k��M!��B�����;�����g�
J{�/��T)0����_|<H�rPG*
Z��W��ƛ���FQ<� ���G��ϯQn�PnP®�Q�U�J�iAz�?�s���!~6����rh�2���Ȗ�A�g$��L���;Ԕd�Ty%m�<��Ƹ"=�'�x����]�@�m�k}���w�f���|ҎPtN2�	�G\
1��[���t=�鑆§���]�����n�m�;����<�N'�o��/4檂lT�Ls���ȱ���m�M%!��^�_���?�y�]C�m�2���(O͖�M9lKx�W.B���{;�\��V����܎�#]k�Q�8�������m�ɫ���+�_�����Z�a|�\����_z�p�b���=���{��件��+�.�,=�x[DQ��Q���h;�R��;}UcĶ�*���RH�����{Gv��ԫ*���L����8غ�^/��S������9*ݝ�B���Q[�őeh�ؤ)d�!^��l�Q����׳�{)O���HGY0����Oe�&Ay`|!/#��P^eMvMT���3ƚ��ָ&���%q1���4��wڒ��ز3F��Ú���LC�g�ݺE�J)�U&�R	�N����q�Ɨ��������R��ز�W%�)������#=3�aC`��7���S�"׶�o[Yפucd��n1H��)�
C�qE=kl�T�2�)/�t��Jħ��S1�E�e6i˯�Qx��G�S���Þ͙��>�髱TS�<*�J�:s��2¬��^�Vdt�f\�8��IÑ�~We����F]f��e<�E�a����ǰy%���kћ%�nXi��efm���hp+�&g�,����#ףs��>��*�ړ�fn��.��/��گ���PE}O��Um}:^���'���˰�,�I�¤�n�t�{o����۽dgˇ��_������tk�05�t{;1���v^�w�G���L:I�������#�z�L���$ q���'���	�eDR�����#���"D��YV�i�*Z��e�뿄��"�C;ݳ^�E^C`_8���OAa��8��"�}o`��
���A��YWq�'�P _����$���<^<��W���$W0��cx�D��[y0��	�	����׍vv���S�����.r�(�'F��������x�+�����GK���E�n:�Ҟ<Ym��>X[j��smv~ztA(�z��E�MC��"��5�e�}��W��4����@Cp��blݜQ�2��<9F��WRF��ޑ��2�0̲	�lԹ��5�qd�%k�~Z���Bx��rU�X�6���+��[_
U�۸��F*]C/����n���g�_�6���f�G�����`
��1.�|�3,Jњ����6\�����r8a��ݟs�G���K9�ǔ%O���m�
.��P	����ϰW4�����M�g�(B|d�?X�\�V�Q<� �-��@�v�߼j6Z�VN��S
$S�e�"Z]濓^M��`J^𩽔���ҁ������]d����=�XC�4S�j*�F_�)�J9�O#�� �x2d�
��S���(6�R�͆Ru�^��8��'��P84�n
�G�,aV������J^��y>�Y;rގy>�l�NsRw�.k*$8�����M�u����v0�>���m��ah��}28Eީ�y@�FC,R	���GS)�V����[/P�;�'~qF�Q�o���n�������I�\TKu��I	Z�c�wڤJ�rH�L;;�o�����Ƈ���ᾛ���(â��L��������=\{���T=~�-F�Wm��3*�ٕ6>��B5߆���(�K��62��&�����S�W\�`d}���U{��oڳW�jIki�)ry?.�)
;0hdit8R\��jd��>_RF;4�U�U�ѓ�3���ăjh
(7�]������)�G�m���mû���$�ܨ�i��4�z"o��W*��@��

w�(�zp�����x�8�hdͻ�eq!�f�3e�^jS6�m6C������Lo��S��~MX���G}3���4����0��	_:T���)����]y�wzeOw�s?Z���\W鲎�����rz^F��'��c���L�T
t�y�=��M#�uoN9�-T1=�\sݞr��|8r�g��!�7#���
�e�<e�� p�Z�߄32�4,�xT?v�C-]7�:�����ҡem><�̘z��c�$v ���3�w��r'g�$�fC#HL����c�t,��z<��}F�xg�;z�٭YYH\0��Nkt���8k �����������������w;O�uS0��c�mfn~^����=3�d����dH�h���]tx
Zm_�L=�7�� �Fʗ�w��O�LIl?+�2��ߵg}�~0|����}&�;D���ǐt8/#�Q�ȱ�q�>9b���oF�1�&���d;G��ٮEΈ�Zo�	v�@��������m��~����;�D.A dm���,��S���ƞ�a*L$��k�?q����ʴH��O=(�BĊ@�4�T��[k��<e�=���n��������Z[Y�oS(�[@�	M���ɣ3��_���۶�{��r�y�x!�<�[�Pc�^�J��?I!.7�[}^�W�'���V���1�/4H�P�*�V~���M�|�4iDs5���2k5�N���:��Z�dë1┺2@2u�� [�j�L���ٚ
8?W��g��g(�{��^ů,-��%��.�E�>7�p�x�x����mȲ �:��!�A�k�TiJ_Lc��NS�`%dn��
S�Mz���f�.���et{������
.����{ϋ��>�Tр!t�Տ+nZz��8�05ƭ��#�����+(6䖳�ߏ~���-C��g<�M�W|yM�A�J�n�����Z�>��k��W�Q��1_�"y�����`��F�����W&���S��`�?�_����_#;�
�:
��@+:����  ��IDATS�Zm ̺���T��+�����r19vrz�vv<�b'۷EI�!M��-Z��Sn�P"���g�dh&���F<�����Ep��e��� &)���8�4W�+,���y>T\k�+��0���5�`�PJH?�0k=��|����mrf���/���D�\Zm���(�Km�)ES��aVyu�%
d�˘"-!���2Q��E���W�ݶ�59����\���n��'ɏ�I \)/Ň���^#�"<s�4��ӟu]~�&]�S��O��ϝy��^a�_���507��At���Q�6y�R�L?��¸z��?�k��������N���+N�Z�^V�\_�=x��/?��V�'���OY�N;�ڢL��S'�ц��sUq a���(���4�d�
���h� �@mu�G����%�������tY7?�S���4�GuƏ���һi�<�������Ë۶��>l�O;���d��E@����PE\*��~%jjf^�̴��$_ؙ�X;��Q$vH,,�e��W_=mk�C%��C��-�7?m� �cG�נ"|�H�e�9��������(�F#�nP��|����O�R0�Ћ8-�����RRV;M3.��i��/aL'���	�Ž�3���d��:�z���Q;Ez��3V�����,�@�Qd���8���?������C;:<#G�	rɱ9���Г.j�pˑNYG�albQ6
�(����N��Ϧ(����O�s�@���H4������X����v|r+�JG.]�"�Y�顼��K���qd=P�f #@ܿ�S9Ҥ���AךκQƌk���
��.1�OC͍i� �n��mN�SWٹ�r;{'��A�;�v�N���c(B�F>�p��]y���xq@]�.���$uW����f��;}������gm�vN��}���=ێ2���8����ЊtX�C�e�¶��Cۼ�^��M7���5��i��4|o��c���p|���|_i���B�$3��]���ׄܤd�£{*��i�c�V��"ؐ�7�Ge�l�����LY5��t�G�nx�ϟ=y�^<}�Vё���uNF�G���M�,��Y�Xu&��<-P��=V�
I ����P��mYK����* ?��h�"�,�zc+в��ϡ�^A+�y�c��[P��@O��5��Q�I
�.��`8�ՉF��U;<�n[�'m��)-���� {�,iH�p���"��@����ʪSJ�}�<���������E%���e8�k4�w �bc/̹����N�L#K��u��Vn�^gR�[�u��GW�Ç.�^�N3VW0���F�~q~�-���s��y~n6�����dj�1S?��C+C��7B��Ec\�{�sʃ�I�Sj��z��[��+y@��D�d�A^
,�G?w���kx��et���ԣ��������妯4���ŉ����_�U��>'2��w�y�%����Jv�']�,������y��ԓX�;_�qޗ:w���[�S��.4wy��{��/��u��x�2ܔ+ȏk��2L��LA<1�&2Æ���6P����
�������*<ߺ���6�҃ƃ;jdI'E셾0�W	�g������/fK��I�?�� у��,�0OG����#m��֯>�l�,q�a �Tt��C�c�[��6��7�7&Ai�_�������q�Qۀ�o�r�֍23�q����e�eh�1
ޢ�Z?�!/�A���b[XBƢ����=y��=ut�U{��%J糶��1����6���&��k�k�*��X�,���S���'�� ��~@�2ʦ�F]F1�o'��읬)�¬�h����)������q0��CQ�g�߅���>���~��7ė������r�V���7��1z�r?Bݏ�m��^���㇟�۷?���_g�����(GƟ�n>~Ҟ<{ɵ6���_n�s��9k�+T��W��ί��rr�P't!%�A�W֣��
#��@9�8=�r#�V{�-� �ã\)]6�_�_���/E�y�y x�2�:�M���f��_�������A�=T!�D1�pw<��Uu8d����Na��M'����c�zf&�SHҕ��(ԓ9����'��+��J)t讦��f���������u����4�\��J�,T���4n�.��� �#��Xw V��Qh�3E^Iv�EY�Ϳ
��C��z�<y S��4�s�a�3��]�x'�X_���,��8�R؁�=��驎�(~T���gr��ʊ����#ȱ��h�6����B����CW(���/� k,��Ny���8Eѩ��Q�g�x~Fxp,�*����E�euu]p	Y�h0S�+����m���rD�n0���Y�i�|:����)`?��6Vn���T���ѓ����i`z.�#���J]�*��e���i��#�J����*�8���ﺫ�6ɽ��S����պЦ�A͂�P�1t�ٶ�si���S�.H8g
I���%x���4&<v<A������˗9�@P���r��gn�p����jS�AXl��J��Jt?�J���R��/ᡩt,`��x�Gкv��y�%-�x-��D��y��g|��۴i+H�3K8�~�3���it:ޝv�d�B?w�k��3�x�+G�ҳ�:���b{��vɣ�<t90�����эdyN։�!���+l,�F�#K6�
!{��#��l���N�x{u3UL����XZ*榕8"��>N?tyi���S�#��=O=���H[ń� �acc���u��u�a���s����='��֖5�F���@�U8懰"��k*��dW��T���;�8uwgd�3�t` �`���ŰJ�
P��CطY���z�����Q��r�������ֵJ$X�2,�g����e>���� ��� Yj�0tXmqQ��E�U��+���i/�]h�!V`K�c�L:�njT��*c+[��@�x�����Ʒ�C��TT�3{i�:����4�NǠ>y_FY5�}�2��ʯ7�¨��/�.D���	�V���1�1�M9�C��g��K}�g�SOC������q��;��s]�����;��mbv�{����ƫ��?���uo{ �\��Q�i�La(�_�&�x��*6����)ȭr�uR�q�F�FV��>;e辌,m���H��u��~=�.�I$��4b}q;I�477��i�fh��3��[���zP�n���L�F��rˆ%�(��4gMy�X�GYBx�;eVx��a�Q��ec�[�����}�Wг�Tނ�R�Iy�����J�@�@ ��퀀g��wtDjfv�-,"[Wa\=�!���i[B>,�=�ѵ���������r����ն����Pd�PP�\'��_}��N	~��$
O꓊�O��l�`�=����2ڛ]�!_Y�.i�]>��:����7��;�H|���x��?�����%��p�J1%(�XP�C�rTم�>��l�6�b`�n��ߴ��u�C�c#�"8?�=�M��}��Y�Ob$��OCS%_�yfkh`I8ΤP��@�� ��T`�{ ;>w��U9�Ȥ���U����k�`�Q�}�0p
�2��o3�si���$0FA�.�3HZ��w��W�K}�6���90�ߴO{�b���#t���vq��U�:���(����'y����M��kG�4.�v�N e��W_=k/^=��Zojd��������[�dk�,2I|�dZ�BN��,Ӽ���T���n��s�i�RD��M4�j�Ӿ����1���vz�
��.Y\��dN<����Ǥ�)g�V��z���-�@�Z�a`����39�v��bp�D��=8<ho޼k����9�8��-��+������G\�lt��F�0��I z�F�#։����1�O +��F�O&1"���"�顗�@��=q{�ϟ��V�c��ѯ�.��i;|�	�I����@y��+�����J{��Q{��I{��Y{��i{�TGZY^F�-d�y�--�/�D�	�^��1y=\�?�HG>�Ki��:%l�8�g�4�#{�pS���V{H��ϟ;2XC�vʙD��t�ό7������U��9$W������֫�����]��x������vv7h���]U>[G�Ŕ�x�SS�K�S.��.[��Ç���U��>2F�}��v��Ix��k�Q���T3��o�=��*�=�:�\��\t�� k��T��7�V��x�wBǍ���*�իb�yu`����1�V4��F���Zw$k��mtA`�@����22eo�J0���rL��)a��2Z�p�C%X��VA�����=x.��KВ_�)�1���g,[����՜X-�����(:
�y�`+�y��uY���,�0�"c�_�O���D�����W�B�յ��,�KQ�&�z�P��`/o%����U0سR��zExR�k__��=�Y��q��~�*�Sn�T�6
Z��Pv�YYumՓ���s�S�£��-����sn��CÇ�y?����lzf�	�u]y�W��=�S�=�!p{,d��r_���k/C�ڀ�#[�;�0����� �k��!F��XO�(�Wa��f��/e`uP�.�F^�s1�\�KOzBt��W�T���p�c{gZ��k�F5y��p)Cn��Ty��:W�\�a��\�+�\���W����}ڽ�i���޿v��eޙZ)c�0�9�.��O��NJ��id���l�_��,���x �=i�1Gٹ�1�,�#��v
HFD��d#<�����4�/*�=<��y����Rz-��@���N$�?8LxaFӍō=zZ1v�H��cE�fn@�M2��(��Sq��Tɒ���0��P*�M�CӔӺ�=�9�D~�!��]Y�)����mN�6�.w�����PZlKN5[u��Ӛn��������,J��"�jfv�M��#0��S�v� 0�V�˫i+kx�
�u��=~@|;���3�G���̺�w�3�j�'�p:���RYe��WѴG?��.�.��������=�B�]�Z����p�c���`��t=_�^u����	�Q�mC��b�� �/���1��g�n����>b\mm~h�]N�k'�M����x��:s���6�q��PT,�!t@��: [�rq��� ��2��X%E���*~�M���a�)~�LCN[�ˈ+펝z��<�,��]���ʚ���n (�k�"5�2v*���uE��P�w�����Q{�qH�~��.��m�
�m���&iDq�1gG���؁#M�~H"^����O�D?�����#xcĈ��j���mow�����붻s���ARt�6~-�v�u�vʹ���P὆)e��]�]؎١
�O��!��&6�3��+}��=���9��:1�u��D�#�G��H��S���I���I�פahdC��ț�����C`��v�QqN���e���]y��m�h@�͈*E"����&:�G����knC�ݎ1N��]{��D�p�x�7h$��oc,�����hZðq$��Ed��y<��ɓ�	������W/ڷ�~ݾ������W*�ۓ��1Z�0�0�0^VW�����(Fܣ�5�<i�^��n��@�^}M�W�_C�N<�[B�2ߗ/��W�G?k|�?z�>�q��i{��%��+��؟�\�̹-��(�@z��I�õ��>J9)����V_�K��Wћgl׬o���|��� g�����vx��6Q�)k��a�Xq���Ȓ��ue7(C�yy�$��]�F��y���mK��7r���B�g+3���g�;�K�$e��&�f�|r��K���VeA�8=�k�`l!�3�:2:u�K��|����.���cL?�nV��-�ہ���?�&k#K���	A#��h�:�� ��HL����%�%��A,o>=�\S����4�D�ʊ�`fRH��4���#�i)KQ��cd9�bW{j-��o*B;I�ڰ���<��:<�j�����3������O�f)l���)��l���8��ji��<�s
º���:+Q��5�w��+��T\C�3��=�4b�)u�m����L�YXn~q�θB�*hI��b]�k/�=<�_�x0��-K�+�u���ϳ�L{�g���uSm id{��x*@c��:-�CO��k�+�S88�@��A����f�tyg#.���F�ђ�T@e(�Do�Ks�Q|��e��u2��[W��=�hJ����e��b��ç��Wh�(�(���I�K/�'x��"���᥷�Z���r��A_����ƒ�_r5�4i���Ժ�W�	��R�M�V�w�b,&�{��.~���4���S�Pq�y��3<JY���F�^��R����krV�V}��òw8F�tOeX�v�&�j��V�F_ڶS��S>�?{{{m��S�����~ʮ���eqz��l�"-CsW�4
��n��g/(-"����Q��Y�Ebwf$+�YDT�uj�����t���e�!P��؄L�G�Vv:�etO��%1��Vr>�C��G�Q�מa\�H���r��Š��Q�>�-�3��]�&�	ӄ�К�qZ�SW����ť�99�&�2}�J���˻~�^5�4���P~>��5����+)�e�fT`��i��Ev�S��-^5�Ow����/�g�⺋�[�n٥���[��͏8Gx�n��a�(ʡ���n��Y���mkk�}x�����{��-J����9O��@:}���ڣ'�2z��b��3%������FFޣ�(��\;��O~+%Eee��8��>=`��<]�Yk�U�0NwN�>��LS#L(_�v�rG�1��X=�&�<��ώ�9:���z,�`�W6w�ۇ̓Z{���(��(���϶G�[����ݚ\�Mgr�m��q�%-�G޼jK�Q��z��6�<a��ҋv�Զ>m����}�S;:pƈ�O���[�4�[q�4<��rQ����X�~�N�kme�������D�C4��P��O�i5]�g89ʓ�g��O<�{��}�wM:vlY��H�Jժ��;�����V�g��菛V�Fi~�@�����q{�a��~��}��&o׮����I���d,�Ҵ54��[�k<�BSD�$�m�(ޑ6wϼu���Q����1d�k���A�&�r�iu��+>j�}�uF���<Őr������"
���/^<��5J��k�|�����7_Q�/�G�5��DZ��z�����`e)ZfXa��O�|�K�����i:���o���0�|�|��q�^�����0�^��fzK.��,G�����<�dy��E{�������O(����Hۑؕ�8;�f���?�*yK�sŜfXg�}����μ�+ea�<!��"��+����H�bG7�u��f��LT��ٹ�s�+g�����\�����'��ߔQ�5H���d�ѳ'ӠG�y��L,�-gU]����h���8��5 P����=#�5��a�w����u������f[��������n6vVG���s s��h#�4V�d5���OzJi��a�~WP{If��sf�a���$IDD�;dOZiD�07��]_Ὅ��U�A���EX ]����)��E{��6D�D��C��m�xxr֎�C�r�� :2�$rG
�$Oo��rW`K�]#/R_���I�i���9e��Ynx�z�H�wo2I������	�8J��~�@4�Q��r�=�_�g�v7����,�F��i�k˙!t��ϟ?��h]^Z��մ[�"��s�K165���S���E�N�X�s{اP
�܉���e�M)@�Ӡ����v{���:E�%m�4�n�W
Q`�t�ZƤNm|�mv�ъ�p��*�D���"B?^���5t�B��b	.Ŀ����m���1��y�H����~�(��f���^F����d^�I
Q�z���I�"Q��H�7�����5ګdwμU� /M:Q�wR��b8���BP����Q�x&ρx	%�}��^���+���e5�_<���DP� �\��y��Ƃ�S)�H4�P7Llʪb�s{�t��p�$w�rn}��.�A��L84���ng�rJ�Ux+��Z��]XX�����gg�����?��?�!��%GRT�M?J4�[�4.��0Q�/{l�v��W�CO��951zӍZ��(M�i�I��	��Tk�N������zG���FA�q�8��TA���+i��f�l�ק��iG��B!_}�����>�?ǿD�xƷ�661O�x7�p͌�#�V��V�Ӑy�@���D��~�Ϸ(X�T55��Kȑɰ��F�#�O��"u	�R��:#�a��]#[N�[������Q>w=Cv��%r�QPZ��%�@5>��1�^����#�0������=ϻAаMg����_�o�I%�ɍ8��Гpr��������?4�GN]��˓�v���~z�>}|�6޿n�����BoЩS�GQ&/�N7Ȕ�/���/���jƀ����fN��x��$3=u�O��^��ܱ<|�W�y_x�0T�ҫK<x0�;�6�lF�M@A�������J����^)�HUFڜ@�%�%�m�.����3h������H��CfSmw���y���}8l;{���l��]@=c��P�CG}o�/�pV���t=�Ѱ;�i�9���a��̡�ԧ��v2#OQП,���)`�i�G�mgk��y�S������C�u��8m�S����F��P�m���&�En�1�����gm��"�)ΑQp(���a��0&n��mf�����n�S���ap<y��f&Q-P��q��3�.y�����e�r��Vat]����t8�ܙA�wJ�$8��F1�'�~b0����\������i[�����D�5t�R�̶��o2Z����s���c����.�	������J�㌂�����#���O�o6|�N�wzz�w�-�O�"O���N�b`�PN���H�Y�h�+������F���S���v�4��|�ǉ��f'�q�来�T�!���������Hsn��Y��MN��~`�1�u6׭�_���V0��3�lya�-�εga�-���3�h�f�c4���*�����Gȁ[ŀ[�?^s��j�Mk����',OA�f@D=^}��4g�}|��mm����-�3:楝��$Y��>�K�(	����Ta�U��6�AR�t�~���/��)f�g7"���w2�NF:w9�N%��"��]�W�╹��`WM�y�6#|tB5����V��M�uxh��<�6�T���mS��[<��������g��"|p�K��m�_��YA��n��;��@!P2rD4^
�ڕʑ,���qQ��=�QlKɳ���ȴ6@�2��n��P��vz����tROU�R@0��f���i��Z�>���H!^�"i�H$�.F�Y�X�י����u��'�1�bP֊�
�"$"�������+��\�۹�c�п���µ���VE�2J(��^�8�����&���CW*�n�.�PR��n��7{�:��Ӽ���:�w�^z{:4Z��š�Y!�H��La�#!�LT$V	���B$ڸ�-��0��|�Γ�8�[�@:[�°���L1z4Re"{3�k<�����S��)Ј�u#�c�iEC|���T>P�S֤-W�%Wua��W�x��/~�R_��6�y�犓�Й�UO���s�i�c�Sw1�����ݝ.��T"D�$~纴/ȨKB���/���C�җŻ�������>��R�[�5�E��NKٱ1��
�J"i'.b.�����w�i������Qe��[`�T�ǭ�2=e�S���\�і?�x0��ڏ?���;����)�6=����ujo~�,~��]�1�X ʟ
F�V��q�
O�Y5��3��I�{�Kp�@fT��<l0lJa��N��%-�������/�&O��^y�֞��?{�=��Z~@�Э���ZhY<���Z�YB��[�fݒ��>��}�W'8��k]�W�Hd�<oV�T��}}9%C#�u�d(�Νάs�YC��&�y��W�(�����j^>��kp��;���$�J���|��5yw��A��/��y�fƻ[�%F���n;��l���Ƈ7�YX[*�n�~�G��ԡ���~E֙����5���>�N�n�܆5t5\�^�:U�x_x�]���L��8}9�1��3�y�����K���.K����#Z*��%)����p�MsTٵN�z�����c6R���@)r'���ms����ҳ�0����E����fV�c����y�(�7:���bISn��&	kW��Ӈgc0cD��?�~��}�����4�#ϗ�CQ����;=/z��C�R9:4K{kG����/�!o汇N�c7Upk�i��,��/����cHծ��á�%�Y�I���Əmau49���b�2W��s�w>�:Sn���:���ˋ���l��wi�rzX�`8�R}bn~|�vt|��~ض��(�g2�c�4�OW�_hh��g�����'�t�L��1�T�C�[�����_վ��Q����ȑ9��.m��i��ck|B#9�,t��Y�U�PTF�{�G�`X�@�9�F�
��_}/9�!�t���Z)�f�ge��� )G�~��N�b��.�Sԗ�eYrr:�u]08��:M!y�m/�m*�ڗ�5�bY.���w�:Vup�5���~����Ց�QM������a$o�����#�9�L#Q����w�	�S�����z+�3�w`����%roX��_xɇ��~�	���t��ZR�8v�G�$t����a�4��C.���f�����LJy�7pj=;�)>�蟇W�Oژ�>F��V��i���wF���3�"�@��^
v����<����6D};wZ�r�;ˤaf���b�sj��l(�ȅ�X��
���Ʋ�V�]�[��GY+1���b+��Y!Q,.��qod_v#Y���*;� ��x�TU����I�R��W��Yy]%��J�O	��X�,^�V�
 ��|�l��4�4�(n������Wnr��8@�"�N�����P�WI"�k��H�þ
̥�Cvn��D�SC+�l@m��m�v&�,<�������(wה��mzf6����r��I�#j���G�3xd�
�R��>�Z�<�]�K���\eb�0�8�I���x��|�C���2�����������͵�Boh{>z�+�V��5��iIc/$c奔^@}id���+�.����.w\O��e�����^���^}��w�z����e��ĳ��gz���
S<ӥ��Kw����T�>6Vrǩ6Ҟ��z�ΤY�`xyyEíR�A�#n��3����;D9���/_р?A�YMϻwo��ׯ�ǏP��K�A?�(]�fᏌt���'�C��24
*o������:�f/?��u
ԙ��*!4�*��t���>(Zb�q`o"8��JC�D.x.��ʪ�W��kO���Z���?'U
g �ſ��T6�y�+�L�Ч�P�)
?��n@�/J,��'��P�&8�G� 4V�X 'UOv���e�MQ�u�m�eSau��
�=�"�����Od+�]N�$מ����C�T~��X���Y�;oǘ�e\�t2j%mc�!��N�r����[��n��`�����7�`��+�O ��k4�9�@�96�"]�=x��~ޖW�(.RT{]]ۄ��^��䝥��X��}�jO�_^�wyn��$�pՎI�*������8�0N���w�2f\w�z��Kg� i�LZ�*��n��gȹc����Y��1X�5�"�$�Fs净
�L`\M�cb��Q�T��K�2D�\�Is78we[{舁[��S�֎����n[���^��J�z;9�G�	��D{J})������v����Dq�	#�vv~���n�0��?{cj��C�eed�Ft:փK��溜�'܊ܩo�Un^����a;=9L������ �͚�]E]�>���X(�]�u�7��Qҝ6��/��w�C�rs�l� �*�����oﰝ�ӆ�o���t��b����8=���bp��G=cSY����A�t�������w/�_��o�W_���"�+=Y��<ʧ̋��茷Щm�,*\˙͖�s�"j�m��+(e�r@nΨ4��wX��H���Э�7Mۛ�Ζ �eKz��n��t��AΰI8�Uv49���t>�_ɤ~j�z�ma
�u0����$�=�����~�W���Ic�5�#�lcd�{�64���StM�ig�t��~]׃tR6@��v2�x�q4�u��7�+L	�3�W��g\a���O��[]��[uK�,�"�:�^�{�^u�� �����hҹ'�й����������K��=?3�5Y���ȿ�W�v0���3hDYAM6z1� ��@J��s8=���ɵF�D<�	�P�
G{?��j\ef+;1m���¡�j�Ő�(��5Ҵ�%���A�.X|�h�=\[I��Y�x ��i�1O��Bpw#YG'�i���Vo���
�'Sn�/�Si!��Jx�)鮙��_�J\�4�{�G�0��+>��0��2��v�o����S�1�<x�b�w��	@É|�*���X�`��$���-���y�+.��Ğ���fn8��cC:Հi�T~E>4������S��CX��[^Ea]\���p�Vi�5��W�^F��K���../� >����|	���O}運p�Rֳ2t�P�YW	�7[�Fn��K D_!%��1�KѪ�g�\-_�ýߓ JkW��PϦqgd�<r�_p�ֲ����ϯ{_��_�#��t�|W!�������"�t�?��}�yv0��ב�1뻧[e�Se���Թ�P�X�bL(�)C��SO�	��*m�did�ـ���j��s�$?I�� �ͷ���Z^^B�M�����>�޵ͭ�l�����o�.�>�������Wc$��Cx�'�2}�w�u�؝�\_��k#nh�a��j�frҌa�"��
���ʃ��y�_۞��
���>����Iv}�����3�RZlT�c\9��Q����%3	��n��Xd���P�#/�.�Qm�7i�������(��s�o�f=jȫx�� �]�+#!�|'?��ͥx�����������ő	�����+_�]���7�E�x�2[��¸�[��s��ϗ����v��ٶ=t��OU?���~��������s�@iK(���*���/,,�kXOx���K�oTb��	��$x�>����D/������u��*�����+>/ZO�%����W�V��xrt�qy�4�u���\.��,�O\�C~��Tjo1`�N�좵��ۇO'=�u
:�@QD1������)JEfN��t�&ƽkw�c���+?�%ok�m��=4"\��T��GKQ�O�O�F���f���O�ӧu��H�k���3�֮��%�<�o�M���SʵT+(h�^<mOP�@W�������R�N�w��u�����H�\[Y�/�T�)��(C�����;{����pC�i���>m{��"��'~7bp�r;�����e�@��'u��7a4 g1
5��u?; T\�ή2�������52�:�ɢ1�V��g�3�:���r�Ww�m�+yJ���>j�+��/������lO�8?Ey�>r ��� �=�I�]]#k��;���꒰�vRG<=�¸=��؇N=v ��OAe0�t���9��笺E���\�$!�Y��\�ExwR�PB������Gҙi�.p8�Z������ݝ�����3O��HW�t�JX�P�Iӎ���e��w���xG�m_�ǁ[��ֳ:�S�ō����s$kss]y�>���;�'��0�d���5������r]�yo�d^��}`�� ʘ��(g�}��Hޥ���nms�'<[=��3��D%����ȃ&�t�ק-�Q��|����Î��X��n#��	���ꍬ����n p4�ԜJ�HV�H��C��2���K����^b3^?%�M<�=����2k�T�كa#TJ��SK*F&�(��S��BM���~$�兄�W��3��@���7���:#YG0�FV?���r�d���-��q��UeM���CgSů���¡�N��rl�s�G��XW�rR�c{Acd�'d�n% ��	����2��ח���	0�� Y���8!�0WzFTjd ���e�Ը����	���z�g����2T9ep�G��8��Fم����W�#�:b���n�R頦����P8XCc"%8~��QP��(�V����G�¥Z�UwW(�=]%���Z��������Mp�'t����
����{�L_Wn}zU>�'F6[C㥷�+S��7D�|܇���s���3L�R�J�{�_��'ޛ\�4	vΗ���w��g)����"L�Wҋ���o1�{�+���㴎ɩ������U@1�
��wg�ꑭ:�s��V�؀׆��w��܄G#�ڃg}(k4����r�͢�IҸh��;4t�(.�4�(�(M��͋O��+ �W��x�/�$p&��ą�5�:���o�����t��բ���j��C����ndW��6����jW������o0"��,G�\#�A�M���7^��1����&c�/GFz��@M�"���~5h`�S�4_ʈ��x�p�rf���M�YY�zE�كyё�#�y��x������1��n;><���ǎ� �t��J��Z*J^��T��ɵ\K�z��+y'D������w�+���먕��/��9FU���R���m[�c{�������yw=#[�G�jXM;J0S[J{��TS33ظ��1� <��^ �W���T�8���"~�m�� .9(��'���
������³?�B�|�ܶ��o���WӢ���N�<C�?;u�9���S�D�W��6W}�N<��*IN���iGg��x�>m]Ү��cLg$��Bڰ*a2�	����$�M�_\G��Ȋ �^I����Z��P��a{����m'����洸}�e#KC�Y�v^�����
aq�.�]���F�0���ŹY�'�.舖�~��|��&�im����gk9��uYl�B�w�;�?�ǩI��%xF�9��:p�@p��45?K9f���3ۑ�9�$��{�=����s�+Fx4�:��f�#���.�C`L!�cP|���޾��.0&&�=WjڰJ��T3fT�]�#�{%��i�� ���[u0:��O���_��߶�����A7�@KƮ�9>>C�;��qO����=�-�$��S��sڎ]����j?����~?�c�S�Iif<mg0�V�$Z�������mll��>Ű��4dk3� ���i�������ީ�G�Q�t�{NdM+,�髻V?l`,}l�z���i��G*C�'|�������(�����;�}�./(;�D�x�]t(`r�9�$.�H�\�����0���q7��$�d)�Wc*�p$	�F!�ĬY^$G¶��!^�m������֯�^�;Y	W����uiv���W�o+��!
z�����b���ȳ���uS���L��q����6Lm��]�wn���1�T�6������fw���{1�N���2�a"P�\SS�u�RU��	��)L����:������t�;���^�ש(�zvԣ�r/S`�G���<uܡw{
Y�h[[���F��.h�J4 R�2������j0�F�{���n�^F�J�����L5�<�0t���H0�*Ч��{�TX�O�Օ0�@���n�>!�x�@�4�7�('Y���+���#���M�|`5�i��L���,�Ճ?0���0����<�;��.�{!�^�#�\y�����(�P��N"P���e8~��V��ܢgZ�V�<��_�VO��b�",d{M\��o[�:�~=XzG�*Lq�!M�r�4�xT���p2؀k|SJ�
�� �}j�W��>�������^�^/}�km�oʝ���g�E���lH��L)���ըG��x��b��ݵ{W�'���8��&�t�'�l�]���{a�7㚢��ǹ�+��J9S���x}��8�(����zW^���<w߲�-�F�FOv<wD�]�0��վ�jM����B'��� �K�9�Yf��twur+l�Aqz�=Ҧ���J%�o`U=�#y�A�{����w=��Y�'h)���x��A9�H|�N��5�ߎ�lS��lŀ-bq�w2��VM<�s8���7�h���_��_}�5X�"�_��)��̲�F�:#��)K��|� &�$�O^�V�C�F��X�4��E��;l�|���?�ZrQI��Dɣ�r�9��
ib	�w��	{�L?D��;j�{�������0��E�n��0J^�FƜj��8*x�1����Ȣr��<K;ښ�"oI�h�r��%4qN~VǇ(_�mg�#���:H�����Q|~l��߶��-�[��� wg�w˻9J��8��[��Ev�s�#��>D)_|B�<����h�����[�	<�%N�&����}}+��.���{�����؅�"I|W޺�<4�����\�U[�v����L)�^�/1�x�;����K�C���/�W�������M�`b`]�(^�u�F�q�,�kӻ��aT���|�F����y[h�`G]ݢ����Y�_^���@[0(��߷���Ȣ��Ù33��+��Ϡ�~��W�/���t����)�:��~�u�v���nA3�G��ݨMe��c�ܵ��::�wJ�S/���_��Ht����Ծ�ٶ��.x��/~�����+.+x���m�C�Z�RO�ĻB֖��,(%Ovݑ�W���Nĳ�d�Q�(�ˋ!o0\< إ�d95K��2]�*�!���1�f�݈����Od��o����M{�l���_�� $@ۿ��?�e�M;I"�m�-��-���'���PA�`��ܴ�����{ -��?|�����������ߵ���߷ݽCj�8\G�I��2���U��9l?�������}�}���@��hhbܩ֎:���	<�������}��O���6F�A�w�a���I�yxx��|���ᇟ������Ǐ����d�I�o�#������]���Ay��h����������4�}[,�4�M��F������l�?~������W��(���q�)���md��V�_�J�_�a�p|� �X7�|��t����r�=w�_y�R'hf_IȋK� ڹ�����D�Q����4h��<��U�~x�=���˘��$�:��r$�-ܷ1>N�d�70T��t�T�wz��BIE��3��l+Ӟ�)isw��S�x^�(�&v8�|��kU�>B���vʙ���W�\[�btNS�d�X��q{�x��{�CVY'W1�O1�N�_�Ԧ7�J1h��T��V�Y�?odE9'��V���y��"
.��}!�}��j��iI� a#��H6�(�K#��j`]_�g`� =�,
��'J	ēE�x���p��ރgg'�s��4��Rg���T�M&���ְ��Y�!!X�ޞ��m'�Sr������N!�� ]�0�:�	4 ���7p2>▴Z�x�ε9]�Q9qf}W���"e�޺��H^Ĉ'p�7BA�	G�{}yY�$O&I�sUm��)�\�)�Y��)��UiV�X�u��EX���C{>��4�����k��s*�}Y����������O>~/�d*\�-���k����սoBo�Q��L�֣��E��zݡ|i�K�Ҩ�:��Nѳ!���Q�1�|��ʢz�g�1��uݚ,�#�K7�� �����H��N��P9�����e�
�=VG4:�{�mwg'���|)�}���/ފ.�ú�1����ڇ4x"�+S�Pf;��gM$�FIɉ���;�Fer=Gs��k���o��XNEQW��Q��!��х۸�(��|�`�U��2�N�S%54e1��_D-�7�<�q���v 仝:c��d�غsN#Y#+S�Q�$�9]�d�x��#���]E��:x��xtЎ0���^ӫ����v2-�gG�PRUj/Ϝ��p�l�r7ޭ�=XŖ��Ӄ�;: �;��l{;RP�޴��(D�D��{��{���o�:����z�p]\Sϥ�LA�U.Vςu��i[9�v�^}�.WY�ƀ�D�.�B�+L�p�>���TQ����<E>H���Fյ���דּ�"]��p|�sh@ڃ��?��i�wg<��Uu����,�{�S�>N�TkJL��%y��5ZjG(�8m��J��y��s�6w����vv5��>
�`��h Kɛ�{|�4��j x�����⽚�*�[(���4.�w�[h��
����:��^���m㮑�������Z%��@e�k�<����i��ͯ�[~�S�v���ί1v~���붶�71֎��|�,d�m��ѶJ=c˩�Xg�";��1 ܖ�N�q�r=�{���+��Nϟ�_��71�4-�S'��3�S�����z�nα�|\�q��i�>�|��CG�����r&�u�(���Q#�̬K��������Q�����3��{�=d!�\�E6b8�-�ܶ٩a�ӵ�����_<͌�n��Y���F{�v���f��Y��������O��H���;`���C���`��!�����?h�:�����~��^���^���}��}����C�a������M�6u4��_c�B�{mg�mm�c�l�Y�������޴����2ڮO��O��ۏ�߶��Q���?������Ѭ�cd��32���C���'`\oo�Q�7�}���{��������sF�5X�^*��B��>�S7�����A�f�(��1�#P>�Uڏ��%�䷤ghY��O�'����3?�ӎ�^}����$�i}��]�_����w��%:�$��4�Z����k��k������z�J�7��,��%�<��:�Ӈګ�����Y�z��Z� ��,���;c�M(#Y
C���"A��mxS
Zk�nC�S46Z��G�IO#K#�w���c�(r4��W�'���n����n8�#~�x9���g*� X`D��1����6��u;:�5Y���`Y���pXa�GJ14������UI힑������ȯ�*�FZݧ
�ݗAe%��� W++��+�V�0]w;j`�/Q�0��nϫE7���)!�;+�L���v�����@),����<N�rZ:r�He?�SU^TxTdd�"��E�z�t��t>��:7����$�4
���eR�jz�M�0��W��YП��Q�
(�cX��U�V�Rk��W&tQ���Fɞ�̃�pQ@L�/F&�4����G�������^k��/���e>�#�hS_�����$��M�L��Fz���`Z��`��K��_�"��F���*�|�+ta�
��8�W�뗤��b��!Ҥ�G���څ�ѫ��u�ᤁ��WQ
T����z{��3�i%5��Yx�H#@d#�PUH��eQ�x�;ﹱ�����	�=�;�;u~�1�#D�c���̹�l5�T-��K��+>��+�����؄
)y��|���l���>���C�C�Y��`�Q{�����7��!�N��ĵyq��k$�3�Tj�
�!��H����ڬ'�[�m�@���2Y�.:0Y���+#K�Qٶ���5���e=��q֑�溚1|zJc`y���t�!;oK^9e�-����m�]�!G�v�?�]�Y7��r�Kc��0��w0�Pf������@���jg�c����i�m�X�)ރ�70���������ow�6o%����Zw�s�Ý�q���^�&���]�t�C�k���Qh��4~tl�R{�xT�!��Z���j�*��;�œ������Ϲ^nH�%yG�r�9�;Zl�iߠ4�Q���F�W$��m�:y@5�R��_�d��H;����-?�-�An�W(�W��>vGq4إ۽q�صRRN�:=à���)+�Trc�`Y
lu��2vᡕ�'�Y�i;o��e���$��x~�S�Iq-/��
���]���p5�u���9 ��W92�C~�;�8�Xq-�|�`�SY�m�(M��X�4�����n �XG�NY��ğ�kKȴ��6�������(R8�ȍ<\gv�|�v(Sܚ�]W��5�ٰaX"��[���nݥOw��
���]��n��nh��f�Z�/���3Q�;G[�'�C}�O�,u���K�О>Y����}��ﭹ�?G���C���+Uo���X���G��>�~\��:u���o8а�>�o�B���W�|:Ű�@z�1��q~�Lp�1��)���!���:<�}���M������������یJ�~�.FW����Х7���G�{G�7�����m�����6��A�^;��>@��Ȁmڤ���a�y�lC�l�N2rJYΐ� :�a(mW;\����-�u���� mC�x�[o�mA6b��y�������C�L\_��]�s���2�ڮ�W���Oy����[e��q������%��u�~򲽵��$� >��W�"=�a�I{f����/nP�/=����=^]j�������7uq����/�*dY {��@��;�P��{��#:�8��թ=+[�;d�D1�0�L�)>���ʀ���C#b�#�����Km~:GǞ<z؞yq6�p�h�,w�>�^��G���5wE95��cd������E�GyN��v$+�Iős)���TD�R�T`*<꣔�ǜ#%a�M!o�gKE�[sp}u�5XY�$xuѭ�r�q.�HFlҫ���6`��i*)�<#���9�����JԞS���ڛM�ը �xQ;Cc�z�OWQt�8����a�qJB�X��-i�u&w���N��l�E�'�ۛ�hVz��+�S$�Rg
֌l��;�+=�5ʢͼ1��` T�e�����m�w*,=C���u<P.S��#� ��kn�g��W�p�:���̓�"(~�=ጰ1w�x����_>Apҗ.07����a�G��%W0��}w�'FG�A8�w����׼�_��'n�Q!�;J4�C�X��[���dʞ���p��r�*��bm��%��,�v�����ʡ�+_�_���hZ��2���#���"�V^9�"��7?�AB��NbhI��#y���(�)ϊIB�H����z����N�gT�E�he4�R�����))��O�x>�ey��7���~ݞ=�
~_��5�I�u��BY�Y5�F�%^�f�x$���u����s���	��*dv��-�:��I�rc����v��hc�������N�6K���tn��hVXz坝:cî#u�r�>2�i�gԕ��G�\��<;m?���^�{����������ם͍2��eTa\}��;�����zW��z��`s���v�7�]�x(��;[�;���1�mg��4.l/�25F�ak`pM/�������]K'�#�F��R�]����*����MEy_o{g2]�?�B�W���e�1iŴ�}i�@�A��aG��]�r>59gL��"�� &-�UZոwd����m���n���#��h`�};J"�C0r���s�N!�"Ci8�7�B=`��~�,�����(3���Y���-�A6��u�ڏ����0_G�=���EKss�ŋ�9�V�Gcf���Y����_>�7�X\X�q����[�Ⱥ���&d��٨��g\g5;G[:��R���.�p��3K�w��v]�U���q�Y��~��V��e�&梤�+e�ۋ;
�r�I�� rM�G��7��ߑB���z9�ʺ��#�]��ܐ+���C�uݭz�����&F�������W/��2��R9G���:h?����v���z�~��n����O]!˷�b�^���㶟��Kt`ې�mn��(#D�߾Ɉ܇�b1���?�H�@�;�E�𷻋ᳵ#�i�����k=�/�����)zW�@��Q�{B���>�N�C�;uU`C���K[ogԹg�jdit}�=z��}�#nb���ճm]�c��	u�+Q��g�hI��H�&rNz�$�d�����������Q��+lo��<%��ī��x�z����a���O��D���D}I�r}�8BU�ܗ��M��-���m��0���j���h�v֙^�$�Y��m-N�)�C~T�L��P�M��+����K��GK�m�3Z���F+��H��;V#V�� �jML�x�)��rb�Q�c�C� �'N��a�5RT��G���
G(��i0�2��@����HT���Q��X��s�*���E>8��ɑ����
¼j������.x$��[h��(0]�v�[(/DK@U	��p~�u��0�cd(�@	򝢽<�<��]Cp��\/Ov�Ⱥ�I�7W?� �9{��"E��Bjdd�z�7�ΤC�*�=#�Ӝ:���mee1���N�
��+V	��el���/�Yh��\��T%���o�=��0�&��JrmL��+1;��Ц����aA�{~Ȣ�o̹#�dz�����C�u�oX����_h�2�5xv��81��k�ƿS��ȝ������r2���׼����{��W?�[ǆ�K pk�A�r��^x�q$��YI�9`��!!�\�V��d����.�<��Õ�|z&ӽ�i��4:����(�y���4���ϡ���DGm�xC����[�C�C)'(".2vj�FF��b��P�Hkgd�I����w2��j=S�#-H�l��:U{��(��R����1[_w����2�,�p�ue�����'E+�E�O��'`�%Y��=g��]B^��)e=.���O�-�uc��Jev�lS?SsS����oݾ�/�>FQG1'���M���_��k`9b�ˑ(��Q9I0r3�+��^�~	U����8��U���q����r8
�(�k��#G{�Q$Ļ��=��i�S(�v��^ĸU�)cP�=O��.r��ӎ �u.$5Bv�N�Υ# 0~��hd9ekE��.��[����v��H;�H�p;ܦ=�C���_YNT`\g&�ӑg821=�Q{��{P�Δ8��N�^}����J���L��Yh���yv�gMˣ�J	�ff=I�_Gy��-���������+\��y\=M�9��[1�����M����~#�h�#K��F��(�4��3.�ى@��8#MI^�����E����:Dѽ@�"�b�k�W��NE��8v��F��7*��S�#�(O{F���)���s=�y:�������������
u���__�˜���l�62e�4�Ww�#��}�(�oP���#����ڃ������ۇ��w�����o~�����_����e@^l�ӵ�D��]#�v3�d�ce�2�ܭ)�:��IH�rkX߾s�܏���>(�Ewpq��u�u���ӨW�{��x>�c�y9���~��q���ڻw��'�,GS�?"���qQ#��%/ֿ�$3&]b��B6�Z#�<�,IrE9G�E[Z��f!ϟ>�L��Vw�����^�������q�M�w�r}O#[�2j�"��~����K�о��1wN�;=sGj�O��7D�<��v��	�����Ԩ��1�=�(�[Ϯ�^qב[��-�a����b�A�Tmu�Mu���`��[�����ݽ=�tg�9�b�;�[� :��@#Q��uV�!Y�/���`cL�5��fm���
�I;����*��.��Q�:V��z��sYR�����k.ƭgݽ(���_{o��H\}<���gm�	neR��(���x��h/�7Ku�N�>Mi���峸P~9���.�>\k/?l�n|��bd�������}�b7w�&���Bq�]K<
 *�j{�Q�a$�,j�⊆ОB�Kj�2d�e8�� >����4����aK|v�b����{���0�潖%
�J�==���m����U{��r�Å�䑎�l|�� ���E�,h���3�,ޝ�@���Ɨĸ��Py__$C٭5.��;~��	HI*���G�J5<Be*ȃ�(V#�!�Q��C�!�ꫳ��<��Z �ߢ�8����im�����=�7�J���w�Þ_�U��=�w��Ch/a�,O��U����l��c�\R.��u
r������'/�nG�=Y;�p�ri�N��Y��gO�u%�F�*�]=}�-�(�Ј,��.M��ř�6�FԱF�uMn�E��ܥt�t�Q��h�yҖ����ѭ�����{`A�<�E�z��k L�k�B�s��L����!�:k��]O�I��D�Ȥ*�)�7��0��]�P��OZ����r�[]w�)�����˵�Jd���_����%��׆&~�5����fZU��(^&֥ۥ_ӕĉJ�x�*&5]Ե��`�}�V|ؠ���1988@	@�� ���	����V�����{A!�tS %�t��-(|U��kz�s_<D���S�	rÓ��QH>}��do����ܢ�У4��u�����7}���ʃh�xW��H�!�֐�)|�1�������4��4ys��Q5�'��5��d�_�W_���|�����9��kd��S��Ho��7N�u]��t��7G뼣��o}w�-�*x΂a��'×���U�hQ\J��
T�N\R>��Q4�%کK('�`�F��??f�|F��rnt���&iT�7ծ��[䒲<x��N7d��1�R~��seT����|zze��5z;���Ȟ~{�]L�w��-iޚ8ŉ1��K٩[(���	����#jL�H���U�h�H��rH���w�{��4(;�M��oנZ��9<�zj;I��B�R���\S�:$x��ۨ�
�����v�2������Д{t��F�{���i��ܐ%>�4.�bwFZ��}����S
vq3��h��m�-�7ۇ�H��X^Sw��#�����I���r���(J��ǌ�^ߺ�;����@�(�@xyW<)��Ip�ќ��.�;�����1F������;ƽs���(�gЫ�S3��E=���GG;m�`��̎��Hϝ�.���?���`�o�ɱ���ѓ��ɋ675�<��sM��hck��bdOalOMyp�<�e����e�u�D*7-������1:�o��w���Oms�S[��8
77؇�1��{�-�e��#�ӓs�{y����P�YO�I\�əm����h���}��B92~}�A���w�ƍ�3�-~�Q�1p6>�F'���I��_�IH��0���;���d��҂S)�7z�z�9��ÿo7�ڛ��m��S��(4 �\BWY�(��m�l�&'��2��h4�c\]�k*�%�|N�b,A�����D�%N̒�;�N��/^�7�R6߾� U�55�N���rJ�����3e7��f��r�[v�D6�A��0�	ϟ��#C�j^�t�_�p<�S�� ���#9rsx|�66>�ׯ��ڎƝ�4d��Cz���lc��Kv^�6%尚��~ur��=��o�*/Iĸ���>�	����
U�ſr��۞��"��)�\}�}�/�u�� ~7���v�a�0����ݶ��1�td-��-�k��@��A��XYZ�,�+`�Ȓ�����	�w���)E�Q�>+��P9ҥ1�rj}�
�&A���&M��W�HS%���F��	��������b.o��+�p�gQR]�*Q�o�.l�u��}�k|��������jb���Θw�����@��e�B���Oi���r���	e}
����<(Wm� �*)��PYJO����=񚆤v��i�NEXʢ��:5B���!���)���Q4
��/36�ЃĬ�0��A���n�ۮg��f/��v�FVv}�]� ,g��(��5��E�477���\|�_p��i�go������+�ơC��Qq�(�aQ������&=��>=G���e����e3���̧�P��sw_�B�L�(���A|n��W|O� U��a�Ĺ懶������(>����pa�1�յ���i�q��3(K��u���p'S�����'ߠ�2�I}Z�K��w�'��������*����}�J�2+��lq����Q	������O;�oLCy��{��E3\z���?�*h��F���2����ԉ� ���F�x�`AI�e��������gչ#���C�&Foc��+�&0��s>~Q�r_��Y��u�q��
��B�lN��tf��)r�Er$��5�(�ݎ��Ֆ�m�}J;�;j?��s~�w������Z�TSe�Q��Eba�SkJi�xN<#�{��D���5�ҫ�q�p� N�-�1�[�TW�)����:��W{�3+@:�#���E��IӲ��$�Z�Ѡ
m�]_wX�cg*�����L�օ?����+��%>��Ӌ�L�r
������^��Ő�����9�(pFxI�.�@8���Hn��n2�C�]#���9|�>���KiU���*�}��6�6�i����d��?uG2n[b\�X���IG�KO[{��?��}�������i�޽�TA�u�_uR���S�bPa�x���J����������^����q�6��2������������������5��Qbא�k�Q�e�d�y$N�x2�v�y�˹Z�������z��R&uDqU8�[�	�I/
�D��&B���B<�S���d~��������l���,;����|IL��.w���#b��L��F��5��K���3r��%G���W���@չT�6����qG�y��uz�S/��~YE��P�eipg��YFy3c#��)��z�K7�,.�Q�}������H��l���0��������{�����	�q�`M}U�!?�e�l����䙼i���=׻����i�����,���w�����+��k[�>M婞�C[�7O}_���	m#	Jl1���~��"�n�q��Sټ�p#M��'�v�g�`�;mT	�)E\:q�"+�J��ՐU#�B���4�F�	5�
��(�gC �T/�0Ј�MHT���:-H�X� �������I�������2�|�Wl�bP�~���{�T���;#?�'�J/�S�#�S^�Z��c`� �������	�8�ZX�N�4-���w�ȘN����k0�8 l�#(2��nێ�^Zi�˫mia�l����؋}{��o/M��"fr��п��k(���@��������{���l����mo�S���:��i'�K�6D�<Tx[}'~lLz*��M�)�Ň�̔�%�`xIo�@7^���|��!�$����s�͝�\�Q
�#{55�h��,�Oc�CN1��|$�4�G�Sh{�}��U�݋��]�I����u��B���}�@O��|��d���[R�k�ß�	Ӆ�cG���u�g_��M䁲C:��=����iiP���?�+z.W���4�I	�Sݦ��2}od颼�xtr���U:��*��՗#�/���F��e�h���9YX�gOe�V��x��=���;5�L+ûQ�J�#\��6���sm�������<P�����|��|�{�R�����|qU��J�\w�#g���Ty
��dZ�F����P ču|�5��~�pթ�g"C�cC��*WK�ꌬ1��q�5ӛJ�ovN` i0i詼T矊[M��s�>�xԣӘ�+N�2�>ky�#�
������sG����z�m���⛷ƨ=ҝA�ס��s�k���t��r}�gx�:��y� S��{�7�N9��Qd�����l�ik���ў_�6Z����GAӑ���t��A��"o?���jȻ�E��ȥĕ�Y��5sbǅJp.�TZ�ب���nt�M:\����꼉����o߶���w�>}�L���0ч:��T݂7��QLG�0����������,^�G�5x>|��y?���U>U���A�y��<��,�
��
�S���t�֣���O�YXO�vp*��_\�sy@�ǎ��q��͚�V:����i��@+��F��Ƕ�9mYY��j��'�^��7��h4+,���G�҄�+�t#�p�,s$X���oЫ��A�av�����PQ�r�q�8�NcV����dgIE�0�`�x��v»|�LӧS1�_O��UU���d�B��}O���S �yթ�?�ko~������u�gw_�Ŋ��]�l���S���
V雷��{g��o\�)W�(#�V�}��dnᥓk){PC&p�FT�c\QW�����G\V��z�$�!���Cp2�-4~>A\�6�q�:���I��TVӾ���E����8�-�P]@?�c&�v�s�Eڣg�g��BGp��4�X�
*�&.B�ѩ��bl({j��k�H�;�c����C���]���{�w
	b���A�ҹ���.a���kY�Ǯ����!0�J9){F��"�L�\/.�к��G�ψs���	�`]�䞡��pѩBb|b:S��ZYZm�+k��ʃ����9��	`�șub#&Cnx�Yf���k=BRC�!TG��'��`o;k�\Ӏ�u���ǻ����x'�E�P�\#��QN}����G��!`w��p��6=qK�7�Q5��'���t�;�}yi�-�η�Z;�s��U�P��Z�lީ�]cH�\��5�(����SZw�sa���8/���q,W�������ť���d���,�|�C�.��w����_��o|��
0p��[��w]�8�������=����<~�pVh�VK�V�]Yy(��W�r�/�sJ�;1�(�+[
D)Nw=�w��������Ѽ	Z ��	��R|���c���VK��&-��2yFC�:ҽ�S�.d&/+%	ͅ4�Y����OC��]Xh������J3�ahh)+���z�;��=n��w?������_�)G���Ɍ~�#���X�`|idU�����aqp��[<P*�ʇ������=���f���u3VA)Ym�l�T��2X��C%W��M,j��rY�*7�Vƕ�b�E�OҊ�g:���%�����0��Y�K���ˮW�A2U��V�(����3���^q	L�!����D�����&�q��B���L|޶���������D�� 5�)~��u'֧�U�X��%K��Ć���)���@F����еt�myy9�T��Mh�s��i��l��\(��:�<�G�A�a�k��~{wg7��u��?J�lԁ�u-J�k�OpH�.�,�����!��I��I�~�뉎b�8J&�h���g��Lg���@u.2���R����"�K/��Ұ)���[��ط�)o�~S�h�z�ii@��4�T>��;��wPh幢a(|8R��峺� �`x��Q�{Œ�0:��c0�u9u(��ݠc�xX��u�Zi��g:������t��BN�*����w�{d�,��SN��6�y�r���s�
���W����-Y]8��M�g��+}'�%Lћ��'�
9i�\�3Ӵ�Y�H}̓�7�ߵwo_���޴��p��j�=D����X�zw��y�7��������}�p%O�=��7�2���M�\�w1���Ai�G`�p!B���+��;"�N��Vu��K�G<�\q����0߆41��PE��8�1��;�d�i�>�g�)��Lrp���s�����Ql@�Wĳ ꙙ��XH	���J(acd�Ŏ�zN�Q�q+Қ����9G��$�kj)F�I!*M^Ǜ^����I��O�X
�r?eIz�W<������Y���K�g$�W�.Ěk�R�q*0�?0�\��{F˅Z�/�I?'|�s0� ^�<P��J�;��$D8���<��L���|[\~�VQ��y�3F��F�r�����5�!�j�b֦#Ë���>S;Ơ«�5:��gG�<�p�������^�a�nO�y4
L7��W�����7W���R���s��j�c�3�у����Z{��Q{��a{@ø03�f3u��M{FҦG�x�
�sw���G��J!���2w����A�ۥx誔9_��{P$���_�pw����%�g��(�\�np���=�.��G�/�Px��T�g/�;��p=hgZ��4�� TP���ZSYh<�i>�����c����%����fe�
����� y��p�=h�oUA6�%�L�*�*ؽ'}a��Ι}od�	�w��ip�JT9*�����̯?�j'(N��٠�wWז�i�Y����S�u
𜇃b`�|����q�~2�hco�J��; �����>�����8�.��Sc��"E��(\�F�`�8eЩ��+�����rS��}�X�P���v���&f'vF���uSƎZN�V6�)�1�@I���vSxީ�5�o�ԵKv�������q͑r;��){�!�z�+#q�_kR�y�qu���4��g�D{��F�֊�X��e�c�L+E�uU����9�X�H`��&L~5��0��5Ů]9��iGmg�4k��0�����m�G�M��K!��1���H�uP#�ƫ��|��k��2������� Y\Z�q����{�k���8=K��mW�x��Lz���.�o�9�^�SGUk�W_�ʆll�)���<W��7���hL(�ɛ��~�[�y$^4=�ڭ���'h���04?�'�Rʴ���úT�����Yy���4�K����ö���F5v�����Z���0r�����Ex�������
�� �.x��<�P���6;;�N��r�;:,�#�����x/Cγ�j��c�rɂ��4SF�4���؁C�s�"-e�f��D���S���� 9'�<����f�AY�����AN�t����v|�����l���6�Y�epgeQ;��2��P�Y���Zo�Ѹ���%�\����O�m���P���e]�I�׉kӐ>J����o'x��޸���샒ׄI�^�`��ύi!׍��9�wֱta��O/�G�Wf,^j�R?�Hw��S����芎A5��"�(�c���xB'��G��c��,��j��8t=P�b=��w�����/BTw~pAb�<�J�[G��룓�����`E��j��ғ�1F6�~�B�S�v�t��[��ޞ��(�Q���*5P��s�o8��2֕��[JU�V��7Za[đt�K|���߻���Qu�׻��!���F߲A�#���o�O���h`A���C �"{��t�1�1��f��T�RV&ڔSh(��匱�"��@�e���Top�bL�gf���֡
J�g8-J�ԫ
�umo�om@Tll�ςW�pt�p�>�0iT� T�g�k����v��؇�B{������:oc�mfj(#Yk�s�ų���7�ۯ�u��/�i�����W/��j��8�G�([*wk��N%��'�!�u�>�����[�
=���$P	���ep����Љ�E)�Q��O:i����'�S�^�wE��P\�\���ߠN��_r]N���:@�s��W��	�"O���{�Ëţ����t.��ӈHoq
e��~�'u�EJ^����HS����(h��T>=z�]����pM��F�)�N�Q���"_��/K�UF����w�劰P�ꍃV�V�Y]F���onF�l�����Y�'.��G	�|�q�t�l����,F�b�@O4�T&�7����Q�"���C ?犃;���Z����a���\� �o���!=6�F�Gv�N��Q=� ���p ��p\�B�Jܪ�h+���� S�+���]���X����������7���F_��z��{GJ f��4�2m�Q�Nѯ��.���ҘS��Q�N0�bdi/����r5^ᬓ5�*��/k�0�]DYu�/��~��I�Ǻ�N�(�I�Mq��%�TY��d��kǧݙXۧ�I���eT��	��
�r�����HGvrt4�]u������4���&Sc��z�Y�t$Z���RZ��רAhC0��'�>#*�c:k���(=iD�I�:�ݑrT7gGx2

��I���]�R�x3��&�ה�#�i�f2e8�Ë��:��)�G��UN
F��ʩ�F�,��-wV�+�����tϩ�s��Ϟ?kO�>�,5y�ٵv��%�w��vj�����tg�8��'Ntˎ
G{T����ų���~�� �a��K�����&{�K��)�ch���,�ӫc�V���@�k�e�C¦��qd)Fun�6k�ԭ�-�*2������eˮ��݂����B�V����^(�rBy��g�߰N{���a��W7���;�{κ:�V:u}����v
9`aY5\���|{L���ǜ��!�̌f�y�/p��:,���o�e[��S�8BK>�Q��$�{=�{ɲ�7P8y�C����yx\v��d�V��R�L��Y����_=gݜ�L'�"G��tO�y�Q*bܑ�q�u��(e�N���� �	 �n��%���N��/� ,�r~�/�;[F�=~ګ��b�f�V�**7L� E�7�#I�qc��[v;���=��'�	�Z�����n�.�[D�������`�k���&Lʅ�
}W%�p�',%ї �G��U���{��k~	#��$��+Tl�k��g�+����R���!p�-Ƴ�E�)����q��e,8���m�����\[^]l֖���Kx�0$aܮV��������L9p~u�C��+V=Y
��γx��%�KXe��}�;N�%�-S�\x��[+{����r�͞��m�l�ӣ�vyv�����lӓ�mia�=~��^>_k�~�#�E���~���/�i��A�jϞ>n+ˋm���U=�Na F�,=5�:q��
#�Ѵ2������)�m�T������-_�����9頯ҿ�=��ݤ�������}@��ʳ�σ�GN��YWٗ�>i��R\���'�����o8�ˍu�4ϙ6M���p���s	��ͼ�N�?a�<��j8ٛ��&бa�����'��j�i���^�������:�^��ٛ]�~'C�O�+���n%�k�Nث�t^G��:p"��G��:��nVg�x|~������%|y���h���H�R�P^G�������5Y� @��PI��ɳFD�^\
�������=^{�?���Ia�uo����s�x�m�ʣ��'cN����5��#�YeB����wݼ�s����c�d?�P[��R�
�un��=�@��B��*#V���{��%�$��������L�3�*]C K��d��
����>�X�*�n�`���"���|�"y�Ɍ��l����z�Q��� ɫ�{���2�r\�[�ӑ;c�k�H���*�'!�i�2�<d�����"�qq{�Q� �W�(��vD�R�.�)�������\�9�u0�&r��*��Q&���VڲC�F�9�@T�H��]�2�F��v?]�'TJ�S�%� �줱ӫm�G׸q������l�蔰�(yUo OԺ5�q˘���\���u�
���} ���</�ꤱ�a9�!��۰1�������2q7Κ�s�o���:Uy9ƈ���Go�ф�� o��S���$�Ө�)�v�O��Ƅ����|{��e���o�ɇp�4�M!"��8�uli3x+��4ǚ%��p��>k0�<|B�,����Y.v� ���`���׵��%4�;����0��]fT}�4�[��A">�B|��G� �������F>�H'z���|FQ^u��ѡxҸ���o��Y<V��hLÀ���x6���/1��E-��_8*Sx�u�b��r�$i�`��>Gg���#�0`�=u\ᄭ��]��6yG��˯��2T�:��]^���(?���y"sMG�q���݃kUiB���K[��]�2��75�4�lM{�ܺ�~8@
�W�(���"��j:�{�;#��m��;���  +���2|됻��~*�B��4��?־����_����_����_����׿j�|����ں}ѡ��)�S&*�*I'�=���o�T�*�e�oy'�J���|�=�����_���Ľ���:�I<�y	�LG��e��C�[5]M�.2��ׄF��,�,&�jhu�T�h��(XW��1��W�r�gb���n�:Q�4�!*&>�w�lK{X�[�:(�\Ԛ).�s�����вQf`vjH��es����C��{33�=#g���`?;�0�sjrF����V;�T�����7�g��0;�,ϵGk�����B{�b�}�����_>o�}�z��a[]q����g����4�J�^����>..��.��V���������������q����������O^:������ +��??մ��_Ζ��u��zuw�ݽ�垞'>ˏ��7��D���8�P�*߾��^�I�Ӎ����4����(S>x&Z�U�{eg�!o�Qf���ީ'�b={�,#��*$��l���14H71���4���w��>� i��o'������)��^vC���G�kڠk��Y;�7�j��~�'�Yc(kS4������@1��t�}��|T	䋾4w�w��~�?���m�>[R�ow���RN��Q�&�w�%�.+��U������pR�A%Љ���*�Ż|7[R+�
�H�F���6^���_�7�������XO�I_xx/���o�:�K=ߍbeJr����֒��^g�I��P�B��/0�ԃ�hI
��/<ë��__�����l�È�d�aFW��	�#]�0F04m�5���E��o7S�e�v^���Ҩ4�I�X^;�4��I���ws��P�HF�//MH����I[��-�('B��K�W�8�������oǐ-��V������w������a]u\<��
�H|��0�[����1nR�ipU���q�����Wq-٦K�I���=�~h�b����+����Y��E��Ōn�۟#h�˔/��h��6�F��wP`�S�����ٖ�{7�Y�w����NL���ԅKV�!�k��mƀ�ח%� T��k�QN:ʄ��%���!v���eCu�h���5b�S����/��0��1GڞuX�=M[܉�·Uǳ�)/4C����E��4g����2<�)4 ݬ%[�m��hɇ{
4�;5nŻs"<�=���3t�5��Jd�-i)�S������r�Va/��t�s���<�L姺�Y�.��Q?g�W�,`�Yo�ˈU�C��򼦈���~������5� ��h��4AG��%��˨"u^�#��Q�T?���
_w���$P�V�q���N� 0i�,��m�B�2��x<��믿n���o�?�������?�'�����O�?�'����_���_���z��$[���d\�E��pK�\*�������T��@����"��%��'�φ�#�dY���C�����a�Eʤ0R�(���H�۫_^�-���qՀ�[�m+V�V�+m��2�C=�E����3*�!j��<���tA�QPlpj
�=���BA���,}Ξ��9�c�)?�	�����!S��)wC��*�������ڡCko�[[�;U�wN/tN��D�,�#3��s�man��͌`@���8��̶�O�0���Oc�=lk�Zx\�o3������������g��8K���N��&M���3����ۿ�K�V��P�ū_\{�0�݅ϻ���r��]<Ӭ�?�VW�/�Y;��I��s��� ֍�}v�,׼8��h*#
v�d�y����c=��Ro$�X+���C$� 2�s���ݞ@dSzֳ���Z�,��&�{�.�/�걻���(E�����/�#����U�)s�(�n�|C���ӭ�~#L������9g�f�7�lDn���Y.�Q�����\�8�/����Ͻ��Q�a W��P�E�J"iȍ@0�	V#H<���
O�M��'���[%y(�IS�N�A	Air:��S�O�E��E����{��:�<��'#�\�˚6�G��|{ެrt�+me�ie��:ʏ<�9=�^�tK\�u(>҆A@��g�[> &�W9w<-J��ˑ�<Wg���������e�����Z�7n�=~GC���(�4�u>Գ�֧
��bhd�6F~+`$.�T�ߪ���tԄnH]��z���TL&� mعS�T�<�}^ߕW:
�w�~�9t@{�6^%~僧�ն+הe�qZ?Vg�O�l�,,y(��.��®�0I*x�]�:��e���i5��{i��j̖�(��������!2v���[r�W�4u�	FI��оf��|�Q"�O��ѨӞՈ�����暮���x�q9��΋���dwձ8�c�D�qf�#;zG�2M�H���b(��$G�2"Uy?�ic�?�{�R�dZuw�q?A��z��~�������+�*�
ѧ����O�s���ʪ�T�f4����j�R�6��z����x���u�ͷw�-؋'m+mck���8�g'V��=O��uC2�+�)v|���Ww~u֜yD���bd݇3 �׺���9}��_��}���?��2�>1��i��C��\���/��F%}z�2���#N��ާr�aez�L�2���
Rhz��*%�FF�Ua#� ���1������m�����k���韷��������}��ad��_�U��������ګ�/ۓǏQ�Qҩ @��Q*!V0�m�CѤ�����s�r�) �����|�\^����#�T��ҹ|3�i�w�
��"P�/�eOj�c$ �	aN��)JN%��
0�O@X��?�!��Ҹ��A{�h�=����L���%f�Go���}'qkh���u�:�޸�xvJ������e8�1�����dqr��C�L��Qb�:Ck�-g]7��9���'G����j�h�d�sm���O<U�BY���f���&'����(�2�Q����|,-���C=m��]u�GM����Y��w߫.̣�#�b��׍?]��m����y��>w��^��n��>�pϯ�?=/�p}q��{���Ջ���������g�.$!"{�R���s|�p��})�������a*#�
�O����ȫl�̆[���*N/(��b�PuՔ]�/r�gv}���r!k+8%wA��^h�0��2�5pI��&�.����ӫvtt��l�ܻ���pW��0<A���7�(|�h����u�E1:�}���؉�����������.��TT�#~��<��}��y�Ng:�-R��*(*'^UX&t��4m�k&�W�,:?A)sZ�%r������;�T�YE5�˩G���2W������wi�e�y�	�m��J[��L�@�k	��@�!$��|;paA�`�MUu����{����{߈�)L��$�7N\w�1��cŅ�I'2���i k8g����:�2x1��w�H��Dj�������ס3��ed�\֫㍄d��Z���������ƤT]��y�) 鱓�y��W��e����}��7�������l��n�����V��<ehiǷ�Hܲz���=���b(t.���}9�%od��g�Ւ�KrA%Q4�{9�3~*_yX���6T>�W�fTHt�iV8�w��#'�VD%�\!�ϼI�^��� ���yX�IdXmX\�JZ�',{-V&MX?x��Q���\�o��lUI�q	�3���\�;�@<Ͻuϸ���?�Y��"6Rj`���Y�b��0+~ڍ%���r:LC�{a~>��4��,p���	��nln��Wg���ѡ�~
4���֔W������EN�U:�DuQ?�d��H9I���u�;qu�H����V�9tB��*h0�8R��i<7M֡r�����34��e�%�"��$=�������UN�GO둗�X�P6(��t}	�	m��"����|�㣞�_�Ym���!�5�O�Au��q���LЖ7���Lժ���湄��p�c�j�z��Pxי5/��r�X���#/#s�gu+��:U�?�����!�i�ުi�g* ��v«�Yy�1|s�a@�P&a�t��L4�\�{!D�WoW��u��IV&���8׾!�"�A�*��s�t{��I���M���h����ߵ��������q��_>k?�����ŝv��b���Θ�X�@�b�d�G\��'��@J��ɭ=)����\Na>����0���9���
�BB:2¢~_�H�8@`�z�/�Vp�݇�p��'0�`~�odf�S�\���!o�y@�G���;2����%h�T{�l+�s0&ad���UV#�59�ffڃw���<h?~�߹���0��f�"MQ]���n�Jlvf���ۈ��G��}4��w�ړvp�q��>���(�C`|��(�����0N����RV��F��*L7��2�@9����|ň�e;%=ǟ;�;+q�TqNw��99����>�*���ri�*<.N��A��>k�����s����6�㥢p���i���C�]R��]�~���V�C���+���A{9Xx@E���a�E��eg;ა�� ء�.�Wǐ��@;�~��o;qխ�6x/%�GC�Ar���u(ĉg�K��BS�Þ�ZX����;^ q(@Iy0�yg��X���u5�Ռ��@�B1/��A��|Ю��&<���E��.��
X�'��5^u���
�E]�tfX�	���iIJ�UH5jO-���gYu�]0�
޷�h� �}g%)��B),�<���{���8�g��:P��!cs�����j��)�?��^���2M�`�����bcKm®aM�����vzL����j�\���ӡ�up�6����=��O���s�����C%P%����<��)tq�r ��PD)�
]��@����:��RBH�k�J�[B���:�Ӈ��(���9
�]g���
�yg�Q�!N�a���	���0�T��uwoil��U������3���q�x61Z{����G�O>o����=��7��g��=��o�G�������΃_���?k�����mx�ĵ ��O�	�$���u8�9�3!?�M���� V�Ԅa`�|�1b��s7o��i�{�������{A $h�y�w]���	�&^�A�_z���9|��BR� �T���$@#<A[��(��&K���"�{j����|�������v崽~�>쌴���v��=NW{�ZuN�)?[�!�$u��5��r\�Sy�B��#��=@�c�YҰ�ظ��3Ϩ�o�T�]8��t��5�	�b]A.{�}��%8�ƸB��gXD#]+����M��}2��ck�'vp&	{;mg�:�%�u�Y�"��R��\���I;>�O�����`$��� �&����b�[��)x؜����i�8I}�@{�t�O���)w�N �3h	��P�rT���<F�"�yMͣKgy��Y>>m;����}��6'��a`0�p�N'isNL��̷���!� �R�q� ���y�?>l�G8�Gf�+�H�)>�;��5ȩ��Ӷ����^#`ңN������6<���<p��8_md��\u��w���,�ƁǶJ#7��W�K @��
�3'@�c�e�q{�����\����?u��������0��i����M��E�E�ـ�����z���ԁ�ҙWǪ?k~N݈�SCn�O�c��I����(;��?��zNy
C�<?�j{��@z]�q�����KK�Y`�լ�߽��{�՟��@ݻ��#���wnݚáZj��n��k��x�~�����}�>}�=y�wwﴻ˷���tW��'���U�2=���!d-�4���� ��s(m�x�G�����4��[=�?����z~~D�؁�%$M��_a�hΔ;�Adr���+@���`.a�M�ˈ�(-
p3�I�e-�iD� 'qb8���"^�g�������g����ǀQ�8����S�mkh��mQ����W�2�+�8:�Ʋ����!����zW%��]���#�H���tG��������
z	 �Qݞ*"�G���24� �ʪ絰�AŁ����\[z�z��z���v��r[�>00�^b���fk�ҏݟ:��I��i�o��0?���Ӵ���I��d
��$�l�kb	�SB[�\aʮ����V`�f����Y��ҩQ�h����A�����x�|Ւ�.�z P���`��ā�u����o7�T�JKh9�
2+��_�2
,K��L�o
?��=�G�ZI��u�!����<*��TC 9!��g�#=;��?�/J�bt�շֱh*��u�]>]�s�Ի;��e���/ׇ���G�#��.!ϸRHڳ�0�=��E1h`Vk'8��Q*1 Ho	���&��T�|�aKp9���`K���;;�mss��b���[ yˣZ��.r/2��Oeg�eγ\׻���Ơ�~�7�A;>�p�1�I�8(���5�x�@�M�ǹ��tP�:e�*_���q���䟕Ԓ��DKv�q�i�"o���:���.z��i�w��=z��T��f~���Ok�_pT��
w�a}�1�[�M�Y��5�N�ŧ
����z�#�;Ġ��P���[�ޣ�8Q���~����_�U��/����/����7�������~�7���_��?��~��ɋ�ڝ��م[m|j.KW:���U!�Ч2�X�o�6V_\SI��D����VB������^���!���{��!��/�w��������G����rd �} ^9q�Z�h�t�a�H��8^�81�}h��D`�-�c���8Y<#��G�1QwH�BV�U^�;� `&�Ua�	MY��,#I��qJ����e5��ty���tjbl/g扒Oɡ�r$�9(����â���>��H��R�G�PA�j�EƂP�ؖC�R-�XDF����=B�k��V3y����"�"��fB�A꺞��R��w�w�o�t���&�N,��b���3�H�f*T"C�gKfd����I���ʓ8���ԟ����|�.���6H+�Q[8�BZ�J���T��%��t8���;Maҕ�q���s�S��<�Y:%A�v�rV�]�r���7�}�s��^�qn��
��=�@>VG�`�����4�O��av�^��e��_�(r���1j�8�F�B�$�q3߽:[���vf����,�-��Gz)������9�G�'z���] 'ԑg~ם#�	EOۃeϕ[8�� <x��>�t������h��i�=z�u����������/>ν�Qݻ{/s��w�>�>}��J19�cx��LC
��̠G�����g7C��8u�3��GG��<1��4"�����:�$f��J��W�}�`M8Հ����{*ˡ�$��C�>|��Q{��y�;5%��Q&�(ȋvx`�f�(FE�`,W˦0(	�.�X�}��c�U��zTu�yX���������$��ȗ�����2$K���dUa.�c��"l���od�0��>��k��C��������<����햋=�TLO���FY��L��-������jY-e
'kvJ]Ύ+ZIƠ��o�p�3���T��S
ɖ!r �\�'Zl:%`���JG*ΉI'�S�)�p)gp��U�f�����i�<<�"n�h���&���-����v�J����v��\-��ete��d��W�4x&�0E�ǉ�%��/b'x�x�F��t��u��iՐx~ӥRѺ�@i�n�m�tpI ���e�S&�ٳ%4ND4�V(Bz��`Yg���J;�仟8x�g��ι'r��)����]�yh�R�F��4�Nw�;�K��AW9"j,�����ՊX�L5D�Bpqch�������ssj����9��1��H۝��7�c�����e��$�b4x=h��4��Å����&�T�h��( �E!���z^bĜ�5����D��CG���UƀW1��?9V���H(��pb�YGҔ>���V:������0�?)e��.�=C��e�I��ǣ��+ZjU5UdØ ��)gЄ�Сv��3�쉲�kʕl����h�?�Y����>��oڧ��M��g�^|�������g~֞����\?���ON�_�O������I�y{���v���v��Ӷt�Q�[��Q�؆'f��-ۓi���5��e�ȴ)�$�s����c�`��	{7����{��>��ts�ÁI8���ڣ`,������[G��4�����*�7�7p����ņ��+�����=hۄ��ch���9���d�6(׀��/i�/�Lx�nY9{A>o&��2z�Qm���Q�Y���.j���e��tu�Í�{�3:���6��1=i��&5$�����.$_��/�2�� ��*nI^�φg�l˷Vu=;�N؋+�Cɏ�t�*����
���Ȝ�w���(��O�joR�}+]k{g�}X��V>�o��>��e�Kw8�!�O'!���y�:?�8
{І#���/��S
�ڦs������מ��C��9��v[�I��i� ��ɂ]]�'��.u		�Y6�1p�l��qTŁ���	��^�;�p��0���8��ſ4~��z�cV�(��� ����*-C+�В�ΥV�v6�W��&�6���^%�t���������G�EhB|���=�-GB�F�B'�x}�|%��s�3/O'�H���*g���4�s?yv�=��z��I�_x��yή"�3�p� ����Ę�L�gOǩY�)����K����3�"��{n��L%�8�:h���P���p	����BQ�3�
�Ͽ����{�^H�Q�-��db�N<K+�#��3���XR�萹͒{4A�*L�����v���u�K9J��k̲�`�G �I�!
˫b������t����Dr��^vG߸�kc%��3�z�G]�:��2b��b\��� ��H9�h�H*ܩSW?�܏%6 TΦ_�M����,�p)�;w�ڭ���I���@��.��N���q���m���ެ)Ҙ��ɘk[�`|��*�
�έ����VZ?�w�3-�뜹"�Cƽ�d�ƴQ:q���4�u#�e����u�t�Tn-vikX���^F;��u��:�{��CY6h�V{�L�l��M# �]���s���v���z�8��:Y�T8TIo���(��s�m��E��מyם����k�*��F��L�tQjQR7���+b kbzͳP��'�#7����6�d��3��4+]���Q5�_��eטWY�YO�yV7����))ulS�w���=�O���K�f�K��NO��U��o��A�|�n�v�C���7�%l�����:W�k�%W��<,��0Ӷ�oc�u�Uo�)/�q�*���ƺ��L�2�Lkl�w�
q���c�yC��g*��`��87���Ň4J�w���*e%��t�)ܟuX��a��o�y��?}��zX6i��J�ցw�o�����"�]=NGKY4��\���߶:ga5�:i�x�N{�E�����?�e{���'���O��G���_'���6s�~�\��&�&x=�|���z�y�|�q�s�Y���E{���g��'�����O����mv�r�V���@��A�A�Q����ȴ+����gA"'��hi��{(�a���:\�^-�mP>h (�:���)��O7Qe�?�_���!R(��:�$�̴�{|zĽ�v�\mn�h��xJ{�%e����غoc_�*���6��)�O��x���x"�r�h�7)��J+��W�&N�Ʊ�vQ��K��W}��N�٥�ӱq�w�L'�?����˰$`�7�X�u��YW6y4q��2�V��4Tߺ��?~�1���vk��q2�AH�K�e����W�ѡl����<���Z6ʙ�P�ؒV���N���k����7o۫�or��X�҅��¡Va3��p���\���'d���D�;��xʴ�㣶���^�y�޼{��W:D�l�@�5�XJ�� �H��r�����CrʵMLe�d�(�����陛ã��;/�9��B�P���0N�Ζ�ؾӑ�n�H2�G�A��J١s`��)p=ҩ�q��+W]Qn�=@�@�|����'8[�k7�/֧>!�wҭ����g��A�� ����;i2#Ψ�
YM;�QUK݂RΫ��׳;��sa2�-*Ãq�$���[�Hs>~G��u�Ql����Gٜq��@���t�gW:V���}�`�`|�uA�ʡ�W�ǎ�0v�鵰\�'�.�QX8��� ;���z���U}�M'�H� ��_���T=S2���D���srl�Dux�1�'+�����Q�O�B�"���	R1�����CLf� ��AA�a}o��_��m�8R��O���#�r�
�*�z�y�%�BgJ�WKG�s�|��$
��<�86	
h�Q`t��"�/+�@x�ߠce�Ռs=0�2wy���_��:�Ѫ]ϯp`]�/�Iښ:�J9N���r�BC�Cp�m\?}4�{� ��
����B��8����!�wV�`%�{�ep%�n8��4�N�%L�̶��9��������V�������B!� ��O�Ϥ���+�7w�n�KsmG���q� ��E�J�H��=W�?,���DC!;O�\Il�T�u�wϺ8�~�\��ad�k[֊j��@Y�i��o�܏�u�9R΢L�]��z��Q����ו� $��n��bW���/G:�^�t���Q�n[Q��>&x>Gii���IG�\�"�E㜺%�Z�L8&(�����M��m�����k�SJ)�J�����O�4��'���,yTw�.��m��2/��VYE��!�r%H��B'���u���3�Qt*�h{�'mk{�mn�=�W�B�!b]�?u>\��J������Q ��vǀ.�����A��R}��P��6x�w��1�<����0t-�l������qc�:�3�,���Q{��q�>��_���"�N���64����<��Y:k��Xa�$h��l�Ghc�mtr�M�߉å����_����=��������ď�5�q��&)�鬻ܲ�'��.�QC���%
���w��Nw#��3K
��"� P�X)(L�ɣ�"�^#����_���<y������-4�F��&�+��8<:ù�o�[:X�m��^
O�<�O�Up=2de���֢��ơ�̃�����B��������z�4�6��gM'G���]|���r��I\dH�����Q\���F��z��K����(Z&)� ����P�d��!/eT9�B����#0�x��y�����'�|�>��q[X\D�a����G_�����������?<��|n���!W����E'F�t,W���ŹZo+V�C�`�V�uR��o�g��w�ő-i@���ex����m�2���X�����S��o�i_�m� u��N��l�g�N���{M�/�!�9�����L{ OC�lٓ�&e���<K�ױ=���{�
Mz����E���Ay�L{�\ �_y��Ƴ��N�:���~��q�i:�0����g������ !=�]}U!9����?���ix� r�Y�D�F]��]�4�!Yy� ��XV�~t:�+9ϸ��t�i��ż#��NȠ3ƙ�.;_��As�����������h�S鰰��MB�]�>x�3E@N�X%p�9����;0��:Z��q� ����e�O<��.��͒˶�:���k
/ c@�о���Rڶ��d�����T��#�[q��Yd�xU6*�{7 ��rh�F�٩�*{��{}JU�5�Ա�
@�NRr���]��Uޣ�J�Q�*����ϩ� ���wwx���C�0�_���3�����1��2�@��1��� \�t)�)�Om�X�+����ˑ#=�o�Nnt�+���fv��dG�Q�cO�p�}��t���אE�$�+���&��IUB⡟�M%8MY4�j&m�N�B����BD!c�	!e�
�ᠥ5F�5i��R���oedh0y�r�m-�i��C�ҋ�0[�Da������͝q����^R�C���g��E���
7����T�\Ĭt4��c�u�0�}�b����G������}h��8���c�q�j+�҅�z)d!ΰA#B���.���#���L���ypXN���e�.t�R쮼���'��	�ً�Ekj�+N^v�H�>�=������*'�Tj�2�.�W�<]iW9������B&����h�|�
�cH9��[ʛ���O�=W��y/�Ţ[�¿�u*���@ܾ�Xl'���\��V�?#q���u�8Z��J�P�BG�_8e�ڲ���!�n[��j[;;Q�
9�*��O�
���!����P P�yZ`|ůz��tNW`%�g��)Ƨ�H]j;+�O�j�����v��������ӏ�a��S4�t���,b����8?8�Y$i�����H��3�[�8���!����B��Yn��ڭ��������O?m����ݾ���q焐vM�/����`����{yvr܎���#\�G���ꃕ5�²B�����O>�S���o4��J@.zo9��'��߇5�] �57���9i;���.�ao�sR��UO�� �+��0nK6�rd�.�r��#U��yh%rP'+��D&��Ω^����Z+�e�����Iw�ۆ�r��r�>��ֲ2��j��2�C���O����S����4�x����-��Ȇa�춶7v�����F��۷ۃ���'Or��t[`�zu=�	�YeH�@x�N�`VHM���=�_c>�<�9����.�a�0��s����C�R�j���������m�0�m����)���j��i�N9q�����ۻ�wݨG8U���_>\�4z9���e��Ck�
�^��}�2�CХ��v:�pX��v��U�^�pϷڜ5�B]���rG���yaio�z�U�-����Ց|"ۺF�.h[��Fm�J�M�$M�_�<-p�J	�7�{����<���#�ꏀKXp��j�z�G�c�� �N��I�8�s��Y��ZMp6W/��s����{:��C���������7[pH�[�j]��׃"SV��F]�W�/��J��X�X�8\ [�3�#3��>=�!�i�����'Kh�׽��L)���>���ƯF�]������Ug�tf0�I�|aM��vw�۫W�ۗ_~���������mscE�.D���+�e>�b��Ԓ���O(T��u�'O��R�����P�^ؤ���y�s_���{���b��G�H7��;���r�H{?b� �Lh���t�Т4��I���+UB(P�� �ע�8����r�;�xL�U}0 ����$]D��ޓ��xԖ�ZhDf��5a+Q�jL�(F��� '˱��83؛eW�x�[���n�e��FY�J�u	|�%n��q�&�;�&-"0�93�"��b��
���L-\��0uE!M��\�����Ңc�q�L�=�lM�,�M%�3�e��.(��r�d)�s[z�B�J�'A�{�=��B����:���$R���}�U�c������+B�y�qVaG����a�`O��^��a�h� �,�#��RoWt,xO(g�b��
�Q<t}�������/�:�V]��Q�H�-ˠ����v�a
������u����q��1�(�Ű��"�f�i�b�����,�����t�R�3}W��@���$�b�U撓eXH�'cW�K�y�º���t�[�1�v��ِQƥ0�B�,<`W����0�p���N���^{��gK�F��{�A$�e���w�J���J�����G��
7��τ�:�F1/ʉ��q��o�
[���d��|���AsO1�+,�D=x�G���g���y�}�	r�t>C��ۈsE���+ͪ,�	�q�fV�3������0������CW}���k���]��p�|�"��ࣶx�N��vEUWaux\Ѷ�T90��M��P0w����6睬2��������	EcX��}��:*�� ~�������ݶ���6qvv]>�zuc�̫�;��9�i�M+�� �8�����P�~!�{�M�N�RG�D�!�>-Ya92�4�Oy�M�<�\��,=V����V{�f��}��޼]�~Yi/_�i++�����U���h���v2=�L�1}�I}�7}#�Ζz+e� ���ol��P�mo޼&�7����#c�ki����r���g���/ړ�O۽{S�C�)W�	t��q�L�˘2$׿��wAü����ƌ�D/#QН�"9�PHxd�5���F��d�(���-4��w��JGY�$6��V*���4�{�5��N��v=7����D��v�����u���3"����hts]�ƅh��:h8w6v�VH�rea�����h樗L3 ^�8��-�OIu"ӤK�SW���y괎�\�]��U�^��vU�K�v%��q5+\N^����FJ����-�U&ȯ��U5��%C|x�b �s�gҐ�MoV�k�W/g��ݧP;�:L6�i��o\���%_����9ҹ��a��6R��lO`�g;�#���Y�W������݇���w�I׆ϲU��m��NCav��������mmc�m��
�w��˰3�U =eq2��C���O �Z^n�d����޽~�v��B`2��#�8(���6"A?Ɛ���m���\����cz��x���G�a4�"�8s���I�V��r
d�/|���/�
t%F��4+�)�C�(��^�P6?:�b���.C���A_`�_�
�Q�b�_�
��lF���R���D;�� "���@��GGeXC@��A��T[�ٸ}k�=|p�}��^�sk�MO
s�g�Um�+��L�L�@ĜMGak>:¶L_8i����􊋬��)Q��a�S#�v�y�1Ht�)��p]�BZI��]�:M2�p�Z
*�%�ƨ��Pt'�C9\Pe�k��u*��t��⤟督B"$ͷ�C�K��,�P��:e+���
t	�j"BH�P{*̀�_{�B`"����q��Wu�C�����������s�3^'ʢ"0����>3I�`�tq���z�
��wHqB�.r[o�ֈuIfES`�ϣ?����h)D���um�3\�xydy��L�Ƈ�M��2��:=�꺧Q��W��%�,��A�	Փ�"��V>���CL-e @Ὲ��W�:���O�w:�1X�o-�%��j�Z������McRn�$iz)�ƹ�sa���k�+-g0�g):��pD���rx�����e���j��'�ɞ3Ȃ奥��?H�+#�H$F��x����H�}��˹
+)Y���@!w��yFG�ʧ�����ݶ6��z��`�]��#��@�� �%'��d�m�(6�-"��{�������v���md�<<E�p��6�_��xY�͇osV��kݧ:U��	}�g��Ael8|IC�	��֠�R���ʁJ[�m�x��oHe+�S.�C���p����ДU<�pP�/u�E�{�PA�P�?��'�>=����̄;��y��fNO����
��8o����8,;ms�mn�탋v�����p1��xS>���סVN �3�\g�O/������	w*dn��Y���;���h���V�Id��|N�$�� Ak�PC�	���Z���������|���t�����7uT?�@��2zOaO~e_��:G�_<��������")p������]����O���t���-�S	�����m� ���gmo�(�#�}i��9^��Ws����R��c��cy�>eo�B50��u~�]�1�4�s�L���66ۇkؔ{ѧ��j�	�\�p���|����-�l��8#g��CL��6;5֞=��~��O�l���PzvUʽ�ö����Wׁ�N�e`./��#���{J��Y�*�5��B����aʱ���1Y*��qÔyH'���:+��}Fz�O�9�W�;G�t:+�L�y�8q�͎.�^��Bd������$������F�+[0̆���Jx����(�eΑg)����%��l9�佰�7Mފ���/m��{�j(�t���w!�o���0=�>��kzH�Piw��q��������zz0�KU�my�m�*ZhKh����?J���<H{~�-�bDn��ˁN\��v�	t���mt�Bd�����6Ý��������8�|�+�I�)��ѿ/�\���db+�8ƻw�/'����|�-3��[-3�b
���ޮ������?���������믿jk�?#�������~f�
	��w!��Nm�,�F��)[�cy({�"�8�" ���ǵ���ϯ��DX�N���*�Z$�,@W�������Re#.0�8��"K��ppU�M%`�h���ݻ�p~1�t�`%ME~��i����J;�3�q�^�J�k��+�L:�z�0ѦfP�M��EBF�X1Rp�@=���5�|�{{�2ˠ�O�YY0-�t��<K�?���f���N�W'-"�����S:Z5�������!|���$���Sm~a�-.����1��(��6��/hT'M�ǨE����V6�����[p0�W�=�uU�#���Rp�w0��8�-JY�+gp��tz����v���r_,Q��n���>I7�A��>A^�Cn�b�'+��B٢ZV/,���C��S���[B)�|W���������^��}v�T�1 �p	�JO��k`gP_�=NֹN���*����ը`�e��������� 8d�o�y6�٧t�\�AS�EEF����� =i�#J&��C~�/9)��h��{K��CCi!���Fe|~�·�=!��N>r���
�⠽[y߾������/���:|�p٢�x��к���%M�0�A��0��]�]��Vz�Ne��YQ��aE���fl ���� +��K��r��x9V��
�Җ�޾s�=��Y{��s�c,:To�of�օs&�v��S8�p)��Uɹ�{���?hJ���wqx��1~��9�e�s��#��6��2F�8�q�إ��u�*v��'y�sEа���k[�8�[8��3�v�Jw�L*�Z~B�ऻ�s��:�yQ��D�nK6|���sW��+y������������������n#x/�Ygg�|tC4��sv��B,���fdC�����y-)NV�O�_\yg���Q�B��H�>{^������>y�,.Ա��C���h����_��������/_���|����<���(�O�-���k���ޣWgl�wq�r��eQ�Ir�����S�����`����ҽv|`�i�v����ԅ]^|�yZ�n�!?�s*k�S�ʹ{8y�p�.䩢?IFʁ3����YI�چe���9�1�f]|e�7���=�}�9�d��#l��l~�qj��HV:V��#eS�=�:3S������уmia}I�2K��9���y��N	���Ć:�8v.�i�I�[�8TW�o���:?=���S����'ޔ��|7���"~c�Xz��r�9�� �Iۅo�K�jN%�9���6�[N�5u���`��@]g�bz���2.���Qtx��n��.P8pW�xUW�vfF؄n;���Ց�R
�3��^B7�㙴�����Uc�k����6vh�O}g��M����2�iي��txۉ�N}�G�B����P�'�A��9!
Q��ƪa����~Ǖ3Ȋ����m��{���@:�y+���<��=�����)gr%���a�yd�7p�84J"
��s�������?��o���׿k_}�e���^6����m��
�My����,QYDV��ܸ6$�༯�E�R?��W��E�.���?���2�\�}�zF)��C�+�	�����r-A06���Tn��B�}z9D��. X��8Y8�� �t��VP(�L3�
N�D$
��.�~/+[��t�KWg��	{�df��Z?�!C
p�l%��ȗ( �"�+�:���~���Z#י�xPB��3�-�Y��P�&<����.]�vff��ty��P{��D˥�Ŷ��'kv�&Tf�`O[�)�uPq(<	��h�U��l��P�!X	/��EV���� ����w�:�N�.hb���&�'i�a�7�*��c:��u�3�/�.2�g>����[D�W�V'��z���� t?o�#U|T��K=��+���pp)q�N���?5L@������D�dx���$�����Z�.S�>jY���"؏q��3��e>@�����N>�/;���d!=����J�A�mi���f@I��&��	ig"t��m��qX���o��W:Yk�d9���P�!m�����/I�apP7|��[xb��f�#p�+uC�[OKf�΅9t��bYF��7���7䫼�Q��%t����-./�{���[�q��4yNP�1����a�n0��eÈu��u.�vu��;�����I�F!W��׽P�Tbtz��,�*G���w���|��f� ��7D�(C/��Y;Ĉ޳'uk+=|.U��ʣ�f�̻sw8�׏�����"�}��~�`Q�ԗ�Ds�����{��������a��B�m}��3:���W�(pȹ��)L�O�r�Vx�����,{J��O������d�e�m�����#���!�D�I�3\r5[)G���&�Ƿ�|�~��?�`}Ѿ��;�֎�\�Q9Z4`::]����D,��ԁ�s�k(���'�|o�N�/�/������n����z��M{��{����7o����J�H#�l٫���FC��շ�Wẻ"�T�H����78�,O�p���f{��u���o��������������#=>���N���K��p�����6����pG,��8biB;G�{��f��=���"v�+�)�T�G���#�焙�ϕ�:>:Z�A��G�����$n@�V��&x�9L�h�m�)�	2�q��!���|�C�пΓN����'Ƥ�x�q3""6 |��D��w
�+�N�-�Rxx�h���ز�\g&S:H�G��l�j����3֛���+�����{^���3]Z�@���Ȝ�W=V��W��(��K}����)c��ql`��Ķ�\�X97.Go�I׳2 u����U���[L�h���:\*�}f�E9b9�5Om�Qር���t��������kmu]����K�0n��z�p���vk$�\��i�q�{�W c;Nמ, Q̕anP�ڟ���&�wu,�޻� '�r�{"hS��ߏ`����2�0�9_�aE�T
fV�B��&P4<�c��h�쏴��!���o�^p�M4�8{�2��R@|^�!f	E%��B�(0#vqA`ȽP�����t4r5x�1�ҡ�0`;��
�#4�;o�J÷�7m�&��R�p�J6�3��A�
����4�߿۞|� ;f�^v	tҐ]�{�h߮�Cul����L[ZXD͑��uU/i9
��ؚjk�-)s<\%��O�O`��-S
K��y����L&x�M��+g)��VŠp�EH!�P�G�eR�-���U��`������g�+[V\8L�q�**{�fR7{G�3���.�8�SѮ�w�%rA��QO̒�g3T]R%Tʕ:QZw����4��)h�������t�4�A	L\�dTÂ0:�\.m;�'�cl�Ä�Ki	%`�axؖ0�8h��\���:c�p�����p���l+Ċ�U��%��de���"	`or�Yașt�d������Cf�6�)l3IY��u���OZ� J9���-�1���<�Z��)�����qJ�D��U��~�R��T=�|s*]]�������������=y�4�źI�s�֑Ao߾n�h���Lٍ�:�T�2P_�ZubC��<z�#�?8�(T8+s}Eyb��G08�������_#�6��. ��L/��YA�+5-,���E5�a<�K^��ᮡwG�
%K-�_�����N0��k��pC<4BΤSJ�zW�r�(�f;�ͭ%�Νۻ׶�޵��MʥA�l��ǟ|���}tr����>�|	��~�Q6~��E���H�C�ܖ�Ω����<�`���k�K�o�!��� �a@B���*��oҔ燑�"�3�.u70PfXu��4�g��:���ră�M|~i�Ol�u��Ĩ� ���3`l�,ҙ��RD�8d=�]`n<eg +�Y+�(�+p/�����@_.���P�n?��,evn�msc����՗_�����u�t蜫�8ӎ�����(��������!	�%�����U������9?1�x�>��"��f<����b�`�63��á!��Jo���n2;�&ы2�{0I�6~da��SWH<�K�H����)u��6(�O���Vu����Ω�|O�o�߳n�U��ߦ����9����6�޶�g����6N�����]y���vw]��lg'�2��w��c^=��5r���64>6�>���*6ر�����JZCo��Fp���k����8t�=�qg�e�߼}�66�IGZ�>� E_:7R�jJ#�[�}��T)s�|��F'��e�Z͵�唝���E�޿���7�h���q��G�����j��Y�����v���	��J&�O�j���<N���j�# ��%�ۀ�,s���o��gcsĄ���Z�=J���l�H�:�Y�ڤ��V'�Y�B�[}���3�]73�
��g�tx����G(/$Y{�6�@hbl�-�.�\�Pf�[Fm%�)[u��v-��\�b�M*�B}<�R\t�\䨆���Q��C�S�f�����RsQ�`Ք#����6�"��1iM>��K���X�S����Cg�Al�NtR,J�E�	�^����md����f��S{]��N[������t���<;�̃�H���Ν����G�ދ�
�jM� �Z1�甸{RJ�����*l����X�\�5lE�D=�º4���C��"Ȭ}υ�!�2���o�i����K�?�������O���]���W/q�j����X��V�)��]�������\�Rߺ�m�s���Q�����e�Q� i&��~=�d�Ʋ���}!!����}�����d	{iI��U�f��3��d�C�Ã�i~Q�J�DT%5�P`�oY��`DiW�zO�ޠ���$]�0n��@�����G\�3�lH
JCG>#A˙z[6`%�Kg:�*��ZD����Jie���"}�hOc�ɕ�$�hJW�̳�ґ��	��O\�]��m>�'K��;��b��ugqH����*�K�q��*i���ѯp�������������O�]��`��q Ntv��8��s,�%��{��&B�"��8����Lz��W
�si����Q�=��[j(P:xt���?y_)���B�Z��U�P��8~_�u�@�y����ɑa~/~<� H[{�(�j��p�JyD~p����[�Rɞ�Kk]���ay�H�n�}H� �x��Z�נ-�x9T�RΛ�(\4�|�V��p�3[�5,/1��0jߵ�߿�����D���HDyp>�S��F�j=�]�.T�;�C���)?hVe�|�h��$'��N��_,��u�e���M�ڝv�w�F��{c��DS�+�=�T�\��Sm��Ν�my�6�p.|��A5s�`����Qu���T����o>�9x��¼�ːOO;\�v[�}�-.��cT�Hg�)n�p�qB`*��p���`<:��u���M�°>=؉l�5k�-8�v����CWrٹ>����\2�`�=�G�&�w�S�>h�2�+���P��%6 �cؿ{׾�����7߷��޶6p�����	�謹_���E�X�@����X:�a��ʆ��i�5�9's��Ƹ��'giT��O�x��bi�c ������Or��"���3�ߚ��|�`�,�#5vˈ3M����P����K��R��=�^k#E&��e�Z��(7~�����,�L͠ӏ2l�[{���E��?�����}����N�&<��ʛ���Y�(;cT��o�d����`T
U�6P�����f{��m���W�͛x����	�r��lׅ'Rw�н<^y]/�v����ޒ��ʾs��\U�^YN<<Yt�Ӵ�n^�z�g~�U'۴�#l�vh$�<����f\�aMs��Ｏ�
��4:x�@)]�LI�<������/S��2p�68��!������}�:�`1�F��+l㭣�l0���h�C!#~�Wʑc�p�x�Uq#��Y�V��o�'��M��ˎ�~�C���9X�Oq��T���/���C�)st7�z��l'�N��O�Q��(��u�Z��w��ܩ?u��}Bt�<Y�8���p�މ�k�x���B������#���6� q:��J�N�?m�*����{���"�'�!]����	��^~���}��o۾AX�y�&=Y[����B�V�@
�Y��Ah�#uI�SU�������ֻ�:��������#ڰɄ<�c�d��Q��)g���C�R�\d�&jd���0̚[�\${ŕJ���p��h�8i�Rx$��_e��HE�$�9�w��Q�Ǡ�������q�#�k�ih��Yc��E���("H�/^�h(bHG��e����[&$�P��̐��"-��Q1�yuפ[�B��g��cۼ�P��&�<�'�!����s����]G�)��h�&S��a��ҷx���	�
[,a���:J�s�#��N�����V;9�h'G�ͺ>X����s�]�p�.g��4����K���3�q�@a�edh�<�@��Rr*���a�ԣr��on���:�;Z�3i�4g�U���j�8�lQ]`����zP���ꮥe��Wү�(ly�u�v��p����)<ڷ�E���I��O�\nK�K{Ewuo9��˥��1ם�O���92Sy	]�&�?�F�L5�$�(���>N��7���߿F~��B�5���fCD��{+�C��N�+����!MPw|���`!���^�E�s�f%`�N��[*<m���U��Wѳ�p{ӡq{1$]|��N��M�J���ёsN)���r{p�Q���!rp~v?��U��A���}]��C�ϊ����o�4����
�pO�����/��%���;��</G2��}����Y��{'�E_vq�Vޯ�7��}{��5��0���?� #%O�R�)u��H�F*�l�rk�����3�Ɋ��_4���d�u�����_;&'�;�qwo��nDw��o���h|����`�`���Gp��/�54u�4�MXZw��-�.4�09i��.4��u�KR����*�W�����yP�K�^FZ���Fz.�P����~�G�R
ኝ£�K[�,��l�6̨�]DA��3g����wp��7���#p�CV^��t�\�Z����{���u�mLq[�1��?��<���S���_��/g�FE9����l��_�Wg^������	�羦n�~x�3i��:����� ��
?�w�	˰����A&�c1��QIt��Q�zR+L�-�e���{^9
J��p9Oɧs���^OG���y��ڃ
�;�G�<!S�hbi�dEd�������ɱi�W��pm~ԕo���z�|f�Eͪi�ƅ�q���2�%�F�fuBj��m*�h�gY�ة#�kX�o� hI.�,Z�3��7=�y���G}ȳ.n�>���+q�����vYI[�RK������!����x
�vp4�a:q��p����8��%A��y|pT�){X�ԗ��A`�\����g;/ʂ��=��yb�X��9���
�'��
���2	���P�|h���Ծ�1Z���J���Ҵ66�+�"(v�q�p����aeź"Δ��%B#�%�T��!7q�p����	�t�	\r���o!�ϯ;,GW� ӖCB��ԕ�T���a�)QI���:F! W[-�������G�W%s�#{��LN�2�8R�#��%_�N�
�����|#uմ)�*X{92fZ�{f
%0�yz�M�٢���5t혚�4$Tz�ڔ��,muC�t�B
�fb��%��u��q��:7O�M�2��z��z�v��JO�A�|�l�[�[e�K[�	��B�B�<��<0�[����:��:�},�{u~�����Nvp�p���q�����*�C;:�Ǉp�V���Z;��<����V�	J8�oC���q ^O��'oPG��Ԟ
�` K���Ԑ��y���[���\4�����a�]�>+!,�����/+�zV�=�"W�wy�ùBX��uG������"xN%GO_��滔��+_��^wi[�Ez�'�ԟ��w���4��+�Q�,JX�h5@ŚCҎ�����n{�v5=Z++���I�ߌ;�z�r��x$mp���^f9����(��"X
�9Y�N�^��gZ�:�1���rw�tr����޷+o#�m��p2X~7)��GV�nqb^�F/`�>h>n��<@G!���h���#%�)[��]�(�W�:%��G�,o�b�o� �y�t��Xı�����};e���$�a������gը�p������������m������~����l�__�jk����#�������5�� >�����k!)�5��2������}���W_}�^�rV-r���s�i��,8��1�1"u��,O٠���2�(�mX��Kc_J�JO��#Я�J��PotB�_<���y��qG�k<r#�F'@G��U�"` �׭�d���E��'˅tġ�*g\�����Y��!hV���;4�"u訬|���~��[�n�{w�;�]�}>�G��}K��^I�HS�"��L��4-�שg��_*����6���Ѣn�#�g�k��l;12E��8��Vvi����n�����_{zuL��A���R>"ʿ�:9q�D=iȷDI��+����B':[�]9���cd��2_�(��*=�7�H['�z����6?2����!���tǰ�*m��Zcl|ǋ{/���:����V�-���1�L�S�9@�0�<�yՁ�\���w:�_��}$�o�� oz��@�0.��. l�X�;z����>��P�\�!ny�=S&�����QR�;Φ��^g8_7�J��t��b�������9x��GWF���}��_N]�^�kQPN�#[�-�$���<*g>*G+�ԙ�s�d(*:�+4��T�̌'
3�}/�zc�����{�auβ�M���=2�3�Y��yC"�ɽ� M:WTxQ �P�4�He�����'R�!��~U�A��ﻪ�������d?�������`��we ���Qy�4��03ugOߋ�����/jrBT�0f:V��ս�"	��gl�á\E��F���ĥ�)�����Y�*�f$nz<?;�q�.#?7�Q�-���:��0��uQ���D�'��[T
nHWg?�,:''��#4k��$5y��g�(�_�y�������I�N�`o�$�蕺�`���rT�-z"��B�r��M��R��y��8����-�)"��c�+��8�ʹ)'�8L��:�_8W�{�9W8>x�q���Ώ��f�]��L�mq&�n��g���7qරޭ�6�F�����ɜsۗ��}O�U3���E����η]Nƿ��@��C�I��}=��^��X�P^6bR��7�']�P�W�F/�P��?�ڲ*#���6T�l:����x��hr���c�7(��G�0�z^y��i�
��#q�˩��5��m����ﰓ�h��E��J�8�D9122	G��+����
F�붶���?a�+y���(`��������zGK^��k
eM�8�$���uD)^��KO��+�y:����9(��A�����𪭯�����$ƨ{ߌ -�ɑxrSR�'���65�Ԗ�w�;w���%���e.�Ԟ樳�
�|�Q���G��-ӯ<���{�a^��͞�9�0{M���4v9�_���ҍŒ�T?��<'�mo�e�]�ﻶ��m��m�����sW�E�_�B� 2$��B86|���1��I����Sޝ;�� ]��)����y�W����[���h��ǯ�h��w��K�k߇�r�Nw��Ip3����;"X���w�� �q�ڃ���R+�]���8eVQQ<�!o�B�D�W+à�m�~S���ߒ�^�L�鹜��A�;��o�%�y(��߫'��Zg�T�.iB�νqnϽ{wۣGڭ�˙���a�6�*��q���*�6����r���{ۋ���>�Y��ŧ���ѳ�����I��^�j/�r����l�#��7�����ޜp�ԭ��pݿ���|gp�|�cy�m]E3��x*C�.ۍBBs���3�a8G���c`�0Z�)����9q+d�d�`����>������vpd+�H汏�� �u��/s�)_�y�o�T��P�;�о�i���v�9G�e+�M5V[�䷰��q'؅M��l���� 9�9�#ҧ��n �Y�@zRo��`��8Y��[<&�ؘL���eϿ{�j��,��(]�橍���D�c�b�p� �6З�E��8��Y:�n}T�.�2i���;:�s$���{�c����_}�V���%c��>-��k�e�Y�];i7��?�GW����kw#&���2p�e/��'txWZٌ���(~�a6L� ��R�0�e���2:��/x�M�w��~�+-�Ad����U��xR�+���c�u\T����5�Ɋ\��F@��B�"����C�����aV UΆ��yoR!��>>\'sሴ��4t}��*O��*���HE�3U�GbtN���-., XGLN$H���O��Vg��p
���m��?tB�=^G�Pg����0%��A�Y�8	~�ɲK'kQ'ka�-p�f�*�͕�1��iv��S�:Qxx���x�X��ɵa�=簌}��5tۃT܈�~�]�4�:��9�|H�<�g�V�2�{fgZ�"Ԩ��Li`Z>��Q�^~��$��|���)����(r�X�+�o���-��v���c���֎9�����v��t~R�Vg8L�8L���=�F�܅޶�m�n�uE,��V�?��JO���Q��o��ǘ.���q���CZ����#�'�#ɳte��xTZқ�~(�ڛ�r��Pq��,ՈRJ"2�P9��ru��r�&�Kw����Y:V[ۮdZ{p�^�L%iϖ�Wr���{���G�5�}O�QX�G'��VY��Y�zOz�� M�b��u.��8V�p�ɴ���,�9j��;ʍ�����J���o9�k�;��9�B���|�r����*�4%Ot���U��?��=�C(x�C,iI�V�^2����C��𲭼���U;:�n�����r�%�
�lp��u���P���e���֭mn�v�@������<Ja˙2�L	ҡ��5���q���O�;� �>T�R&dK�0����ΕM����aWh��­�QRtl1�k���j���w�1(�}�޾�&�[v�[���r��y�N���;2'C����:�� �-�7*G!��}�^0�N�?>:�g֠�W��n_~霠������������I8s��qd�χ0T�E�$�XW�o��+Cyg�#-�s�y¼(�d7�\�u�[��������
����c�!�Ž|8�竡�w��}�	�+:5l0��Q^�v9uĈ3��}�s��]#>��|>��8��ɓ'��GeO;�^	�2z�9����ޞ�3�q����=�Ct�����ً�駟��?�Y{������ö�T���>XZ����K}���	����6��m]JO|K_G���!�gQ��d�W��(�t��_���ƨ��ߓZ���v����)��'�g:V�Q�N9�q���sD'q���4$�샻��-�M�;m}!���$m9�P�2/��Ɩ�lK�$9����ؤ�h'�N�6@"�v��Dx�]r
G>�V̨�4�Is��z�����᪈60�{!���<K���X�	oy@�Я:�&�G�|�uJO�~�Nᡲ:B�����O#��(��g��4|�c�уeOE�tw�Ly����U�9�ynv�_�!_�n��ًm��n���9�Ps0��� �ܤW4�T.;P��.��>��*[W��H�9�J�^��X���!,�F�Oxh�ʣi��Z�!�t��LX����A$��U�2�L��A��>�;�����J��$�J��|�Xr�#'`J�
�!0kr2D �m=R8I�{5\�bk��J�^�PG��Y���q������ �y��Գ�<�e����g���7�t� '�� H���#Fu���s����p��(�ސVv��̶��		�C�qt��W�sN�D/q
7�̸����\�e~s*�)O�,�pV�s��!j����^��řvky����8Z3c*l{�Pz8Xq�\a'�?ʘ92�N���*�!���;_
�2�8�k*�t�Qz�`�\��0!4�OFpPx1���<5��m9W�'��L	+H[qxC!Y�RJ��Y�/��F�Үg�Q��H7TP'K�ͪ�]��,�v2��,=YN1>}v~�,q��;tq�϶S��1�9<�������^8�k�k�y[8i:j	����"(p��p�	�z�!4�;+Qx(�����t�:>!��rid_ʧūy�蕐�4��2wp�vw�14t�Tf:�%g��:�
>��-�̙��IxO�<S/ޛ��2�>�!G�$���4��+��$$������C#�]��e�4݂�u]����)��ߞKׄ>�@f���N��a�#U���NCn��+���o3?�����
��^�z�)��o��(u�q�ïy���� ����S�։���aBUy�!��ڄ�Ӹ�I>׉�7���l�w�j�}���������Qe�@n�sn]!̤������R[Z��u'�;ohXY����̐AR�H�4�W�t��	�]w�3�Ы|Ч���}�_s��<��,�H̵��}�8��iH��*�Ց{T���r��p�-���U�x�V	k���ƻr��g���="s�@M�4�)Y.���(����M��ޕM�p�]('s8y��fW`;<�M���Wo��_}۾������oڻ�k�C��!��h��z�r�v�
���=��/��c�s�KG=�ˏ�E�V�f�Z��P��_l]F�ِ� ���o6M��r�^����y�\�Up�RVp���5ܾx�z�;|��8I�}O�?���Ϟ?k�|�1��g��>�9z��ݻ��=�%MxT}JF8��>.KG���:����X�]De�N�s�nV(\^^�q�zQ�}�G9U2GY�<)������q�"���8a9~���)/��K�
�[�T|d����{��P�j�;M��#���R�g�<��g��ئQ�|u�������+��HP�@��g6�J��+[�4/� �F9l0���v�}B��l��a�8���[�HA8?�y�ɂ����=;�y�V=��m��OP��s���99�l<��׆�g�F7�w���~;8tz���#���1Z��,���� �ЙM/�M�.���j�l�6�ý�i��='��,����;J��N��j��6�qZ��ҩZ�ϋ�i H�~y���k:��8Y�O)�|Q�4(����k�,W�We#�q ��y^g���:����p��ѽ��L�Q�R:}̏�#���w���F[ݰ��X �r�e@�ۍ0E�=%zڢ�Ve'%+��H2��-V��X�0�D��ي*���`�\lm����1�H��y[{�|���Ǚd��y@�5ԡ���z	�5xG�!�.���ݵ�m�О�7΋{sT/��lzւd�崬Fp9��-V�|)GbhD��~�%�� ���me;?ߥnss�C9S*
&o��5D�r�w:��n�裇���%�Dn�m=:h{����=c�U�8�2�x�����C�J�����h�:�cu�!�|�a7w�dck���据rh+�Kr^1�FCm�2�J^*xp��ȼ��@	I�K�2�x�Ϗ
����QIN�h`.��?���A�aL�3ʮ�eV�3w��-?���m�M��M���+-iz�}���4�w��C0�bR�(�dUdt�O|N�I�V�!79�%Y#��άxlp�@���8Z��.G{�c��D�!����=.������#��Ә2�*���7�!Z:���(��k��%��^,
m*T��}����g¦��-�Uk��C�q��D�"@�kҌ��h9ֆm%����0202�9:#1�ɵ����oJ  ��IDAT�x��x��s�|��㚼ő2�C��e�5�5tf����{����>k�+�V���j���F����.{�c�<U�H}�i��.9|%�H�W]4 '^��~��G�L��F9j�#G�5�>*I`���=~�j������o�����O�4	�zG��G���!��Pq�[����|k��ux«}������/��7_���U�?��8P.�c����*�-�iń�����?��-,���4�D��tޅN�4]zAZ$��i�o=��u��������'G#X�f��+t�'����6:u�ԙq�����:�fx�����y^�S�M��lAGz�'r�+G���F�F�G:C1��S�Г�g�|�\x���pv��vrb��a�qks#<�������/����+�N��q�Y�¡_���ad��{���d��Kי|!b�ԯ��L)c����>=MA�T��L�g��8�Ր&?�8=���}����s���^NIW�O^�����S�Ka�����ؕ��H���yZ7���F�}k�=F?������������t���f)kt��ѫ:�ƛ������j0��|��NV�otQ��A/��j���T�"N2�(0�QSʫ����"9jϔ�䰾�n��;���N�{0�
g�G���(���5��et��w��<Kdx���w��:�(�W�����*M_:dT�=k3Sc�u�=zx�kz���:iۇ������z��ܡ��1�rJ��)sޗ���]�|!�I�668Gԩ�}�7/��T�A�������#n�VK/�������v�9���Vm�#>+��ҙ<���q�)ɀ P8�Z�Y �V��i�+4*��]|{��'O��/u$�>mP��_�s���mܨ<�a2�p�?p�������ݺ��Wuzj:=�.�'Mڨ�=L�O��:WY  @߿��N��r��н�6������L��\��S�����w�]�?uXG���	�cx�tB{F��761Ӧf�+S��kS��a������9�������_���}������rLaA��ak]�5����x���H����vۤ���(l��0�K�T��-lω�~��!�8`�/�8#1ޗ�z�`}��GN:
0�� F�A'�"�����UC�D���޶w���8J'Ow8U@)6��Խ��ꄎ��0L(ZBC�/D�
2�N��!"C�y�PꝬ=� f��TV*��KVǲ�BÈ8��9�aiq�ݿw�=����C�*J�߹V��m�8P*)�aK
X��bg�d�`u�L(S�:�G�"!��R1>٦�I����o+�8v�r�4��ӄ�ʹ:%�aX�9Y�)��O�C8�]2w��&��2Re	T�Q��\���=?M��DK
�ͷ���v�E�t����P+|� VY
FF{'�#.{� ��[�d���&Ť
'a
d�Q�N<�I���R�c'K��I/��RO}4��%,��Z��ڐ��ȸ	�'��}u�c
4P�Z� E�	��DfL؄��*mf���:�M�������������9`(�Սw ��d	lt��R%�tk(�b�P�=�� ��iԆ������x
Ho�����o� n<�\���*�\vxiy9y:�G����z��}[_[Ok���!X<O��9��vC/�M^�������gF�s�v4g�Ut�l1����:��P+;���BW~��qzeg���|�P+� ��JQr�pN0B�z���_Ή� 4�8�`��6��s9���`'�=0��}���`mn�������J��A��|MK�g�J�3�S�np��i.{��s���$|�d�д �����:̹��q���:����9��yZ/8�d�U~6�Uy��%`�
m�T�������.&p8&���c�k Kw'-NVV�����U9{sܠ١J�s���}�(�E��x*|�� d�>����p�V��~��o�7ν��M{��C[��j��F+�`�L9���Z�,,���IqA��h u��Ј�?�{���4��=׼ŧ�.b�I�K�&�|S��w��o�i�v�_5�Om���\�&N�J��ؚ�8z��ni�%���	�������>����W?o�xў|��=��޹��ՙ�aZ4'�e����V������h�r<\��F����{=��y���{4�.C&�[�@�V�lσ�4I�5,/+'��xBҐ�z~�0ۆ���K�.��R��������=�g:YPq�o��r?��(rz8�^�w���K���)��$v�{ �_���d�\�.��eOq������j�G���CU���+xxޡ��i�O�Xy�
���Q�w�gj!P�#�Qv�z�x���c���=�}}=Θ��z����KHCG(���OX��A�ǻީ2]���g��rD#�rF#�W5>P��m�䟆Hu9���*]�KWMvOčߧq�wi�vUGq��d��ͦ����[�����e��Fԁ��m�����p]kcE�QW�/��i����c��x�,'��_G��b�����t*~�[�M��N�YA���>��5]N�����?p����봜��ǿ��w6���^��uVV
@��;���p<�C���ڱ��8Y�TT��_J`-�c ��b�a�_D�.�!� :UD+�éᾀ�so�1����'�r�{�6��ç1()Ii�	[
7W���+�K,��p�d�p��s�i�B9YԊ�������G�!p�9e�JE��x��F8���>�|q��eKBY�1F 9Kh:ZD�`��;ZA��	�
�E�ͻw@��-�m����i�,��!0�������pu�8�&Ƣ�8����°�FeIM
����([�&Ł�7N���p�ys ��F�i Z�Q���:'KF�o?V���C��r��~S=^*;��7�-N�J�g>���p
S8�K��/W��ɗ�U��V��gm����3�,�U/=b�'aP q2�9YY��Շ���4�w��0�sq�gֻ��Y���"X�8Y�Öc�\�9��s�N�Sq�xqj`
Eh��;8�vH:��u��_`'�34�Q!�l�wZH�҃e=0J�
�3T)����]�������H���T&����I+��J�Q8�=Y:����9^+{̀�"{Sc�?i�ѸDad�Q���UHʉɻ�?� #�����(�۷o#4oG�oY����P�ݹ�~~'�uK����}�K��x�s�>��W׾�?��+N��-��s�#�'K>���)H>B�+'�!�!��Qz=T��n&����K��0�-�sB-��|��*�1&�r����������=��'�\��:�M[y�2�ߣS�S�C��6�L�A��C՛��3ʾ�e�,��Y\Xj��ϐ;�F�f�Lz�Έk�1<4����@w�a����ß>:H�����*�I��JNX'J'��Υ�������j;�߅�1y7�L���FIi�5>3��t*t�ML�����$��!��3�k�w��1��iM���!h$�-��Ycc��.��\ta�m���_i�߼n�~�m�h��˯q�ނ�u�B�#*kNI�xj��"�R'�,����f�u0��z߫l���D���8<+����$���CgBY�ɢ�����!��\=�4��>���;Ӄޫ����t�4�6�e��J��`�<�7�Y�������_����?o=z8h�� ����k���9�����a��{�.K��p��G��t����@�6�P5��wLbK-,d薺��d���[o�9p���&�8Y<Ϫ���9L.�!�i [��i����-�S�
g���:M��g�Ţ�՘��c�k��4(Djp�%p�N[�a|W��h��q`��ٚɪ��E[�{g�N֛w�mm}+���м�R>���h8d�F!yPRɦ���a�'ǐ��w�k����W?]��@:WSĝ��x�V�?9�?k�!yDOQw��a~s���2����gp��}śN���x��u���Z�!��B��4��dQ$��<��-_?L[~�:�xS�*�\��s�R٤\>:X=_ȋ�L=�^�栵yh�!���o�g���\�B�����Ӽ/�$�ki܎���Z�Ş,������6��)8�&�Y�I�ҩ�H�'�A�^C�u��G��8Y�}O�Ll�8Y8�:Y�-'����������+8Y�ܵ7��Fh�C}�z�n�.ځs#� w!P�ƀ42Go�	|Y���{���  y<=�ё�6��w�~��Y{��E{��i{����죏�f��ťe�	�]ʘ�Fh}��Z��l�N�>U����޽h[��mg�����W�N��p*e<��J�Zs��8w]�~!�C�3��� ���pu�b@۲�0�3�F��/1�5����+y�8D(���1YK6;�%Fƃ��.r����R�$,,�'���h�q�vQ��da��TT,�2BZe��f� q��?TZ5R�ԯz:�n�x[��� gfl-��� ���n�ZRNd�6#��aq��h&�Faߛb��{�B�D�!���ٲ�=����zT뭂�R���s?�鉙6;�H�б	�O�4s�p�q����w�z����B,F��Ȗ*�{���-.:[�_R>R��X�����)=�^#��T��q��u���rueO�.4��N�\��[ma��X��]]A�W�ouL�p�I��<@�<.�
����J�h�y
�iDq�Y#?�V�����rh�'�r���18�!�ĳ�9��JK�L��u/��B*-��xVA�1�R#qlL%b��s�e��Fa�pD� ��^�K_t4蝓��?�	W�!�s��e�!+��<�h���0�8LM�"���ގ��U��g�8�z�?1.Hϐ\��4����ɹ��^�� 8���A�8�|}N�2TH<ȩ�h��C~��H�m��%�mlĉד�3��l�u�X[w����˫&��)���.���/g�+�cRI��`�p��adBV�A{�Zm[������mm延��m�Z_�q�C����%_�Dc�2:�a�C�Sm�v�����C<�s<�2�f�i��&]
�>�_f���t��&�|Y/��x3t���w�����i�Ġ���Q�!ƹr��w�����x�����QA��d9�r��cp��ΰ+��@�.p�jc~#Ϻ��ҍK�A��<W���:�$�#cW�=��=�o����w��������m��B��v��ޔ�������޼{�޾[i/_}�޼y�c���c?ll���vr>�N�����pC��m���	�%�qd9�=P�vA��t��a��܆��Jn�Cq�~?�Ɓ����{�"����%�E��k����1�N�N�[�wi�h��k��9�#��IK	}�	�<��C��c{:��j"���ϕE��y����'����/ۯ	��x��<Iz��!N�B��Ҏ�#Oy���!����X�~6({J���4�S���;gԢ[��S��:��]W���v��6���vq�׷��p�& �	d{�b�# ���^.[�9�#U��A766���`c��|����>RV�+�T��9�Q=؀#�ހ�L�;�jq����!��(�Q����H{|�����ὥ��8�&�ؼm}� �����+msm��R�	����ʹG~��a�"Oű�t
-] ����'�ۯ~�i���g�S£��1���V������jS��<�i�?y�~���ǟ>nϞ>hO�?lϞ?j=v�H�r�R/l����g�?��>��t�}����1������8_3��������	|z�}�p?ʛ�[М�]���+�3���'����6��:X6ꄮ�O�A�Z���S6���l��gB���P�0����V�C\�biѽ�n�9�2��(y���c)��C檟P��p��r*�ΕN��Ѩ�2dpg[m�g.�Q�U��6�E�^<��3���qTV�K�����~Iv�&�	f��,�
liQǙ�H;>�#ש�����C��5���]�r����	��FeJ0L�w�T��`9�
� Q��~�4�?p�x�R�����wB�C��0ć���"]�����g��>����ٳ�[���8z� �`8�b��1H�iĖ��p�*G����U�۷�'�쫬��ep�^`G�h���'����Np�� ���Ǌj��ƴ��΂
5���c���2u��7u���.���w�0����!�r�8Y������&F`�r�-Ň�mwBu5"�*��-��_��z(�e$���9/UW[�h��#�e�'0�2|���A����E�b�R?�
��F�� FY�٠Ů=EO|E���DeL[t\�ұ�NL�gU���tg�Ҥ�Tu�%��O�J<�3��#�0���u��mcHom���q;t�-H��j�K(
�`H��a��p�T`X�)���,�)��N�UZI�⑜BL��3��B��w��loVmD�y�;����[A�\�q��Q`���>8 q&H*�*l�G5B�p�F\yɠ�^(yY6�G�g��.���5�,P�T�J��{))���w Ö�����퉎F��P�'��%�Z�L��[��e�����l���Rϡ��$�2Kެހ�����������{j~jk�Ʃ�}gg���k=���z[��Z�Ar�p]���8}�k��-G��s�u��e臗�,���<����*�����Q�	���S��N0mp�WӲ�!�������a�7�+e��~��c����<�s�����C��mm�b a�c<�"��n���
MH���뤤����[w۝�8�n�x�ո	JTe�<����R��N����O�����s.|�.=�U���`h}��:B�>�����l���x?�l��K��T+�ymZ�4y��[܉{����3GÞ�cx'��\�˹Շ�X�N��tx��쿵���C�1��67���ʇ,p���a�j�!<n�1=��S�������N�)����� ʫ~�e�����t��,�`��o���� fIO�5��}�|3N�8�McP��p࣢^k䥬���T��o�����,+?��?q������ �Vz�����ϟ���9��sx�|o�]���߳U^��͛7qd߾y�a�>�f)�3��t��p8�����:�p.5��E��'kjz�m�l`�}hG'89�0�'�^,i,0�`"5����.��e�3ؓ��%n�l�G\�	�ޱ�.I*�����T&	[m��#���Au�=7x�i�©X��l�����W���w�2�X�Hb˾���>6�姽�Br�ܹN��u�����ڰ\�q����\����/�_�~����Ƀ���=l�[8u��������ѣ�8HOc��c���O�p���&��<DF�nK8g�:��ړǏ��Ϟ���q��/��O�\=~�Q{̻k��9Wtn*�{K�(�kH���.h�C٬3��2l� 0|dP?Js�:�:X��9���>����xօ܈7��+�$���:|�ӳe���a���@���h�g{��@��?�kuS|�qޮ���p��&�@�EW��xD����o~�w��\�|��S��S [���q�$��rE���36�a��d�n�\���kO̶���ayr���@ø�1.U� U�t�F�����R8_�=F]Q(+!�c��P���/�е�B�n���`	O�<n�F��_�`��s�Y���1֎��Ę��T��`�dMb(���f)�ʆZG����:Y8X�����B�d���;Y������NV��#�QuX��(!����:8�N�=
5\Pӧ/DUF*b�ƯP�Q^ꩣj��F����8[��ԛt]�����-��L�sC���	����$)��_�YR��~�Q�X*�!�ُ�v���w�~q�:G.C�٪/��d�~o,	!��̕"Lʘ:Y�O��kYe���`9���s4���⪘�V˞�i���T��FX�;MO�(�-�
潽������ǰ�E`T>:Y�jÁ���v� sr�2��]S�X^�IW����ɂ��Ѯph���%�2��x��yW���.N�6�}�I�{�OC�QH	��>b�R���DA�VϮ%VERC�zB7�e����霬�y� ��9�RV g�'פ�� 6Sw.�]�����75��~//I���u��+��]lh���CWf[��o�(
Ex��E|�uN�QW�Y���PI�K��q"��;�������G����J�ʾ�}'޺����bե�T��O>�K:>��r`�¥B��<K:���R�ʪ�ǹ��1m_�qol�@��+�'q/����qz<PL��搡3�!�!nF����(Vs&��[�'��=�ФO��[�	��P~���{��������m������h�X�ޘ����4Y�Ӭ���s�����|[�}��",��aA�H�,-m#��3:��+"l:��?�����ßq$�DB�R��{��R�.L;�<�ɒ��p��ww�۫����a����rɞ(l}��w<�U9��3�+�38r@T�Y8:�!�6����wb/r62�������N[]]��:&�t���.�	G'+C�ϥOe�21`'t��GV���ٍ�����y�����X'�d�����C���8�:�!bWO��F�rJ+�C��*f�Zh:����7#qdH��a���8����)G�T��ԁ��^��s>����7�Wi4vH��t��[y����"F"���C�8��ݻ�8	8�����񩎖Ԅ��M����	�d�Wy��oe��[����n�7C�����d�^l���_���0���hz����]	ZY����/읊ܰq�F��O�����<υw�� �k���9��	ŔyL����J�8:e���{�گ~�i����y�sk.��\�.�^�2�lXb�RG*A^��pޖqvn.�R&M�S�#��;�׿����/����v떍ٳml	GɅ�t�޿�S��=�az�S������2�^�����p@â�/��|�o��L=��}��q��/�n����s�@�A��/9��֭%좑��c�~ãvVs��ʌc8��9cna�T���;G���=��M��Ɓ�7���AX��ޥ����^�^�2=.����R[��֡�N�й:����
��ۙ�X[ذ���W����|�Z��=>S.�EN�om6��<��/	�P���	-�����\��>Lalr���/g	�~�/��[]O���X=�����o?p�N�HBe�ɩ$�:�oo��?Ĺ��ىBHK���01P�^F��4�5z��XS������1����/�����_گ��D�f�K��J#�$�e�G�V"�im�vn��A�È��";�l�ty|:L>�(�s�g8��dEl���G����c'��Ǡ@ݙ�����d��ʐ���ɪ��h�E�\����kY����OA�1�<#�,87m~��k�A	��´���W�d�̩���'�T�d�[�Xjt¼�$�e�.�c����PX
#�(#�\�:
c�@U��%��uR�q9R�e�*�{�Gb�+��.��?y4�{'˕�4~ŋ����8D¥��Q�ek��S�6�(�)����+����#��Pt�1�
D�I��d�)pq�f�,��J�"�O,
qY��!@EO�1��f�1>�����L�#�h��9Yv��Hd1
!M⼓fᱜ�~8�G	Y�قCc�*�� A؅������>U/�A���F5<�O�Ϻ4�5V�9s����SO�#�A��ٴu��������¿����u+~�F�w�h�#�:�8H��Y�� |�3C&x�|���=l�I��q?�I#M�1�?9\P��19,cU4�ʣ��iǀ0���郇,�{��!x�/��Flpn����^p�}'��)�����;&Br���R��y/�ИF����c�JPe×`�����'�Zyf/��w�O����s��G{;� ���s���m|x��?�m�8Z�x�[�CPT(�ʻ�V��t������E�,�e���"N�ݶd�/V3���̳���6�^C7�N#��y���zH�ٟ<�pW�Õ�b��/�)�AI��T�����z�E&�_��0���/?�m��`��7=�; x��wDB��<l�p��sh��������У%��#���5x���9Bm�uc���#3��B^�@�bC��Ut�*;B�\���^� ��lҬ����m�\�s���ܧ�2�u�_���K��#�.�	t��a���&`�#a������"2Fi�T�,ō:�<ß1P����vy�����%��g)����T7���o���1�gf�M��y%-T��	�3WO�J��8��bhj`jlʋ��C���u���ij��^(p��^�#L㪼Zu���Ł�����_�,o�[h �hs8z�_�I��N���T��������I� ��G�:��N�<��_�:�� 0̼`�	#0�����57�FuS�v����{�#�W��8Ys6�kH��U�0��������	��N�L8�"/�7�vN�zGmfj4C��!��ϟ�p�w�#���IW��6�L/��[˱_u���u��e�������ӡ��Q�ns��䨣;w�q����ot����2���42����&q�n������|�.]���D�X�0.ٯ�V�QM�(b{��6�	wG�8]G���V�rԌ��������+/���%_|�m'&��^�ǥ��A�A�J��X92����j��ͭ�̷��\�R�^��t3@��W�$�SuV�Q��bٺvGx�'�ѻ7ޫ�st'�>15��u+.��=�;sڝ۷���N�x��_���}������X=Y*#7	tn����/8�B�[�����p�L*�` nf�y�� [Aj���t��(�V��������7��w�}�z�I=��e��� 1��r�����S #cz�,iw�W�謜,{�vq�����s�d�����A������ԇ��a���GQ�䦐����O2+'Kq�de��9L�RQ ���\h(�� �m*bE�35O�,8A|�О����;G�*#��:�]�b�L'K��AꜪ�:�m��@���v2h��D��`Ӏ��S�g�ShH;e�*VLP��4����8Fi�|'�&N��|.�d��a���|/q�����A[-�vU�,����1���(rT����밭�m�-��C�GF��:Y�7����3���S '��:��\ F��!	B�n� ���,~��ؼ������n�	:=�ɢ�Y���j4[�({B��R�l&�� =4���Ç���Fm	
�2�W`#��`�0J�S�5���K�ץqH�uo]}ZGw�Wtp@o��!]�EE����qa�s�^�s����^�(���ԫ��4�����e�Iޢ�9�7��IߖA��4Y�R?{�����r�CLG�A�0���v�X_[E��du���4m}R7{��I��J;�?�p��WY�@�p�]��AX� s�(ɳ��B�.)F�d5�pMԴ:��°�n�����̫�q�w�������ƘF`N�!���H�S����61ڶ8UV��Ԧ���[�˹��x�v6��}���z�� /�����(>^�UU-e��tLP���N�Ƈ��5l�z/�0�-;�W�9�0-������+!w#�?u�P8����G�����K#�?�G�S�s{��3WX�	ՙ>M���U%lZ6
�Ou�8N#F����|����{52/�o���%�EB*D���_�G��e����>��6a�m�_�����I����#*x�������'�NL�,G?�HU:���=�{y"�(G�1T����3G�h�8��}�u7l(�6�h�e�7L����ڙ��ǮB����Z^q)��ۢ)�_ə�˫ccC�x5^�T=���O>~�>��Ei�+C��D��⧽�6��v��kXk7�C$��]�yX�*l$�8�s���̾�U��y�9o�"_�~_c#�de�=�q�v9!��8�nW���'���'/iCX�8X����ƅg���j�J��u�"�/�V��E�m��������X��]���h/�>l����_~N�?x���t�v�ή{���a��o&yR~\�ܹ� '�Shj�=�����ϰM�%���!x�\����|s<_�w���\���C�dQ�t��Ϭ�uu������Q|.���:�:b#�l+��8]����<u�Ơ�҇�ll���L�,��s������M��vX���p|m�a��}��Vf��ꈑ,�ei���;����]:$��s�ͅۥ"���6:��ār�
sq�^u��>����:Y�Ngl����S�C��	Ҵnq�ltn u)[��Y�3(�>7����[������:���8޳�m�����m����u:ߎJ*M)b72� ����UNl���2��Ŝoɱ��$��2�b(:��F�	�/]�!{<--�{��A�w ���qpp�p8C���j@���T���uy-�e*f�gY*�7:B�P�z�{x����SG����a����rܼ���=�^)F�e���,0���l�'�pP�r����Tݨ��U�et^*K��^$$A��8$D��LG$A'�yK䍀�LT�*B[Ӣ�BN/���
TQR����3�6TK��A�#E���!�Z��m�!j�J+�K'��	r#��2;��Q��?q@�W�ɒ�(s#
;a��mqU�:���{B_*(l��ڧ�P��:ӺkD�C�Z�G��9I�d|��|�Q=Y�� ��ܥ�(@�\���ßYj�i,�k����>�|���Ҟ��4購�Ը�o�&*�*��o�ۦ��wiy��x�\��Q���`7�R-m�I��!x�� �賞v�C/��	��<�Uh�뛇�A���U�ҕ�����d{�m�ո3���^�덊5��;H��W�k���6�G��}N@)eJ�u�g���)��� ~�K�´��5�U~r�7���|�A���ui�(�����K�������I[]�n߿z׾���������o�h��߷����������_�/�����_�����}��W�/~������~���������]���׾��ߵ������7_������:��đ8�dme�s,_K�1�{��PG���E�ꀷ�r���\:�X�� ����O�;K#��f�G%O*����*K|"�����S�����V�;��^1M�+�k� �J/��-�6xe�W�`d�=�=|�������  ���8a�n��j��+�|ptM�ׯ1�_��w���Ɩ+�6�����vx���
�Ǘ�o���υ9�K�4��m�Ơ���� T���p9qu �eh�Et�>K�S.����mT��1���s�]焣S\�ť�ӳOB7����Pނ����o��
?8|�/xQ>u���\y���7�w�Woll�����C����̹z��7�{��F{��EZ�j��-��)�B�x�˹r$�.y��W�_�/�������O/q���|9��d z�C`:M��o>U�AO)ϤTm	��gW�sD������SI/ 6�D�AUc@��eC�i*-S�~m��)=��y����K�maq�MLI7�x�2Rzѭ=�Bn�P.�,�� HD|[�*�>C��hٲ3�V;A^��v��mg�����Ņ΍�`ʮ:LK'6������!��;�ɉ˖��SéCIO�㳻c����WTT� �&4����%�������g���=>="'��}�2?#������J<�yh�� �����ÇqW�o�߯�ϵ{�}'�i�^��߾�����&�|�����xG�Kg���n�@x92�f�/�̆��Fo5k��*\�!�����G��7�͹�xX?G�i�H��r	��(c�ɒ���2&�}�r��޾���Ն#-� �x�P*�u�N��H5�G�VKU�*̥��FeEL=.Q*��V=���c��v�?�iG�8���7�\��������3~AX�v�H�<�ß:�4}�s��>*n.xȀ�btBU���
�*נ�Z�)(�Fz�� ���V��Dpi/�p�寜(�Te��O΄~Br�P��X�и�wJ�ri`Ce�f	U��|,�Q�r��_�o d\�W�Q�Щ�7NGO��'؛)��2:G$��MgL�̝��f��B���;k+�J�m`���K��;�;t�F�>�z�>�Au�� &��&�ly*E�qzCN��ӏ�G����b�N���8�6 �oe�2�i15"�HB�#!����T��8� P~L/�Y�OL��4�vu̇)OW�+�;y>^&P�r2O�|��ƵG��G�Y����y9�ų����2�iM� ��'Tu	���]Z��<KO�|=���n:GһB�a{h����+}̳ϧꞢt唗��N(W$j���7n������pت��H��ŅÞ�k{�	6`�R1f�Kt�t�t�j�+F��r}vn��E��>��� Ĩ~�G�e��_�������������ߴ?~�-�����n>���{�}@qn8#����t0
֛𸝄-Ŷ��6����54^�r�C*G�B�a��a�T=�e�G�qj+��������/�u����/��qmY+\�Ax0��Ňy����=D�������'�Q���h�ޛ^Z�u���^��ӧ��Q�Ѳ1�غ����a{�a�{�}��j�������N��v���S���c��bg]�݀l���)�8񬑜��6�a����A�Ҧ#l����QdyB�#�/JV!j���;����K��^��*T��1�.�E'���0�S�|����	�X��y����}�N�A�FXQno�+���w��3��0(G�8��՝0�j(.1�gfgg���۝;CZ�܏�o5O��AR,�`a��	�9{w{+N���z�����{׾ǡ�c�Ç5�ҡ��Oy���F- ���`��M�r�a������U�a��O'��U;%]��.���Ξ�����@C�4l����O輣�iꏮ������w�s2��[秗'ι׈��Ơ�q�I�Ot�mx��I���c�������v���3�u	\i���q6ۛ��mee�mn��ce����$e���s���+��!|���7�2j��P�����G8
avr|�V?l o�k_"����e;��Sp���"���	��N�\�^��4��O7���Z��e����w���>��{t&��=�62����[�e!�~�7GLػ��q"wkxl90���NW5�,t�ٖ��ٚi�%偅���U��u��B=�^\?���'m���ҙ�t�Gو�@������5\p�%���2:꼕�6;_���n��p�%:��R6[%�k$X��Ka"	Ma��+����~ O�>n�x�>p�Y>��� ��w���F[��4�
�㙧.D1@S����r#Z�i`�O�@R��9k�ݜ�C�i��;��\1f�G
�������=J�8��&�)�li�b%�0.���,�X�i�~_��U��pV���o�z�Q�hSً�s���)�
֜�	�.��OVĘ�t�>���D��"�t]Т�E�P,��/�T�)E"ê���,kװ��q�a�������tЙz��a)�B��O\�U�T�Ywأ�!�xO:rr��W�A�%m���n��⑎dd���v��<��nރ�3�i�X׸�G��d�A����8'g*HǴ[;�]T`�2!=���	�n���~!��t��Q��=8�W��U6�p�pXOJu��-��ӣ����)|Lb*�]��Iz��H7*���8|�+�^�i2!
e�B�0Q6!���{4:��i ]!��I���ԇ�"������Uߦ0�z/�x��B�6�(\�N6�X/i�^t�e��=m�$�[�u[�v��z�3���T
�1�I�r�+?�R�C5bT\�b}xok�۶�>FE�^NU7q��� �Ň2P�����Ƿ��_\'P�]+�.��~ŗ�g�>��W�g�1I��G��Pe���,��a62�ak���F�o�GG�0�6�(ăݽv�<�?ωo������01���=��R������a�4�����vA�����/��o�V�i�(�f�]Uu��Q���a�w�g��&U�©;|]Qn��OF�>��z�k�9��'��^\�����*.��Y�u��#F=JG	/+�Wn�1	���\$�a�z��+lz�#�zd���0i�ԯo��������~��mc(/q0Du�ћ.�9	����A�B�8sֻ䒍y6�ڠ�ӯ|2��U��rJ7�'���TT$�$�Jf��J�%^��s��qˊ4>�j��E��)�Y����sE?i�tMK
͉���Ū �6tMYl��Po�n�3��ߐcY�By��T�S�e����\����D:6j@:GN�^]�Z'��yԏ7��ki,�MC\��������LH/��7O�a94޽�v�i}�u����E.p0����x^�[���ġ�eu��	�Z�����,��c��(N��0r�tlD����aЉ�ђ�O��i�[��i��Ma3�iϟ}�~�$IC@�n�Ỵ����z��3x��F��!{����Η�tn�6��҆pȝv�Ę󠔏C8�C�@��Xm��/�㰾ko�}���)�Ii�j5��w�q���A����v���v�9�y�y��ZG���O������՗ߴ�������E�8x��(Xؠ�ba�4��id��]�ys:ͺ�Il��7�E/�i(3����pdtN1B��:/�9x�m�C�����OK����Y�0F��sf�5����<��4SqL>�+�7���Z�]�F7�bi�c�T���%�S/p���P�8����r�&Dp����<6��P��H�]Y��}W�\�GT��������/V7v�U�lz��f\���mm�:�W�:�!��c�����J�, B�n_����(]�a��g�~Ҟ?����ٕ��iƵ�a�}����w�7������X�EX���F�x5�Bj	j @�	�:'k{W'��`0��N��e$���M���)�܏��BdnS��@|��9Y�)��d9��=��!�`!' �"��e3A[HPq��d��L�/Չ��,X�Dr �.�"«�]���|^��iL'�4TD:;q�"0:�N�wN^��N�%.�	+-k���L*�	C�c>=(�1�[���V9����W��-��5�k"�+a�)Hlvj��)`ht���V pٕ�ɶ.R1�3� ��F�P��8��:�6v�1�-9DA'K��w�,�F�-m[�2'k"Ck4�zC7 ��]����}��DX���¹�j���Bg:Y8^*nC$>���)�p|b�DX$��\�W�Bu�bY^P�γ�z����|3���˺�ꉤ=p��ڢw!�v��n$e����CDˮ|qN]�����8���S�9��k�u-� �����\��`)�T������5�䇲W��`/Y�У~s�yh)=�qЊ�im��I�'���F�L��E��C��A$�J��O��0G�+|��/w����1�#M�8�����9�4�j��J�4r xa��xMa��ė]��2�5�:���t%��={�p�ڡ�F�����\	�cx�)S��K�ko�έe��P�I��rd�5�\�R��s�UvA
�D�P:?��̜���t��ߣk�1�e'!�:����#|XG@�H��'c���J�}���cI���]�Ϭ��#�ܿ����w�Mx����(�!*��4�=��u�.��P${O��Gqr��� 	q���8k�d8o{�mlb �k��su�=��.���c��=��v߱~T�F�K(\z��'e�Q�N��A�-�F��`F<���])1x�h-�y�����Ёu�i����rP�Lx�)�h?
+�D嶺�{�t2WG4AkɷGd�B&���P���O�B~�4C���*��<�;n�#,.�E�(�l,:8��
]�&qġ��[饝��*Ŵ=|^�\|~�gUV��ſ[��t���1/{	6���p�]I��H�B�\�p"K���W�V7LL���r�W�������0�u��*����#]��{��Ֆ������:�BJ��)�����Q����"���p*>=9��8�>��Q{����
�����U[��o߽^i�� �������ꢼ$i �0��SæmT���8/�wʬ=�z�s����^� }�����ߵ/�z���W���3��X;��؋�Șml�u�y�n��|�Ҿ��U����S�7�,y���;�ǽwp�����6���M��߿�aڿ��{��$MV����R�֨$w"]�	NV�0��C�	��~Bg����ʂr_D)IcRS霒[އ��Ǐ�P\�H0~���)���?�4n(�A1��yR�L<L+m�1F�8�N�Ձ��~���e�����1(R�d����)U�f��[~y��aO��4������5��8S���qv!��+l|Wp�W�����i[;N.+"�_����ZVvyk�QӴ:��h���_ �Uܥ�I�I�*�)X��D8�9a�铏��~�y{����hG}rv��	������K���_�x��o-�Nː�R�h�@�H$?e��O��>̱cOV��Ӷ�Ԏ$i���CF��^{V�fX�)Z/�D����B$ԅAb�څ��'KcP�.�2�R'F3�C�w
���U0ֲΘ�8C%���pC`{��@�k���1��. з��Äd�2��L@q���:��$.�.
�2(@���Tx+�u�B��AZ�-����:� X%!!��(A�����c'���A���"���`�2O{�g�"���;TС�1&�S���0�8Y#(y�f�<����@�ͭc���C�Ƕ"iD�x؊f���dzN��(��_PH��N�%B<C��d���i�7�GИ�1p6���p�g�?N��d�Åf�4BL��x�{�$�`it$�Ƙ�N'��:"���PH��u�~��:Xn 8�L�6��v�LyC�)n8�P��
%�X����jy����)s�Ҙq�1�eC���Ө�Y�{�PWJ�:Y���3��d��+眤~�iy���Ic��r)���*��<]�VZ��"pL�]���w���J���J�>�5���H�O؈*߉�ß��.��t���U�����`��5���AZ�1���,��9�fE}��VpP�2y�B�rx�6iȗ�]���l�1�N0F�+�$r]�RW�م8���r5pʒ�aM�g���`��	�4��am�~_�SjșC�g�D���6�򋓕�����x^�Mi�kj������G������wU�Ks,�(�RSǟ�0�ٳO֦����@s8YнE!2��C�^"[��8��j(:|� �Yl��s�0,d�pS7���6&.;wpԶ5���3�cӍ�wt����}�����3�
{���A]��+�rYtq���Q�����ټ+���1r��cѪ�)�w�9���芒EE��eg��+p��#�}��rf�+�����D����;�y˹J�)��c�S��r9���_�5(E�� �rߎ44��q��@��KP���p��t�4B��<��R�jE���W�u�~U��9:�Vu�G7���:X��vHֶ��8H�\ҹ���v�??��݀��)q��q7`��ψ��əȅ�=�t�LBY<���k�QV9-ꑠD�4~����2��������{��9K5r��3���]�<Nt��h��meu�}�ݛ��oۛ��`�2E,�h��AK�@˱a	%�K�A�5l������u���n����ͷ����o�ە�mum=��8\�q���՛���˷���^����)��e�����ն��a�� Y��먽��޾}߾���o�_���~����ng'岧J����Βy!2���;�\]�Dm��j �է�ՋEd�ڠm�;�׃�8�ޤË�E\�������VB��N��K���>�A5�9'W�@ʭ~o� �4������p[;L�]�6�y���]�ިBֻ����Hʅب�ԉj�y5�d9�T�h���K�|nח�]��J�#����R�A�6�1����8Y�BƝ�5,�b�aK�v�ݫNHe��'��Z����+ �`+�I���� ���$
 �����M{��k���o_��w�ݛ��f�Dh߿��w`�I��6�ҝ��A2�&���!�b{�mn��D�LP"�0��V���$�p�L;�z����3)�h��+��!B�õ�\*�;�8\O`g�.��#dw�Q��#�$�_Th����(T�(N��\- �14����Sq���Jx�J>j(��U���U2���d��"�vfI�KTRj�bA��(�c��G~�P�'��!&�w���ft��i���q)b0�ÏNtz�"���.�F���;F�jy~���"[��,�8���U�2���:��/�v������˶�u��6Q>nR}�n�;�mo'J�Z�Jg�S�E�\�Ѣ.�Ӥ=��KϨ4gv	�FqX�p* ��P׋�穑u�4����^8GI^Q��g{�3Q<�r�%�!��Y��Z!Mj�A�C�!�EtN��8e!�es�F�F:�b�^N^^��[l�s�
aC1�@<���G�\g��zC�B=7��}�B���f�_�Gu���Eq��h��2nP�儭�e��^�M]�QMz&�{�S��R�@J��C�UD~/t�d��5�!���������
q�*�e<L��%`�:���J(Z�˽�=�M}�x�CU�$��PT�G�䛢��%N��$u����,��gWL��1����L��������&�9��#��y7���_�u�a�Q��p�
��r��,i�ߍ����4u4-L$3�u9#�k�SW,Sz����U��p����a��|i���~�ga㊽�6h�i���Gg�B2UW�7��4��"y��-��"��%xm�����(�ټ�}�����X�8_�w5�h+h&m{��oW0�^#w��*�N!:���?�;W���vN@�N��C��돡,L�un�n��x8�j��`\o���a���y[]?���[8X�m�x��M8�d�=6l;J��C<��3>2�̀w�4��nv��I�&22�ڢ}a/�88���������F��2�κF1ur�`�����!�c����%:@���MΎб!�4��p\y-+2�>)�5x�\\g���1��,ϥ#�����S=�}�㪤o���k�W�8+�x:�C�7���:F�F�������N�8b.g�MpN�[���\ϳ�zg{��&���ǚ���^���A���Cw����ct���H;BqA�ĉ6<}��_���u5�NN�z�U\����=%5|��y�U|���#�����6��w����A{�c<��C�0p��:�����)�A �&{�u����:J��S�mjf�4\�e��_�i_�kDx��=v�a��[�H��.��E�3mxP>X�����ܧ����n5N���Ǫ���o��������ŃN�׺y��՛�[!����W+|�}��N�����\m�`����������M9X�
�N���xՑU���@9��\�gn%���Q9�\��ϱ���ay��0I�G��H��wل�N��-=�a��$}�'�6З���9����ӛ���JOWæ��ӤSU��6�6SBl���VG�;m��{��> �ٔXz?�6�;�J�)�T��|/���+g�W=G�D`k�u�O�GF,9��>q��+8N�-g	���4l�s�G�����vqz B��'�?�m!}g��J+���m��d*�J7� �KZ�� �t�^
�E��]eBĵX��0��>��Q{��>2���x��~����ΫW߷��u �\�{ia�=�������L�ތ� p��4g낍L�k>�C�\��@'��@w�'W(���!�����z��PPtX�	����-"Z�X��=00d��E�Wc(�j>���ڴU4A8��=B(���ٚ�r���9�uxL�O����N�ecP�_�+ϬBw�	,s�b� ��x��i!#��9����x/cس�5��Ғ8�t��	m��YL��R���P��B�V<�5��A{�\ahan1CG�O+eg\U����Τl=xG�$xw��E6��>�6 vx�ʺZ�N�[�u*Ӻ#Qt�̈́C�0\b����J��=P���U��x )x>:|;FZ�+$�S��a�'�A�Xv�~8J/H�Q�&
�>N�|���P�8��^����U�p|gg�0�M�KpO"2h)i�gjn�,O�f��6B�|V!-H���8C8�6d^�JX���U�g�
=r�Ғ7"\6`�Р�e`8/��ҁt����|ÿ*���*Y���T����9�N��(r�z9Y]!�_���Ǧ]�o+w���p�{x�yҴ�>螥l����45
m��� r�+h�,�^u/�0�.'����@����DP�r�tRJ�_�� ��`���[�M��q��N���U�����*&�&��#�K�(#,3�HM��%�#�\@AE�(Gp�'��id�v�����ٕ��)��6��\����H �<��B����?�Ịoj�^�H�7�\T�j��¸�C Ma�ool���o0�>@37� g�����B����Tl�w�����a�������b�cw���G�mxܵ��ph����~��`c|^ \G�)������ƫ��@B�&�^|&�h��PT˭!WF����h��v
f%S�<�Ƀ�s:X�c�u��<Ce�o���ҝrм�9�u���fķ�d���~���r�6�1hp�'#�A�q����3�A��u췯���;p�*kkY��=�ֺ� \�}�mm�*��Ȝ5d��z�Yښ����kH��\�<�t��l���ԧq*����L��z�yX>O���8=Y���.���K8;�_����G�~��-�q�&�'��W]!�9�h�_���";|T��[������A� G�,�N��n�4��vEM��lpX���U{��^,�o?��wޓ����j	 ��Ϥ/K:�Fҫ���<��_��78H>��#�Y�e���ݥ�]�Q<8�m\8o�^?�C�b#��(�4��[c� =U[�-xoO���BK~�N9Yf��8�\��Ϣר���	m(�ɲ7+K�=7���9굸�ׁa������sūp�>�
�c˨�ã�,�S�2{a�ٳ�Η>�x�{K�؆�ӯP�V]���@]�=nT�+7%�h͐�S�~�H��g�u�v��f]��v��4���"~̃�&�{�]f띋6��7��o߬��x�{��Do��w��nq=�X`$�~�n�ѡ�:Yz�U1��X�,A���io��
>p���ۙ0fK�im�����^� ߴ������}"dt�ݺu�=|�s��F�tz���Eb��c������d���*�2A��d1D�Z�P����!Ir������?��1@Zk�Wy�$}!��,Av�-�qԼ����?�둟�� v���"���1�d9,!K��L�0J�a���1xiT+S�Ͽ�>/��3��r�nr�@i�R`C�2��V�?�:8�A����4�%��y*e`�`U��=~zz��C���lnKy�ޡ(���*KK8YWY�U�G�e('��ɢlap[�x��\[�����p��v\�R�g++���v\�!�'�u�Xؤ'$�PRW1
7[��x �`��h�P�/=tN�����?�PZ���Z����Ca˝B��.��yΐiq�J��)pKY�sqB l��� �WO����k'k��M�g�"� �8Y]H�4��q^�,���<]��I�y&p��T�oN�C=�R����� p��>�4�H;�M��ټ9�0�5y$���b��ܫ�t>�1��r��@�v����і�R�.��˧I�Ô*���ԛ��{�"0'�>x��{�|0�?���h���iFv�`�W��0V����Y��~p���&�I?T�#n�(�KWɫ:t�,ύM�M?��aސ(��3�U����Qɻ��MH	^
ݒG���!S�C�"����	�cLZ�d�/�����O�-!�=�H�}d��:��7� 
�}�|T�wy҅�����Ht���C^�8��< ��M\iN����O������rm���(P�9��=��^�"e�&lpsI���0zܠc�
����I>N��N���E��}f���kh੭��#��v����Trs�U_O񑡢�s�"1Ղ-̕�|�Jڰ��$u���ENT�G����"y�N��'A4C�����P�ǜ��0�1��N\�0@�7] �����Bk�XU(��a6wg�W���d��:ћi�fp����|΍͵�T�#��e��0e��:v��)�NM�?,#{��F��H?F���j�n���S��1
��f�3���CM1�A���(_R'�"����.NU���=��"���<�u�z����o�ᗆ�J���	-��Gm��!pw���3������ɳ{�����L��mG���7m�v�K����vM��|�2�+�l��@+6�;j��M�U\��%�4�Fq/mJ�?\��߈����`:W�N�F��o�����C.h�^G��i/[>u��ߖ�;UV�����\=4��Z�Qk��*L�(@	od5���3�'/�A��i�vw.~����\�I�>���HA���y���MR[/�a��4���C\mԗV��^Y���C��dy�\��y-��>��)��w���q�^3:YKw��$��f�w�9����.^y �z��D\�[H�����,�`_�����z^��x�xV��V��M��~H�S.��ot����Z��K�λw+mmu= Q�05Ysnz���� ��y�7���E��<3����Gwm<#u�<���s[Ő�}<�����d�>{%܄]���x~��KW�V)���7B�3��D��Qa�/� �
d���)&L5����rw8ˆ��
��u]���Pc��	rr�Al����
�|�5}!�M4o[�Lە#T]�[�Tl�ȷ�S��ʒ�����P�Y-2��A�)T��LE98&\�������\'�Q��|���_KP��:���2�
����L�Y��?"���_��Bz&bh:�9_S	�^8䜨L�E�åT�W?�-�ܼ)hH~�_��u�^7�t#�iҞm��s(^�4��Yߠ�Ҭu�v]����:NSpไ������2��:�����]p���u|�B�<?��_^�7����tp����3�{9��c��q��W�-����߽s�p����g�^�y�=��.�ů������K���yZ�4������K�T	���#�����,RB<���6�����sR�jF��	����ûp�Μ�a�����hw�CV&x6c��mힶ����N{�f��z��ެl������yԶ����1Ɯ��t�g�k�x>��l���G{NZ;�a�:�Qj��A�ʷ�1� O������	v�I�hZO����
#u��Ѳ�*�{~yT(�<��G����_�	U�F�/E��0^W��ߧ�{���K���iϻ�Vz	��Y�<�`w�L���fH�Mf��t;���NG���E�±Z�>l���+nn9W�
'�!���j���'����Z�q���KGF��1�l,C��s����Y����#�רM�uB�bx8��L)�4r�����/� M
�r����^\���u��85]�N3�]�5���e|��"���ʍ�1f��C�5����{���)u�1A���#=MЩKU����q�C���а�q��j�v�H��52��b/�7��ҷUOc�bȚN����`��n ��sY �!1��a~FK�Ҩ4 �*^f���U���klq���§�	g�'��~%�a��G����#�v�2�jo���min��Z�isScmrt�9:�����Gq�ƈ3�&��(t�t/�)��⊨��x�tR�K�mDun��d���/=܈�9��
˽�-�euX�aP����|��W�{wx�<��K��:��:�!t!=F���lx�FH��E��[	=ژ\�Z�K�=��R)k�A,���<��Wֹ�!tgi�B�����t��M3?	_w�4���N{��ɟ8qzS��ڑ�)��LOg[4�kѹ|Y���U�\���ewT�s���{�����u�����A�9h�K�&F��W|�#�9���[F����5a3�}B73�\�ɵQ!�K
`�E^\Zn�o���������,I�41�Zk:2"Rg���A,��3�]`93;�;�}�z���U�]�]"Edhu�������7kz�{y���9Ǐss3s3���R��L�ίW��"(H�
�r4�4$R�ɯ����_��8`�������W�O���Ǘ�����'��U�����%�g\Ю�6��������U�dj]=+��\?���˞`{]� W�c�H4.��Iߜz7�����5zr"��'o;mtA�!�v��̧��{�JOqm04�lL<�>=��,V+�d�#�c\�H3���d��P��r��S��<� �N�9O��v\�1�u&C5}�A����(�Dfd\��_ʷ�k��x�w��T�k�w�I�Tm��5Q��g��4�=�(�*Nn���~��/J�T���GΪ�Z낺E��,�9bL�x}�Å8�h�d�e��0��1�����R�
�bh��+��B�x��z��r���%g���tR���6Q�(�0b�K�o�|F;w]�6�n��,�V���S�vVL��pW1�hQ�ʔ �]�� ��iee������F�^�Ay:xKt��z|\7q����{��^�y����4(-q`�g$��uX*�5U9�W�0�"���g������<N����b7���[cGyco*��V�Cn>m��~����=-��篷�ӗ������������n�m`,�aDa�s}�����c�:�8=�s�4���������ȆCY��8gg��Y9F�d�\�>ęm���G�����W��TVa�z���w^�+���>x'ms���ѥ����7��L���F޹�j�4 �1�C�!;�w��ݭtY����5�����q��1�c��a�b`�gS�-���9Ɩ�m�\���>�����q1�H��4�5��R/��t#��u�j8ݳߞ=�Rg��с���IY'YBO����|�r�و�ߥoT/��9G:�y=�g0i���J��7Q0���~�����H�5�*Hɇ�����w^���{�����%�K޲U�8�y�o�Yk[������o�&��Z�23]���Q����S�mEG�+�t���=9'rf6Jl�}�"_�c8��|K�9c{%p[)镧́.O�\����O�4i$��WI6l�:��@u�x�rX/�<e}��#��뮹kd���4�[C֛zy�S�K�N\m�"�1��e�ҍ�331�f��,x1�4}�@6��)�����6
@.(����!]U��;�D���]�U	��(#�|���Fm�pҚ�î��1:���鵎�h�D3}i��H�pq�����N��Q��1;л��m���p�*����Mu�W�u�V)��M��P>�z�:o�4[<Y���q;�V�ϧo����j5�]�1�����H3��O���/6y%�>��_����r]�6��.�[�]�����'�L�)�r�x�o��R�<�2�l��U�qg���p!�HR	0�(���3�R��;��6?����n�;������Z�n�e�:J̃q�|;��DA��2�^X�)K!H�sP���v�w�(�Kxdh����+��K.�s�h�'�X�u+D�f:K�o8 $\�U�ma�@)��]�����r�N��/�3 +e��eo�F9�Q���i�h��N���n[ۛ���*u��5�R��g�^��r���l�ah۩uМ�D)��<��[z*���?���(�=y*I�H�MZ�VeP�Upn<"k"tćF��ZM�#�q�.(��H�Ο�^��_�T�1�G�W��.#�(��bQ�������wD!��p�\��?�Ϻ�uD�:ze��
�=�Cc�2MS�c1�.�#���UJu�Y㽦���Ak7��I��40�..1�4�F4���F��J�\�]�Fe0m��_Rpp���Hw7����%,�ϑ�׏
�^x��S��#U�*���j�֞@q�P�)�#�q�a�@V���]�o���2�r�89re>��4~�5�M���z֕��sd�r������W�%��E�i(��4�'�����|M]ؔC���K[�i���jl��!�UX���|LKG����7C0b#�P�I��dX!�]z#^�I���N��0r��=�_��������a{�n�={�۞��k/���w���NƠ��v9<Ӯ��17��௎Gi4�4����0x��>�3�E�Ș�r�����F��thk�:R�����Ҡu<Z��{�������Jeq����? �5�*4=`{w�����]%�	mS֍2ɩ��#F�$������Lf��!8�?��U�Qg���I{������o����C��Ѷ�7�vv����q�&8�Q��R�k�q7iڈ	��L	�E�f@��)��1N��
�V��5{�k�[�
�<��n��]T/N�w�G�;�bt���;i5�
���O�<n�t32�b������bG�}�>�&�<�͜�%R�(E)���SֲM��a]�~͜2ǚ�^�-�9=�0���wy;�:��5uk�p�/�ݺ��ܹ�hg��&xw��s�د��C��.���?Κ�[������=�"�I��l����u�A����S�ڹY���?�M��k�q�|SF�r���?��%|01i�k�3�Y9�kB��4��c�q�S�e��#�i�L�/��~�G�&_�735��V��Mr�Ҙ�4q��҃;szΜ�t����#F�5���	�8�e9I/�!vg;�N:Vu]�z�{H�Ԗ:�ʷ�|%�2���ӓ�a����YG��;�B��60k���/|�Ͱ��G�s@�V��z��g>��dCش���0ҏy�Jdz/�{��jC-G�	�^��ԻΟ�q���m�y�˥_�{b$�\�RI�{-G���o>򗎇�շ�����q�s^I��������	���g��Fǈ�~h��3�u�I��(l� ���nu��=�%�dPJ2A.H%a��D�V�'�MaP��|j�ޖ��*������۷ncd=��p��D��̆	R�\��~��nfOy;x��\�`|�F!�2�?���]��9��*��ӪP�j
�~�>SBR�)�d`Un��l���KE#p2�/�NX�2��bn�B�8��$#sen6�g�%9u�~���-�u�ٚ�P��F����?���.�a�2i�2\Mՠҹ�&i�9����������a�*Gnn�+�C��BB�7a�^~ݢŞA�h�Z�]#m���`�H/*����:]��c���M;�n���8/�a�/t�q�i+*}8RvsC�E���!� ,SZ�4�0`��_k��1��Ѭ�hB7���9�"��3:Q����2���U�,^�ޫ��2J�)��v
�i�9k(ܙͩZs0�Bw�ĥ6��5���Cc|��p�۳N��߸$帮n�_�&�D���m�4R��]+)櫟<b'OF�=�-FV���o=�@e��ef��	��j�٩L#=�2���!󈈥�Z�'.B�����ާ�A���#��)~��:j�w?�#��
�'4���:|��1�J%�6�;�{]��3{Gf4Q::7<�nu*!���6Y��0��4��%d�ʙ�Z ������mcA9\Oa�nO}vfSI&�9�_�k�΀�|h��\����ݣ˶�{�)���ap�9l�_�����h�#w�t-��!*n�;G]kt��n6���9Sd�q�rí�=(z{{%�8�v\�*P��.M�q"jo��KCw����o	�K����+/�qE���.UFwv=���o<_�Σ��lg����K'�퐇a� ���Ĉ�T;gm�C�1������Wm�j�p��cmck��F\�w���xPBҾ�}�|m�3=p�;(�|���Ƴ�-=�x�0G�(+M�W4ûГW)�(����(e� *#	�#�w��:s�4��$�nԁ0��%Zfc�I$ySE�F�����NA���|N=-��s�K���+�	q+�u���`�q��Ó�*�I������_�/p��n��Zi�Km^�C�Q-ː�w�i
��)t���=nO�<n�k�ѯz��vS�� �(\�5�e	gu�!����sSH��$��(��U#>�G4����g��ADd	,��i�I���w��mc}�{�<�g}ZG�QR�{�x��f��	��^L�J�=](��'���2An�4���12�AP�$/�GxqqE-��+�8(�>kgCNe`���T�m��uX�F։���XxF���O���'� {�
爻h���ۧ,�p��j��t���e8V9���<3�|�A�c�;��Ug2�q���;�_����~d q��I�z=���HZ]��G?r(u��=�2�OKZ��׍��[�g=��|�g�>����(.�f Ǎ2��6����X�%���ioɫD��:�!�y�;db2g��F���1���{�Y		Q�_@dj�h���-WEIL��KZw0��{wﵕ��2[� ��tU���^^�`�z�y���^W޿��T��{������<���i7J6�>�/�*ܸ�M)QVJ�d��)d�����b|�'sW3�Ϟ�s��"@�ӯ��4j0�~1�!��jh:1�bh����Bi�q��d_��ʖ�(��+���@�IGy����� ���S#U��it��*�<:+;���s�a�sW�>�T�Skʖ�����2�4Ԝ�`�T�C����� �cF7�Ш6{%=q�#xŸS!�� <�#�fjU-+{�('��F��o B��+ ��Ј�C����B�)YZ(S�Z*�*�c��̓�=�kH7B8�#����G95���hS�u���/ݒ{�m��q)�VS8��Z�T�aGh�/��4{��ޥ���t��Ы�W�>��tB�8Ӎ��[����)��S=����(kF��|�IR�i3"|Se5��tzW"�]�T�Rg���������������G�򸾀8��z��Rr���}X��9
^�Bgh��)U��Q+RY#�n�{^��t4��P�O��,���X�B+
𘍽��?�*�4���]p�B��p	o��
����8G�+�(G@s�I��]8��e�����՛����A{�|�={��^��k�>��nB�a�*�[�1��uZ�K(��Ցq9�H�[��o���:;�������/�������o�ˀV�.�<���^}<����q%)U���hϿ��"�\��"��A3!�w�.��)�����������=w��w�ĝu�/1��xnm�`�jez������+;d<3ҴA�áUtW:Ĺ�|7<�걗���:�4�t�ۮn,��s�=/� �J�Cv �4�&4����]d�M�#�� V{iz=l��V�Oc/���P��V^
��,]�ha�ؿ�:e=G�2.z�2>r��Ƴz�_��!��U�(>�g��n/�4i��A�nꥡ��矷���:w�������4�ez�<K��c��#`���K�2�2����/`�p�l���\v�����g�t
?��¥l�K��)�	!3T('0��pC�q<�1��ք]��7�6�)�M�U�%�l��|������L�5ʷ:+�^����-��N:C
#L�n��H#r ��I#f|�t�G�D����U9�K���7�݉�n�_�ӊ&y�Nm/�+��J��޺N�th�h�CV��T��$ԅ��)��dA�l���p$q�����f��v�S��X����d�p�{"F�q	W�8|�K��;�W��3��6˫��hQ*��tq�w�U�}�_ҁ^��V'Ewy�����u��o��yx/��_�n�_p�������U$*T#&0�V)���h�6�p�L
�2��.7@��S��T�B���p�7Gp�©k�4u
����v���ދ�c�u��i4�f�$
�?\���]g���J�q������/�=�{<�w�z^~�"={rh���S�*�D���^R ��.��U�ͱ�*�:�;�FLod9B�P%Z�g��4��`Ùj�R��d�x���[����{�Y��j�~��J��y��ng?|�N2+EN��F�zW�ghLAk>ǰ�����_�4&�z�� LU����\d��Y�!��w|	={��1F��=#FW>H�m��l#�5P��9*h]�W��)i�ǆ�q����L��5_��� �C��rT˵:�Q�6�n�;9=�Q�;*�9�����j$�[-��`�*�3�"G��<_#�c�1��&IK�@z�4js�7K2S88�\`��@C����!Y/�߸����M�r'���ۥ{3|�Y�����M�c�u���/�z0����1b�O8${��9�����i�n߾��!����z4ȯ�w �%m0����/��g�����k�ySq�[�
�=��4��ؘ�H��@=6�6֝��_��G�T�ª��a,id���m�UJ�.�4[�9
u���4����.�(3R�8��ʡȟ���_������Y/7������m�Vܛw�z�iP8jU�{?mM�Y��I{�/R/�޽mo޼��޷����9{0v�%櫊J�����_�߿�U1���2�vv�;�i��B��E��^qd��~�#�<4xck�}�؆��N���%��>��K�����6wlYwup\k�N1��2��:/��$�����i�Ϻ!�r���	�9�4���#RbŉMiO:&Y�����s����r^�[:��@~�ؒh�H�z�>�a���TF�iP���������I/�G���@��D�laK�)ډ�_7�i[����W�-���������Y�����$J�� @�jl}�����駟�'�����+���K�����yaa��ah�A�ky�7������",~i�-?.S�O���Ň2�ܴ�z�X]�N������w&�4�ͨ����X*�),H�1Mޝv9F�1r��1q4�z#GCK�j�|2 �ȓF�4M~I��M�6qL��4:�#h�_i�&�_��l�ҏ4��%���~��5K?��w����@hd�87Lt1t�,��-t���s�a�ߔ߸QGt'141}��/��;��O����ͮ~*m��X����{I�)K�2w��H��L(�yp�x�Ѵ��;�u�U<`}��F�.:RGW7R˯��4�өo����<�O�4��\	�=��u�ݏw�*g���I���&iE�s�i��Nx��o���^���HR������2^1d/X��B�P�Z��� ���L/�^�,w�S))¥�n �����1��`ؙTanYz�eˌ*��z�*d �k�Z���?���t	xųB���A0����c���ҩ?X#��-�ROm�Y=��T����S0�� ��{� <�@��������Qr����cۓ����{2�z��1���|T�;��S�GpRO�����!��C�� �O<Yy��lL�[8�P�a���,�
�Ð(e� �#�7a֧Ǒ��L�;-1#o�����M<4�=���c,�-�M�T�3�D�Ѡ�
CO��]�����\Ik�M꧃'�j��0�9��Y��&��e䥑�"[��`hML�bh�h<\�1�!����܈��D0�NC�*��E������1�aM�P{w���s�\���k��aI����_���f����S4��{� ��?��2 F����9&�<�k�W^�?�~��;8��j)�U|�l�~�����N��@��ƽ�-GH� y �����=��(�^�CE܄�]��e7���{5��|���Cg(�Q&m���'#c�o�GI��u�i��K���zeKJ/6J������g5`���W����5����uλ]t�ȼ�d}��0���N1�0p{]��-�����՛���m�`�W�3r�H5�l�,}P��!��4S;�������-�4gw�͈4��C\[v�.��q2 �?�*��~�o��է[�?J0��R���yG¹�_�Iq{dV��z?����?�������`��+�s�~c�������]dx�;D�����r�i�n�c�L�A�����L����lGT���EYlsP���:������|\ѓ~N2�R؋�2R�������2�aL��txu�1�-��X��'��w.J��dy (۝ ?���z�T�K�7��G��_S*��#�]w�l=/����a�'���/�ӧO�˗/1�w����r{�4�/�l�՟�i�����?��?m_~�U{��af���Tyw�SR��q4�����ق��q�����WX/�@�"�U|�q%mtm�#N1�iNk�aQH8R�;d�%�;>�*}��ް��9�˚1�V'<N���R�-}�0B�̩H��N��NGY�2�Ǹ�0�1�9{���>/��}�z��k�/��K\�{����!�|�V����'���*W���0�i�� �\	�Q��!wu��K�&�Hô��_�e��*Ak�n��墬iq7�տz���4�*�*a{��UZ^��^g�/����v�8�#�'�%-���^��]^/��ڙW�����T�t�s��l|3�^��]:Q6:z�.u��җ�����W�x��>�̨�1��0��iz��]I��K��	���dT���O��dEz �0# 0cw��%����+GB�%!{S%�^߿�n�~x��dyy�ݽw�ݻ���g��&S�g��r�s:�F��hE���`�`�m�h�m��=�@Z����)����s����5)QdI�������6a{�Bp%�@��%��O12r�	yd���z� �NiR���Lg9�;�Ni/����A'����L�)����	�0d���S��M��Yp�Ҏ�>5Ax��]���a֍FM���]Q�4��B|�]A� �(�	�[0gKq��)��M٭Ņut,
s���
L'�u�/���<�a�"x���`P̣/@33��nʞ��������/~hoi����]m���!4�l������^�iv.2������v
����w;`|�t\�葸j���
���<��Z���X���T2D�L���uw��:R����43u�2{>���
a�C�]s���l���ws�Y���6?�����$�M��,i��W#ViN���ӆ&�Z����|���f�Y�(�g،^bĹ�\gd��:k6ue�u.ui�.P�U�M���PƤ��̈�1�E�4�6:.)>����H�����ˈ��C�]����<�O�SV}��:\�j�B�6~ ��4�
��yw��n��k�(/%�e� ����v��ٱ�z���|�hJ:8�+;8�"'M�����J�rS�7l�ROOɃ����=2���R2�κùFF�3^��l5O�)�#;HK0d�K�ew#3�l~1�*�1�Q�nm8߽�����8-<A}({OΝK=��`x����=Y��"[��!�����}cAeʵ[��;�w�'z��9�sw�P7��1��;��y(tBD{�����8�<�:O�)����>y#�8q��J:G���w�w�C��_���'��ͫ���w�a\��ܧ�1MNbp��m�������6.i���aC���w��;��n�q(����ap���vL�O��`��'�R,��v6�h�(ߑ��A�׶���*�Y]�L��i�z9M:�hS����V�HdxJ:*�҃�M�<���&���?i֩��ȳ��5����N/<�A#٨T�M��;49�{n��<� ʂQ���,GX=�^]\X^���a�=�	��u�e�s:o��t P^g @Q�re8�b|��K���v���l�@���kۇ�����j�cD�o��ѱ�d�6ک�K9 })k��f�1b�i��i��;w��[�i��$y��E{��Uv�"�\�I޶����9����۹������\�h��8����"��z[\Z	^�j�a5��y����qm?�;�F�t������NGt�k@!b)�+y��g[;��tͱ��v��	�@[3�併���G�ɣ[�ed��H��p6y���C��<l������:��@f�)�9@��6��܌#�KK0H�$T��揍O�C� }����87O��l�Aۜ��9�27R�<����83���6>B�D�k�V}٩����x��&�k�(iY�*�mw��D?��m'�k��{�w�92�$�C�{`$7�i+�Ľ��lR�c䨿�vY��:M��\kӉ$3�x�]�u^�Z�߻ᕧҺ��ʬ"pmW̸�Q���A\˻9V:$�r�v�;�2�6�KU���J&x��_���<�=�e�oD��P���lC�9tZ�PF��Ó�] t�v�MtfѻV�,�0J99��?��_��؎�a��& ���1�2�-' �=.��P8�1�ɀ)��"_(��u�Q�U%]��ȅq�k���$����i�T$�7o޵�/^f]��^KK���[���b�AP�K�f#Y9��We9�ă�߿�4�����}��t�T勨�e�@W5�%4���g	��]��%s�^UY�<��,T����yp3��L���l�] �&�d��WcV�ĕ�$L	��s�Z&y�SI� 8|�h�1퍝��S�mCLa�h���\���4ŷ��P��s+��VY�T�֡�8Re�K�Qa���khē�b�ʕ��
� �|΃7Nm�壄|��1��Ν�U�:0a��ei��ۻ�iX�>{��3�y�2 �R��4bG(ȇmc�(kvQ`1��ZZ?#������6�pm�K��gmM��b�+��T���M�R+i�B�:�ӛ�덬��#D��Vi!M%	�+��a�h<�`H��3�cc�ԇ� g���n�M����GF栅9�7��e]��S�%m��dL�� O�X��\޻+��W�k�
���KX^�/ك[��^!�.�o�uS#�N'�n2��H�u��\����S�4��|F���o��g��`?
�|�7��������4Z�e��S�����E��0J���,��F��C��p���'�^6�p³��E����t�<䒼������Hr�f�%��y��?A�]<�I�q��T�|��em�k��O/��^(��F��]���G|��׵YB)�Q*�K7���Sa��a|y/��uMnؠq��$"+�Ѯ��RI�����JL�  �A�>J� 
4��p��8�R�
���%�.R�]�ԓ�1��s��V{��u{����������2��P�/ol�ͭ}��a�S�l���g��Ä�
x|���8
�R����4_`��S��#�U*[�@��
d�l��1q�3�����t:�:*9�<���{�2[R�o^�i넧�~x��2BT\�"����:�?�r�� �ЦD��{�W`�EF����$��7C�I��N�(#�ju����$S�U�mG��VM���7�w�,5ãx�.�s���l��j���L#K�N���I3�@�/r�mw2�����Y�|����� g������b�aݹs�}��'�.��;�������^�z�4,�#9d<�ybjz����
~"_g} �r���OCö�Y����K��s7�2�Oq;!�y�
u�7CA!�4d��ęvFR��{O'�i�(���y4���%��jN[[�o?���k�(a�up��?<{՞?{�i�v�؉���1�a�����C�ſ3jRǕdh��QK�I:�^�e-i(�K�BX��#׫�1-/8��YG��}��x���U�+�l�<�փ��c2��Ϻ�{��|xVގ0���KKnp��)��O|_ʤ��<'+�
�i7)Gd��#YYo��旎G���\S*mc��^��脝�6Ô�� ��Q_3G�H|���e�?�^mM���>�*��T�}���^�)O���f�S��]W:j�F�o3��Ҳǹ,wz2�g�z���c^�O����Ň��4Xx�����(�)�h6sq
�Ea�8�2�,b�*~)�*T��
�bX�`r.�=5�kh����;�,Bl�j���mks+��dw۹s�v[��ܶSH"!eҗ1����ɩ�-Wi�bd햑���p�I����<�J���1���.�h��.�{z7��xC��'�FU*���S3��p�a"��%QK�c���H�MϠ�%��y��ZX�]��3�D�d��"���l�������֯DRF�,��g�e�����͎�`d�.&P�J�9�J%�j�+_1��8nCg\�lX�M�S�#�e�(����I]ڰYƚ��x����w޷��@qy�i5v\^�A�m{���?-ee?8-��.�����H�G�i�nza�*�
/F�Ʀ�0��gV!;�Vsj6|l<��}����mx�g�ПP4BZ
��N����_�M����N�NY:��,ch�i�YC�g����|܈[e��O�V%�|P W�����u���/�}�{���O�ZQ(�~�%{;r�ȲQRɣQ�*cʩz�@�u�����o{i� <���,�ʯ�C/�I��3Ô��jL�Hø��
�Z[ �������k��`:	펺9�e�<�/r���i� �¼Г�8�} _h<a����Y�z<?_xSy��!�S���%�T~��gᕩ�^IS�>*�J��@�L�'�}����{ё��/]�=�V�)�	�ߝ�5H'YG�۵;C�9�TÌrz?���PX42P�NQ���Lw'NvEQw���&�kF-%����ڲquЧE�.|�h)��r�$.�K���*��e ��99s��
�����߶�~�^�|�>��L���l��ư��)��r#��V�χ��s�U�����B��Ҫk��P��,�P�U�b]Q+�b��T����ST�,r�V"'����Ѧ���顔��Mѐ�m��#;|��� �A�Y7vҦ�$��c��'A�T@�,��T)��_���2qҽrKg���n)�>�5��$��ܞ��.A{�'���S����8��a�0��1���d��6��]��_�}����@����Q���w���V��mom6�O1�z��IYe��<�������]��wӷ^��l�����3&0x�!����A�Uh��W��1�����"�L����t�4w4U�^���Fe$3GV����2����� �6�vּ���X�{ųN�^��ёt�)L7���7E���K/_�i�}�<���]{�EE�ׯeN�P[���t��4\/��8��6I�#P-+YS�
D�r�2Ag%3(σ|ҁD���Z�S�2�4f��˒%�G�(|��H�ɂ�
c~��#�t �ވg> µ�vd��z6E	��S�1��NC۴��3;��9�K�%�eR�Š���k�#��q��*�%W�k���O�28qV[6A!��i��~��T�X�^BZ֑�O���':�`�u��çry'�_�EB+� }�KT�WF<��Lp�������.]FVMu�h
�k1:6,J��6�O����Ň�=���|����d��S�)b��%� >�X�u��+x�C���6�4����>ʊB�
�p�pF�ک	Qa��M�������W���j[Zt�L���!�L>��C�i�]l��K[6`(�� Fw����l!��#�K��x+��5��	Pq�5P�����7~�37z��{?��)�]/_9���l�<���%�D����S(���NN�x���h��e���|ޝ�9��9��8��-z�r{����r���kʕ�%
��n�d��*��.#[�3;A�!��A�S>l�K@�)<���"4l��f%*Ϯ��a٠!z��]{��U{��=��#NO�0�F1�.����� -+�BnE�]��=���S�RD���43{���7�M$\�dc�" �w'����JD�V��QJ���"d]��e�����*?i\�1�S{��0�f�ct�\w�0z~���F�<�Tck��_�� �2������zDH�Y_r�� ����y��t�Rn}R"���;Ji�@�b)�5�� Q�:�ݍQ2z��)�H�3鬌yI�����A9Dzr.0�t�Xg�=7���b;ty��m{��{s�t��߽r^��u�u�G����Vڢ\|�� x����aR�r+�)G�%�iL(k8F����1��r����r&a��b�>���?�V��J���ݻp<��paܒ�5�
G>*�� �7��5��1�j4� Cc�g�;�P��NjGԃ�S�
8�w�i:��h�-h4��ɻ�,��K�G�作�(?]y���Q��c�"G�;mc�=F���������k?��J���#�h�p;nX�w���{��nv��iu�gm�{g`�)�G*�ֻ��}:q��m�RN�1��Oeyz���LY��2�E1���s*}�'�9�Ը�bF�qD�7�ad�t�AY�AcPY�+�!~3@�8
���z��#͚��,�j�CuҚq��_��Q���SɁ*[S��y��{�[��BÁ-���6�=����>�:���8 F� �>�����Ж�fJw���=��#��gGBmR�������ի��N��J��1xQ���r�#�LvF�:0��N��37��N?9�A��5�MU���ݫ�Y�R��.l�ô��F	�1��[?V���zQ�+��4դ�����ʃ(��<i}��t��������c�ru�~���������w�?o/_�C�;H�I����܃�K��v���9�: �����չ�j;�ᡄs�GF�O�l���@R��O�`�	��O��U��FV��ޅDr�]�����'���d>�Z6�s�27�:N�&�D�J�2W����綫nQo=��d��M�P�A��y$$|�������W���ؑ�N�� l53E�{�	���2��ָ�$xPv����l��l�҅�*[��+Wᯞ�{՗�Q�D�0]_��»6~n~��/,��������l[]Y�h��,��'����֮;�ۚ���i���fޡ�	R+0UMݹ�K����k��tN�+L2̊�8�Q��gff�-,��*(B=�;�і _[]m���)n���� �F�LC�QEb�j�Ȫ�?r@�F��F�!^a!"�g�u�P��S�Tw�*�*\�����]Y׿�XOT!��R����`��&�X�W�B`Q>1��Z�i�LC�S pG�Q�nD����5��LUSS�`�%��i{1f��tz��R��mqe��h���k�q|�ɡ�0�r6��3eS���@�ꗦ�)�,ˑ�����vp�����:0f�������v{�a��}�!�kNQ�Z�Ww8�ưJx3�79��c�_Aw�ٴNd.�0c�x���v��
82�QJ�j&_��V��z��!�A�����kZ�g\�$9�X�F�zO��2x�a)8��Y��C�ӫ������3�jG�b�+0g���&p҄�5�R����yƫ�	�|1�.?)`3�ĝ�lhG���Ҧg?��ɩ����F����%��V�T��b^1�eő^K�#6i��~Ҷ��;�V���*0�^�̆
ڭ��HVa
Y���|�{�'a��?W�X5���$�c�ާd���F�&a�!���/ezJ*����z�Jㄷ:Z�
]�0�A�a��a*ݼ'^ŏ�E)��#�-�pT\�wS2Ŀ�'O���[��+��(��y�G���#��CœL�r�R�^��)3��r�Ur��*�tV�L��dO�֕9r��h@�U	,3o��nX�.=K�������޶�?���}���~׾��Xis3Bw�xNYF(��Q���a��d�(�P��;{��)��+���p�;�_d����}u������W{h�����T�(��_��2yi��EB��}�~����81��]��NM���*e;8�͹���АpV�e�&]�3`�Nm7�3p[H�R��!r���K���V��T=�9u^�7�_}�7���k*�|"��w�#�m�$�(Av}�T}y�4�G�v��8+���#{�Q���k��|S8�m�cڍwvw�ۖ�[�����Շ�M�ӫ���۶��I;wN-i��ʽ8����t� m[:�ѵ9v�ntצоV����X��g�q'����v��+�J�QBZҌ��Y7#H��J֥�o����1��b�{�Y/|������M�����v��j��q�7e�F�a{��M���i�_�i�74L�(�$8vj����NhF%�C�#}�=F���g��U22��9.:�0��p�s�Rǖ-4>/�������q��!c�t�O�1����F>�S�g�c��	$�{ë�i��z���ܗ�-�SX�~m˨�,;�m�X6����A� �4^�h�Bz�Y���:�x��w4O�Q�{����Z�L0o�����xp	C��'�2X�_���r�{U]�M�C�u�y��:��aT~f������qya[d���[OMg	�v��pjÒs������v��m��:]0���=�\ef�u2:]�U)E{u�4��@��[�!�TE�El��)#�J�IDNu��)A����Q�ԝ����g����63喡��HxI�<$s��A�(�.�l�{XG�.蔋�3Ȟ?b�8���׏���)��ه���/e�)���㑝��@�$�0�4:D..0��E�EA���Б��ۓ�I�JN/�� Y����jz#k�g��2b�1=�U� =���@!�!5��I��O�ī��ͻL^HL07��@?pR&�mf�հ�	�K�ܳ&��"L����&����컙	�~kg�ml���ť#MӔg:����'nra���a���赳!��p���������ܣSi���iH��e4˲Y\u����Yr�C?�tPxH:ꜻ=H�d�C&F�pЄ[�R�&��?����f�r$c�J�ڒ���_@��������1��Gbu�I����]�xW��?<ɧV�-w�z�fB��v���*R4�����jܸ���U:2*5~)|�t�4f�â�0�c���ܥ[�("V&~ʟ��,l�Sǡ�y�F�ۃ�F�F�Z凾�6����-��sY�{U8x�?��_չ�{Y2M88Կ>'lg����{���(��M��{�ª?����t�:~��ԇM>�[N�R�f`�JgR���K�j*�odNb6hNgO�А�ގ4�Z�>WY׈����	rƩ>u�ώ��ɦ�RS�B�-2�R(�ZwvP�.G
��Qá�ٴ<�_�q����K<te��JN�wM�;�F~�ó��?��}��w�g/Q�qfD���O4��ݰ�u+�(�*�5b��Nq�@V��z��I������0E�4�t�]����"{)���c����u*���|Lå�s�g���*�ĻrD��$��#��{�5��+��F���o��ತ�(.Y�LY�L��2/åmLl�E�G�u|�w���x6Ւ���Z�	�=��ҧr	�d�^�P�&�O7y�>�6�������{�nqF`sg�;u��p��9?�����D����5�<���tfw�q��ݽ�_9�,){w�ƴ[�(�G��6>C�z�M�T}gJ;-��^�QA&�שN�s������PZ�6U��,t�)���a���D���O��	�a����z���.��G���ng�����(��޽�О~�}{�n�t>����4����Hg=k�'i�g��)P��e�N�K�uu����[��[q0��3����c�:�����2o?䟼x���{�*ÊC�ϓ<��LO�2��<A�H�\�
�	�!`��a�Q���1�H>#[�7�*��O�>�8)~(�VVh7Lf��D����$};Lm�]7fGT`6���l"���c�H1�*�!���Ū���_��Me��;/�#�͇�ħki��\4b���3���|[t���
��:���NegϵՕ�����?��Y�ۇ��Y��u��+1lUZ�2�� ���ˢHr� >HY���9�F�*��v~���%�=������f�]xn/�|�Y���eA�s9'���0�o�
7SB�.��<����?�,�ګ��E�h��R ncX�nT������"K�����I&�.\��1�����Hc��  +3�a7]�LbO�s匄wIHa�O�S�wH(�m�lL3�of"�H�wJ"6V����/ӛ��(%B��s�>=�
Z"����_`�S�yi��i8�^�x�);�C\�GI�F�����5����k(a�1��ux|��r�v�ak�ÅO���]X��7wq���)B���[�c	&��)F���4�p�Q��0�`uZ^�f��ާ� \d#�X�<��b~�[� ��:0���u�D�HЀ���P�]}�f�5"G0���ٺȃ��ҟ�����.\>�]��g�&M��4��ݼ��3Iu� ���#p�xP1q�Q��NN9�ꖻ��\^zf��E;���1�jͨ�_���z��C�@`X{�ԡ�(ǘD�HCc�s^��n��������<Z�.ڇ���!ge��h��A�Ұ�}:�_��K����0��O�[�`\.�%��K��)��3n���Y���>�<w���?����w����A�Q`����p�T}/��	k�r��8�Y�6!.Đ�i'���4�܍.J��?�g�T�t�+3����t��#7P���1�D8�G��% ��_�y�FiX�M��Q�wpi[��:���#O��-�w�ً��o�}�~x�T�����N;�w���$�tF��Vޡ�+ϱ>e��L>�vR��������W*�JH ֘���K�Q�J��}]��������3�O�d���_��^�4&�ю�?:6��L�wsQ�U8i�'�>IC��C����*�3�{߯N�LYqQ)��4��K1�_dI���J���I�����R)�W��n�{�,��K^��cG!%"-�Q�UQu�����
A���\��F�]��?�5�*��u{��7(��Zٙ#��y��I��/�g�}�>��ݺu;��Ȫ�����5�vZ��W�O:�(��J�U�i�s5�)�S ڕ������n�� ���d9��!�v���0ƃ�����svX:j�Kqk���fq�z�߲>�0�w�����h�"`�?�	g��QAt�Q����������'��Ź���:I����/ߴ�0��v�����'�/� GQ�؀W��Z��yߩMX��3W��*�c���	�rWJ�!!�P�7٘�td5�'�>� �#^h���F��R�4��!D��n�:K~{�W�=�3�ƭ���n4�1:%����0��(!�i�����V�oҲM��H����k���;������t�(���J�vj���8�Ԃ�V㠹�S��r��<ß�"�������K�����ϕ�r�R����X֑�H�1��Sg<���ŵ�~�3|��OD�r߃�����@X۫Y��ocd�5���?���׆J��"N ���<11��3�%*�9K:�Q�r��F�$���*��w��v��:�^z��Gih�=�6=	0��)�Ư2΍
������E�����Eod�졔kd�g���%
� ���սG`�u7�C㋥�����Uo����?=ӳ"#�i�hDr�D��2jt��+0
7Eإx��%$�GV+�TJ���;^�����S�NQH\�znP@��^b�.N^�|m���r⧱d�]k��y��xC:�hY��4ȜV�W8��T���zI�PO���Ը��#<&��T ���u���a�quy�v�n�:�2C�a�ꕒa���W��;�p��f�0���\��L�5OY�
|�IA���-�����������O���-�tNJorr�1 4~-xL���#��F�ʔ)7�vM7P}Ёc�� '�3��˙\�Lv�3����3��o�����$n^:�ܸ�\��A��Lq��B>(��/��B#ŵ?�
X���`B^�#ϸ�N���ℷ�P1�(���4!�ʖ���v�֝(1��btI�g��⼵mO�2�zp�]��>}��S�I�}/٠�Q8����K|�ٽux>�n�D��²(5\�Ϣ��c�2���A�����A�p�ze�
��j������D'����,㨏cˍ?����-�4��{����7J�U��t�L���͏t�}�;Ǯ�G����5�sjag|�Q�|��aw&�ǔxwjU��<$L�?��1	.�&w�"Cwj�#P�-��y��=�}����7O۷��О���Ӷrв���(
)��#V�Ϻ�n���|����o���5��J���!AyhO�GުH(�;E���&j�W���)�Q��l*�
'����vki��_�2���ʙ�J%Tyey�Q�9|G^�{/���Pw�OZ��4���,W��K{��R_�P�|�7��-�N>I�we>24��T;�OE��?qa^^������W�v&��r&Մ; b��N�|S�FI���©YZ� �2\ՍKU�-S�V�3���Gq��6��.<���ՙn߾���Ͼh�?��thR�XvJ+�4n�w���/��`�4؝Q�t�Q�3E�'v@P&q0<4E�q�~bdMz�k{G�v�q<N"��M�5��C�M�֩�f�k:��;�C��B^_b`] �7�~�KGU�c��4h*(�[��������gO�O���k�͹-���$�v�ڛ����F���j�D�e��GB�)Q�_�����r�s�\șq�p�&h͸����7p��vN����GY�����5k��dII���<�O^��/_�o��8������NQ�WmO�W>�z��w서�t�t���LAN���� ���_��֟ƕ0���5äpX<SƖ�)x������6�T�Kgda�����b�Lų̃-��.�"�B�х�ͽ`韭�z�'�-m���	
��Q؄�����ƤtgܒQ�!M ������n�v'�ce�[{���]���V�_I�5f�����d��������z,G5\�a&5�"��"YVde1�Q +��Q�D@8��&�@��J� �����O#d$�r���₨����L_b�J��cdY��m>�B�>�6�5����|�`d�[�.G#+���B&����eȃW��r�=Wj�������ܙT��K���H%S� " X�3�S5�𓰈=<T��
����K��z�$f	Ⱥ*b
8d��0u�{������"�����{��m��uG(���	B�TK�̴H��y)#� ˠ��%���*�a"D9��`�K�tQ�9����;u:��đe~������xדI�J�F�;���i��ο� �	����Oa��.4��u'F�JUz�T,:劲���Ĥ;+�{W��4<3��^;���$��'-�T����bZJ"�Wp��_ē��OЅ.�nD�fC�8a4q�A#ˑ�ж4M=tkU�#���^��I9��H_���z֛��r�K�W����J�*и+$�/���b�F�������څ4��ڰOA�f�RR�ƤI�Y�N�8):�� �f�!�д� �C�*������޽��u�-",�Y*�NUt������f;��@Y&�6��9��S��kh����T�=�I$rN�4��g�Żᕱ�e�x�������_ڑ6�^�<��p�[�d={�?�5H�0]8�a����/�|�F�w��XҜ�<�����SF�ve=�߻?ߔ'���#G={�����h{v]O��<��QL;���`6�@�|���7u��:ȼ�:���ـ�{fo 'bP�vy����o�}x��3�^aL}�-����i��[�g���7�ݻ���{��%�Զ>U,z�O΄�+˒�v/��Ǜ��5����pVQ�j��چ_!�0䔯�N�˪=���fS�!�|!���є|iu��%��x��28�c***p*��J�_ַY�<W�=JͷR�1�R�*]�C='���N��/��J��Ҝ�Vʓ��Wh�<��H�Aw���R|� ��'m�
'p���QMd��:�<:t!=d��q����I�j���_߁!=�d��  !��saa�=|��=z�����X��͛7��۷Ƚ�L!������_��>z�u�N�����t=u+�kк�}#�M/4v,�p����;
��灅vP��`�e&A`�$������1�Dv�����.6=S!k,�<�+���w��g�-��s>�ߡ�lw��y�uiB+��gȏ{�R*ހF���������>k?��gmqv��5��u�ov�v۫�2%w<�g$����a��TLϳ�(�냓ɋ:)c���n3ʦ�����Xh��䫡�L��u4�}�X)'q<y�|l��Yt䘼^Gީ�c��%5����<6�~�\��v��2�{.ڒW�
�~U#���e9�gG��sJW���[�q�@ݹ�u����Z�tHt3��z�q�e=��l��?K�C��!�c\�S�~"Sݨ��d���]*�Q^�߲&��R�mRF�dE'��	��|q7�5כN*T}7��.�az?�VuT_)��s�]���,�n�m�kGG'�ɆYw�ܤ�)��1Fֿ��=-ޓ��2�@(�fCM�P8fؕ��AZ�S*X,u��CE�pVFh*��ݩK�Ӛ?G�9�������>��I��Q������ʬV"NV�D;5>Dz��uyXɢ����1&���S&7��v���,2FFA؄�h��F"�����;z�ӫÿ�yW8��� �|�DT���%���Ȳ�S�8�ɞƪ�Q��DlE�G�@ԻB�rK����&Di����=�.�>DY����;�"|T*�����ptr��E��1���K���sz�A���_
+�X�ՕK��@��LQ�����2^z��1㚛-KF�����N��zn�Z�<pZ#���=����8w��ۭ�����ڍ�g'�;�dd6�I?�[����ۤ;�5!d���^�ld ~��zZM���:����ோbi��~t�����fU 9���ȧ�r������!�gyod�������48����a����M�w�|��T�+�4��s� @�S4( W���O�)�i�,�S�t`��մ�ť��*�ehY�6d**�tEA2%
nC��\�|��apҟtf�:!�G3-��rgdy�ʋ��Bhz�n����o�>ʌ
5�2yY^�<a�7�����	I���'��3҅yE	��y���ݽ�w$<�OC�wy%yq�F����>y�����^m�k,%.��OA*\�|]�������4]��X՟Pq�F�t]��C^i�#��4��_�P��S�Bˤ��D3\Nſ\�6m�����?�c�����ٍ�����i}[�������{�?��>`@}@Y���F��9m�ͫ�Y����ٳ��勜y��n���={�2�_�6��B4�<�6�wcd��M��6n����:2�\9�?{�Je�SL�]��)�r�w9T~�X��#�����g�%�"��%��	�A�:�3�;m�#5Vh?��)���Q2;G[?1C���/�E��d�55�7�h��}�MO����IL`��7�(��NOCy���5�m�m)�J��P�03�W��Kd�x�P,��E�S�  �k(�DCAgcv�	��kG=�V#F<ͅI0[��#|��e�Ƽ!�L����ԓo\c���c�����"��Y�,���'ݾ�9X�e$kmm-�������7�f�a���Hz�֦_ /S�ST"%�wt״{��ds2RY�M�����	p%����m08_��ᑣ4gQ���g�>l��Yz]B�<����ᙛ��jy�Qa}P�v��4��#�v�`v~.4ggZ�;��]�����[+�g?����O�>��C���O�6:��g������vx��i���hp�Q�&v�e�p�(�	~ �躄��5�4t4�=GCK�����%�/�)22wB�k�%�,�ou Hnҽ4�N�F�5�)����)wt�AQ��1�>�w�k\���ai�ͣ��7M^�=�x:>���11	�ܿ۞<~�n�Z��x|���v�ch�@ҝ:�SPm�/�m�r�vI�-�$�p�3���#��;�0����ö\���D�.�"(xו�Ui�L�|xOX]�y�z.w�*�v*rbpU"�lW�Ӟ�OJ<믱뚫���������l���7���0��*x��݌de���G���?��������6ĸ�A��a�A�,
+�iï�-��<LM#9��Y�"m Th����g6]^xV�߮���J���O�O�����Ob-&��N�K�F�<��8SMy�{����p������8n����mWm���=��Ȟ>{m���!�V$�^���(��?yz]W*_}&+��\$|9�д���<	�Tf�i���s��+�ѐu�2��#�^pL|Ó�#�e1}�#P��K��{^�B��%��ڢ�wz(F�w��)3Ntڀ#_N�?����z�uM�yrS��a�83�@-N͑��S�YVi㉩��ڨ�sa�o��x��0�"'������.�c�a(u���4�N1��.t�`v���s���5qr��w�%e�ʢX{H��@c
�L�E�Sg`|�ا�N��On�������.���H����`���40�ʠՑ�B7֧�e�U��z*Lr�ϸv,�lH�G�zHt�(tEk8����U�L�a��ǵ�za� d査4ҹN�*��p}Z���Y��9��r�<xt��PdW.u��^h�����)0��Agy���)D�JvL�n��=���(l?X6�**���=��!��nO�b�Ӟ-4q���և��ͫL��`Zy�?\����Z5���Oy�ݺ�s�_�#���y������J/#�ٲ�mç$�j��J�S����l G{!kx�eK�;LB���*��n:2b��T[��Jx��DإM0FMy� "i[F�k$ف�s!藍��T�!�.�Z{���z�(,"}��� #y���-ᆲ��[U{>���U.�r��&�wE�������eL�x���=��sϞ����z�����m{�������A��v
�� �.��g���]�.��^w���.�8�*eo�Ӂ��~l0�0��)�ȐgXz,��:�P���6f���;��e�)'l'T�3�:��0wJ���,�Y9�3��C¦C���R	�J�IH҆�z��{�c#�U�:�L���#���]���Iځ�!����a�@Yp��РS�RL��̬�:���-MJߣ8���3�.���f&���,��Ɍ2�?��p����6d#�������Jl7Gs�K�!�����JeAJw����(�����r彅��v�ν�~�6���=rktg�g��c�a�#1�T8z��h��ͯ�ӧ�b�:,��/0�?��#QZR;�D�A^R/r$�g�u��0������,��_n�>A�:��*zR�MaD/ͯ����v"k�v�����s#G��7���u�L��:�E�]��'�U�!�=�s��C�����Se��i�NP���W���y��{mw�i@}ȵ��_���>|m;��y譵3u\�9>2і�pˡWGOQ"4��V��
Z�҂t6?��x��>�w�Ecg�:s
���Ϊ��yhz�v�e�$����7tYK��K�H��oSm�+��k$i��+�T!EH@~8��}HZ�m�y	���L�s�+�95R�=:lK��㇏���>z���ww3k��e��ٓ���3�s-���C�:��Z~!��������'=Z�+�����%}�d���$R�T
ġ�{v�������q�VD��tm�;|ɣ��vA�����J��Gi�8�i��U.��Q_�s��ν�ڝ��Eg���;�3��m�:x�Ν������v�БLg)
&]S���J	� q#1��_����<[*0
E�@�v��d..��q�["�d׺�H�!וѢ��V�)��˫`������;7������w��=s�1�gݫ�}��@������˨:åg�
uc7X��ɍ$�:d���T$Ư�bV+���|��g�G(������7����3}�{��|�^�H�y��޽�l�]����ۍ��p3�����׍x��t ���! ��J�֓=j6�s�% ��\�23����r{�ff"n1_�$�`zY�R���;�ã*�ԿJ8�����]���Py��{������t�0/L`o�����P���4\��h���NU<���C+ӷ�|����'�"����s�%��s��̰���X2>�eZ�u��7�O�?�׮K�{�}� *?C߼�/ɻ�?1~3|}��x�>� �~�S*��_p��dM���,�����\+�+�ou��k�T��A���we��b\�Q�מIx�B�8�$�-?��"���?1��낊���LF��g?�W�i��xMgV���|"3�W#A7�v�t��i��q3��`X3��'��WW=$-�ƽG�W�����O�=N�J���~�-i��]ځ�w��|+����C��{��|S6��S�ʮ�w(��B7���7ߵ�������~��}�������_�M�կ����W��������/��������Qv=����r���c/��n�����tn��t����SY'��.��r�n<�M8��򤜖\S?*	ٴ���Zi(cd{��SW�_a�9
yU
s���g��͛g�!�����C���$��32D� �J�i�G#�}�u~�NE��Aa��o�Re�kx���0����3�	8q=��a�4}V1͋G���3F'��w�jz��Ʉ;9
�*k�rh����ˉ����s>�~�%|���=[*����ى�n������������}��Wل�!�\}��7�o��1���!�N�MG�m����8;^n��eDҜŖpQ���~��)k����IDW��i�v��-�S*w6��m�-�Fi����5ț����1L�:Kx�K�pƳNQq����b�qͻ���ꜙ����=�q|�4�5�(���4�xv�b��/�������;��m�C�h0f�V�h iI�6�]Cҩ�N'ՙ�g��ay�p�m�2>�'ǆ0
G�M�(*F�z7�<	���0ZP�J�#a�QW���F��NC�������?�8k�<`���W7Cgs|gM�2B�Y�]�>�	��5@�����<Q��l���llÿ�y���7�۳��'rGN��<(Z(��~�9ַ�G�]�eNq�Z�������_�=��A#_�CknD���e	����$76�i;6ڦ#���9���(�_����D����"|�p�'�����^�\�P���,�܈'#N�|vX��c�����;X�
��M��e&����:� �y��Ue��WH�Qp�w��g��w�2�p�~�¯ǋ�q�Uj����1HШ�cd��OC��f��)�Z�UO����4��Q3�jР��z�%��B�m�7�0��y��k��ڇ����S;/�1�w���������C�t��CGh����Ѝ	읲G�h"�V��ϵ�%O�.7�0kv���oZ���&U�f]e��Y�������#���v�-�b��;�ӂT����@��pd��n}rG�eJ$�۞�i�1�2�5a8uŞa�)t$����~��]52}���\F����K.i�sծ��ݟ��3x�G��MDtߒR�|�o��#~|�.�/�ūB�Q�ho�%�r�DA<^�A	��!*N��@����4�t�:���K^�쪲���jZٌ�;���7�a=�����kϠَ0��	�Vy����䝻W�����k l��I<����r�4���U���)n*�2��+�'߂�ŤOZ�g㙰�o9:8t)��K�7v��x��N�:�.]Ջ�}=G��?�7>�$=�.g�]ڹ���-�JFu΄����S!���I���GA #w���ms[�����m����0�^��j/_oƽz��^����N{�a����u��<Bfz�i���:,�Ѭ+4;�I/#�Q9�r�(��/r��Z̺*��@ed��e'\M�ꜳ�gZpF��>!�(�<�um>�[i�^p7=G.r�!�vd9��c/L��!kDiT�C�2�)�������L�h���}�3�</}���ؚ��f���S׉��so�i��a���`��]���g��,��h�8�?��0�>��9�州���r�)���D�x�Fw�LÅ���\Es���;i�g���ّ'GL����w�ݽ{�}�q��'�d��4�����7�������?<m�;��a�LuZc<`d�~Ϳ⎺��4(x�;[�g`�
���	|y�_Z�Һ�B3ⶣ���k8��P9 V��H���GM��h��}���j2�Dݔ��K���w�7���C�ֻ~���l��ӳvX���:x���\��yq����r#�(�5�$��)��s��1\�XjKW��ը��� f\�/G>�z/\fs�Fث��vz��1��.��I���H{����NZ�;�~335֖����L֙M��-C�A|�$�K�pD�ul�WX:��i�N������uhG������jV_\\j���O>m�y{���v�ޣl�07��.>_����G1�<�*S*���~�;�+��N��ru��)�:��0��NS5�-�.�s���t�
�/�1��D�(�<�:�Iv�ȻD��=���w���$��쬰~��ǹ�)�;�G]f�@{.O��d�$~�j�`���Z���N��mnvX�3�as�%V�э�?�Q^�����>�g���ŋ�fl��9>A�!� �4|V�w�s�*V1�d�^$`���0�w"�\ߢ"��X(�yK�N|������O��{w!�J��
c���y���B�P�U����. ذnY�� �]``8U��F����{f
i��UCa�dCPMN��)�H.K�%�s�����n��/��������� Ҽ�l8�{ J ��Ɗ��G�'AQ)`2��^E"\��k':����r.W�ш�1�=w���i�����,��Ų��ld�,(F:�|�8�,  D'�B��K�YHl/)�V6]��*Z��qʕ�':	��;�t�4�Lu8C�q��s`���CK�5�A��+G���uN���%��Mp8c�M���y�3��#�,�|�C�����K�q2��fS�4V��nx���IHPD]Z�T,	W��{m���������p�Ϭ���{�xֿ�^�+m��J�%<���?���8���OeR��`7#�^�1� J�#l�iG����N%�C��W��t
���J�Ѝ�9�<w(�뽫����m)�2��K>��xW�r�J��{�ښk��fӠ����/ڳ~��z���iS��_�/8Nb<w�]C�W�ED ����'��^��2,&B/O�Stx�z�*�1���x�鍡��_���q��(N�bZ�ۄ�*9T
����TyzC�2DV�$���,^׉��ۿ��;p��!I3��r��V�+�Uv��>�7~7xQ���|�cQ���\F�/T�Z�I�]+[:����	�x��i����:@��#-��+�Q6gJ$�9���܋�vx�~��L<�Evp�w�'���4����y�]��R
W��7����]��~;�j��ګ� ������	�g
bD	[6]������}d�x^����A]AC���4Ӌ�FX��-��%���o���@��pZ�r�)е��(ū����";V<7����k*c�gz��	�pDD2=��)^\Ǜ5���I�H��Ćm���˪���K����6<��V�P1_�4�4�����ߴgϞe��rQ9�����|�q���ҕO*���� �ވ�3�5%�I�����2�N�4@��Nk}rՍ<o;-�3�RYN�׃�쓞[�S�����&�"ێR�&"�b���wJ�߭�6��a�����=����]���X��a���l����ؼ��)7rm�F7q����x[X�m�+�m~��|�m�o�,�)�z�����X�sS��JXU����N���F/+ˋmaqc��w��y��xҀRo��s��Ѱ	ڼ�Z����Yj�o��{wo�;�����<F��'nw���|,��v7����Nq_]Y�fM��_�[N��N�O�3)mr昻T~�����{��(��G��F�����G!ŭu-���T�S��et13�~v�h|#�����t��,����<&�@cZ�Yt��o��_8"����8ɣk�9ŷt�»�O����7s]�u_�4]�ﮝ�K+m=@�,;e�<����Ch�����}�n{��a�s�68��n�h���/��/^�z�^���q�)�f���S��F��0(;٥M��}�:Pp��(�-�x嚆c������\v����Ĺ `��\�����i��q��#.F���A�*�i�QF��\��(ܗm����b\mo���s����b�� )T��"�0ǫ�[���W��{���Sv[��Q�z�D��(�U^�ͫ~{%0J�@2���D�xK��r9O��7�ɻ��r��ۘ_��O�Ȯ�K|h\Y����5�гAD����I�����	
2]�9�<�Aa�0�cc���:=5�����!��G9]�w@�p��v�q�,g���p�V���P��pb/#Pi(�O�#�9o�Թk��5N�1��;�i\�XW�wYS�*����h�{3�3�	�GV:������T��N����U��SIy�W_<����uwk*�� ��j����KN��^;�z�����4�І ��>��-?���5x�!e�!���^���ɿ.�7?ס��*�`,u���Z]�TF�B����J��g�%]/n�xé�T�i4[9�o�N�����R�M �@V��-X5���TW�p����}׾�����ݻ4HI��$�º#ҕv׸�oq	�����p�o��.�����I)yJ��`��'�ރ{��ǳ�7i��0Uڕ�y��2�,�tiя�_�\��r�@��{�����b��dg��ӷ`�S���&-�ﾬ\������N\]�>a��t����K<YO������s�,+��Z�u�iTu��L��\�Pe'�jd)S͋&`ĕ "���#\��L�2��)�q�o	#�ƥ,i��6L4UZ)�w�V�^�.��Kٽ'���L5�R�#3]���3�&G���4�4l�j!+U�ٲ��k��QI�/�U����ƻʙʝuc'nFb='�|���SZv�MM��50�����ҋ_��p%�t)<�|P���]��:�)��]��Ub�����&�8ů�����g�������Z����WF��T��G[J��.���9�ύV��{���|��������W�m�MCe��S���h�����Vǌ�[r�©"�S���HΤ��	����ư�-����9�C�X��cU�k�A�H�#ԙ�9]K�9kE�_�����PpwG�%�k��|���>y�)el�5z� xD��X�@Z]] 6��i�$�Qpm�G�pݜ���r�s�v{�������Çwۣ���#���z��n0��f&1^'c̭-/�|�}g���/�U�]�d�Օ�v�t?��Q���/�g�=i�o��pZ�����h��9���-�϶����ڧ�>i?�ɗ�O���g?q�q�����o{�Iw��AKĿ{{w�|� ���O�W_~�>��K��(��͢�Ўf��w-��������s,�]s͟u$�X�Z�5=X\�8��)������%]]IWY��y�A�/�ʏ�2ꭌ�Oc��2����-Ƶ�#���Ԙ�l��#_�ZKj�U���>N#MW�.l�g8`��
�uf�Ԥ��T��v,�/a䮶��լ�t�q��z{wD>�����8K���r�7���>�Ud͡����/��ݟ�u���y�~x��v�h-\y9!�����¼QLPG�����B�Eۑ��
� ��a�4�ȴc�SQrU�]ܾ���B��A����vbY^^�N��t��<�q��^�߃��xii�ݺ����Zh8`�y��ٞ����w�ڛ����Q���a���a{��}��k��*�Xʗ�1B�yg�ĠI�BV�(JkڢR�*o=#�Sf���"suq�_��C�\��FK!�����("�t�`��fA~�Ώw�gI�j~o�8IpCT���J���<yߘ~�h�_�ڊ�0�4J�ò 0C�!QE3J.��Nw�$��]��!�A�r:��BO�m=�-̴���MYC8,#�f�eF��F���ݵ,�%�Od�=(S�niH�֎^4*�ry��;
5�s$�5|�Ũ'Ώ"|���^k����{��l����!ʀg��O������ڴ�,���%WG�T$dȡ��61=�&1ǸѰ8��z��D�q}8Jj\��`�b����H����4"��^(���P+/��(	�>G2�9���Ж�5⦟��
��x�
-�띫h��7]k�*��޽����ċ0�U0h5 qu�Co(DQl��O)�e��i]���&Ǉ��1hb2��n�k'��	mo;�tҐx���%�t��;����c�訷�)?�S���*P�h�#�N_u��W?�Y��p+Vq�����������/~�޼yENaEՌ2"*fUf�I�=�g��U� 5p�NϜ�!E|�y��K՗8vږu.U�T�3ZG�>��[���F����ec�k�e���̋<{Ó�w�2?��M\��!���_���*�/y�gQ��;�ɦc ~8���G� Y�<�'����b ��c � ޴��e+z�ܨ��@J�]z��.߄M�WY�4��~2�<&�W�5q�l�H�z�i��3�w���OD	qq�P7�%ޥ�.?$՚�\Y�y�E���^<����1����h���H3m�7�І4C:=-%���2�_��s�'m�����NHO�nq_J�!] Ӕ�����ށ��W�㤥��873��֥�Vv�C�񰼬v�Q�*ez��GܔS��Km�]eQfҭ��J��I.���G�R��d6M;ԁ�uq��A���2r���rđwD=gv:�쬍B|��
�9%^ģ���&k٣n��Q�Nuw�f�8�	�Wd�F<��h���m��n:qh��W���s���L;<�ʆg���G&�14<	���"�!u��63�E�N�=Gʀezc�T�������1�)[��i�Q*���\��e�u`ҩ��5N<�Ђv��7�(c��@�:��3��t�;+s�g?�����럶�>�ظ��f�C�������/��h;;�u:ʴ���L��o�n��^1͈/��wwFw�#�]��w;���(�:|j����q���ťL)S��x���ɚ�����5�B���˸���Pi �k��-���������v͞�`e`�(�n�3وÍ��)��nj�N�o^���3&=GS��}k�=���쁰��D\ef��w���7/1��`�?�.��[oѧv(+��L���AYY�Dnp��Q�����V���k��#j==J+�񍛙��N�5���Fr����#�:��i�2^��{��G;-]ɑቒS�#�kL�a�l�)t��,w�[�S�n��E������v�ӎ��Sb���;��G�`��-�S�]�F�_�Ȃ�����T;�0W*�E�(Ced�e�sv�Y�J|�da[H
	 2��G�����;����_~ھ�=��^�{ûNgxXA��v ���^��߾F)����ѽ�ѣ���,�9,fxW��x�^F� ��>�ng=jO�﷧/���Gm�Q1�)���/=�b��QN��R�,Gj-t	��'��ĩP@���B'�Mh�+L?��������"�]�(:�d��qw�.~�>nW�*��jh� ajd)�F���۹�ed�Se�-�s3H�!,�S�)}��m,~���<��rw�V��@\b�ȶ����lF&�V��!��6;KE�X����!���itm�C����=k�v�R�v�rv��,�$�l��)u���?���w�0��lf�D1�=^*�ZN������V��S7��a�615��1�Fa�+���(��Q��p7�l���*]���Ti��w����m���u�O�;qg�M���@*$���+E�7�����ԍ{�y^�8��LE�x'�gR(~�v^���{e�:4��x��S�˕BT��F����c�d�ny�Kq`oϤ�#N����܎)hS�<9ޣ��n[�[1��#+ u��U�9�2�.��r�x3\�ߩ4� ���N�(n����'O�����Obd�,�QWV���c�,���ܶ�4cP�4�f)-�%���g�{��2��y���'�p�ow�o���R�������O��$3�Q�3]{5��_�%�44�aĩЈ?�L� �^~��ß����^~�Y6rB~wJ����]yzg$� �+��z����+߭�"�x+Hťt��1c˛�#͊gL5��������\�v�7.aKR����Ti۰�c�q�u����O����e��q=:z#�(^Bj8�C�7��
�������;!�[ꢫ�j�;�U~�|�lؤ�_��� >�� :(��������)_��'W���aC�(U=�����Ӻm^��\E{��>?�w�*9%�W�+`-���Q:�ݲ��,��G�S3�p(Z��z��;v$c��<�Rxh��;ιk`9e������L�]�����.�W�q7FwJ�`���m��qQE�Mw<��z�#�2r�Qv˔�&�|p����ʹk��b��ԑUQ6��jD�#k~��it%��c�Y;	�zG�#3l�&��F(��� ��iS5��'i+�Y��L��]��<��g�HB��!'���#�F��3N�wɂ�(��N��3������ۧ��o��|�~����٧1>����347޿k[���Nٛ����uD6�s�:-��
����g�i���7X����)�/uGs��7#8Nw�N�[�8ګc�h���ꨐ��%/ʯ�f�L��S��m�%	�wch�����&�C������d�鴞uv��X����o;Ur��z1�)t:�y��(���oS�_֕3�hk�7��wI�>g�}����?���(��	_P!�_�ᴣ�І�8�&��<C|zNV�;�wu��-���Ҩm�9�C]��H�Pg�.ț�q�Ç6�4ҥw�	�r)��BHW�v�5;킳~��i�� I0��L!I�iK��ʻkf�A�'f�P;����$�mu=xy��Y�7F�N|��}{�&���<2��qGX�����-.s�ӭ����p�Xn"�˻J���֬�����}��� oC �t�j8ĿCe��w��C����tA�L��,�e�]Q��+��@�[s驟L!�?�t���Ӷ��u� ��cdXp5m
���L��?�~\�J;��Յ���}�{]�a$�z��N�_��&�I7=�6Z�+j�/|�Z&%|Ot��-�]�*�
#�����k�ɆQg�&c��;4Ous�a�.⡿nx�&S^���d��Q�aMF�,
i��L�j�B�嶠�S����s�E�����)�kj�e�^����v��vxp�P���jt�]l��y�
�n%ﰸSJ���16:#+nbCC���"�e�
�N�E��9,����R.�럾z�'V��3��o��Ɉ�8��z(5��Գ9�����w�r��s�K~�$r�>�NpU���.L�/��5W9�%���#�U��W����4-|��kѣ2,�Oy�s�z��봜#t�W�7 ƴ���Y��D���<N= �v<�U<Rq4Z�󋛳,��fz���md\��yI{����@=S|�&�{�X呺�^ ��7�I���TXc�C/���<�ʧ~���6`��a�JSe"Yqy��,�E!.Ϣ�7y�V�K�]��^L�2o",�	�+Ʀ��k�U��_x�{���R�M?.A�c7������p;��p��#���̳����Ʃ e������(;	�y5���<�^�z��K�L�v�N�RV�p�~��;�S"D*X��#)P����Ea�qEG��A��˂K��6?o�$�ş��Q�Ы��R�����|��IG?��-�64cT�e=�u\�'�|�ē�4�t_�S(����i��U>��q���� 5��+!���^�� ��L�Buz�����xҳ�H�w��jȇ��/�&�&7����ty�k�l���$kE��G��+�dvD�J�24�&�=�]�3�a�6�ۣ����������!�H�3L�.�2�\#&�Y���aƋ+�Nё��D*�����M�ܰ�d���`�wM���F��L=X�%�K��Ļy���R�hk��bE�aݐ*i�F��4��+L�:<�;ީu��#��U�@'ԁ�e���J���r�¥�N^k���.1��xfv�o�m�2�M�����4J4ǒ#9HΘo3��rf��|[Z^h+n�W�:�o���*�|sf�*���`�.��z��U��:���Y��w�ޭԫg0�VVWR���1�5�Gǭ���&�/��wV��{�������x����j|��/:��t;e�8F���r&��ȗk�t��mN��_��Y���xG���<fZ�N49i>�U�њ����I�����oS�|��F��ML௑�R��^83��(e'��]Ù#F0�n0�KN���� ��	�[xQ~t���3k�0�W� t�'�NN(ץi]m�#ܺZ2�����3�����\�a;�5�g���J�[��>h�<j�����kK𣆮Sx�`�i�35ꈻF��7ڻ���d� y�����ꄌ�[��$�3m�L$��9�C%F�E�?���\��p���G!�� �	��G'mk{��z��}��7�w��C{��-�d��ݻ.�P�W��K~�Q H�
�C�霌d
���i��=ˮO�K\V6�荬�n�!9�m�r�Wʫ����n
�z�e��[��p�[~!k�x�p�o�pN���-a�6����:��P��]y��K�n^sEYT�*���w�o��
7�����*�1�g����>a�,\��^O{2T�u�+�xa�i��@ѵ��(=����a�./���4�.�<w������F�a\����+V�x�Ѓ�a��4
a�	}t�鈝�E�.^���YN��������.�w�HC����EIY����t�C�(M\�R^�����C��FO�
�����/W�?�Y��7�.��ԗ|��Dr<	T��%?���2ͮ׊_B��tN��V��S#�S��V�^�Zd��T����&�W��W���u�oj�_�U@��\��d#�D���������iu
���tly�f��1˟�잓����i]��O��ϳ>�+�$�~E#�\�����+�$H޽2u���O�q�W}����/P�1�rWnW��)x2Z�3��+<
OM�"A��DyJ���_5�2˃[��'D��y3�w��q�iY��R'?��/��9Gy�i�ȢZ�c�B{�=0��xi��wϽ_�����W���r6�\jCʭ�n}PW���K$�~�%�>t�g�_��VrFA���t��+t@|�H<�^�+�*\��7���)?�=0��pyλaBbN߽���L�J��KT�@;��6��'F��'�IzWɗ�{���{E�8����='դ_��QQpm����)�	�C�?5�X?r�>x�Y�sy�6�W<��е��hT�	�҆!����Vd�|b8��!Y���>���v��������F;N��:e���I�N9eۛ�����(��b}{�]��Z$��;f��D�Ri#�Q�R�-;���A�S�h\�x�f��n��q���P6��qA�q�X7�ig{��ۺpʜ���c��p�q��F��g�/qַ���N)_C|��n�Ri�8���U���e����wÌb��Am����e����4a�5��1��;�}zf�ͺtb�)�v�bH�^9�3���IWҏ�I��A�mġ-�~=��z ���O�C7��q�r;�/����9��<����ؙ��Ø~�DTpV�r���=Z�?�H:��sT��B?v�Q����+m	�5Xas�kaa)nye���i�k��ާ0@4��29�!2O��9Ϙ�&�g���*��Ḋ[ɳk�&1�4�zy�Ƞq�xb��z�z��DiZZ-� �����Z�N�W�X�k����&&1
1�&1�4u����Q���B��5��w��:w�WV׳f�Fͭi���)�	  ��IDATL��� ��g�ÿ��+����1�Pp���Bj�J�F�?���D��,�f������Hs��Qa
�L��"����.�޽ݖB�{{mg�!�W���߶o��}����p�4|�޽�+~m}�-�k�X�r)V;�@��0wt��}2\F���<��y��V��$Df�@ˏe��ս�B�%x����l�ޯJjy�u����/r���:� �K9���[�����g��`Jp}S���.�
�� %��Q����J�A�:wN�	7���c��Y�x��Y�j��F�(8�������ҵ3��h`��$[� ưGL�Z�!6rvZ'���J!}y9-^`d����Q;��:=Q��d|��:"=o�@~%hۛ���0�[��LG�+�l�s����"n,���P���~u�#�o�?��A�w))wn1�(���'ϩ.>枰����o��wWh���k~�ʻ��h.���<n$���;C��L
���2\�%��ˊӅ!�kZ4A�xG$-�jh�kR)9W��~��L���
V�2�4�2%�3myû�̦�!uu��D^�e�tn���z��򳼲BC3p��;z6M�K�*�ֽI�̲W.*?��?��/5�#`�{�j��t����>�/�᧌��/Tz�kPa�oy���I?W�/����Z���;�R;M�^D��0�|sz�0!��˨Vw�F��~t��Ge�>/�1��~����/��~��M�|Vy���.�3_� ���J��4|��p_���0�����Ye�߅��C��'-�8���iE��,��]��ܓR�XTi*AC��ܠ#^���:�&4�.�WC�<&e>]��7��x{�*���o�4^�%j#�H�����8=�(d�條�M6�\E�"~�EE�����!��� ����[OwɌ��o;T��w��$
�:�&cT������A{��'��3	�K^�'pj9z$N�ė툺��1�Y��ˋ(��/�?o���ߴ�����5������Q�gG�7 @�>���y�p?<��}�;A�q��5�Nks��[�{wGH����BYG��v�Y.��h�@C�޶=x�#Xe����t���N�R�pI�g�#�9X��b`�cB���J.
����j����Μ���9>>�f1�n�G9��2�5l�K$7�q�0 �C1���;{�ر۳�N�^��^hG�3&T��d�2/�	C`q���5p�!�5:nc��Ņ�N�"K��
�����1��#���
c��9��4Fn�."�.�9e^1����C�ɍ�N�m�]Kw䎟����FQe,�����D1���E����H�0;,��.�A�;u޵FC�Xkk�r��F���h\i e��D�JC�{����53����C�];VF���J�p�K��:���64��0��;7Gv�cSv4 ���Ю�i���h�u;g@��z�t�NH�Q�W��uƔ�$�����9��s}�$F��y1,Wo�i��}iy}]�YP]�puH\ �j+�q~&=�2������kY<d{�@�������a}�j�Gƞ7��I���,I�:�ŗo$����f�Q�m�^�� ��z+�M`�ĝ�ͭ��o���mm춹�嶾fo��R|�����6��,$o�%��:v�ֺ�r�?k[;�B�������q���b��.RL!��@�Rϟ���Ռ���!�
���"�I 8���s}Ux{��G�t�¯ �`�0��1����������Y(�M�ll���`����#O��&�,R �@�)�����z|Jݝ��#��:*���6N�N���v��c}������8��h�U;��6���Ãd�X��^�|�e��H�>,*���F����i�&0�hZ"L��Is�����)�|�A�6����4���z|��L̶ቹ�!��|�n���ێ���P`Y?�κ�9�һP9�Y�SDԏ�
�7-�w��H����k�j��xI���u���ƨ{��K��#����а��<gD��?N�S�]>q^u�xJ]�-NO�HQU��Lm����e�_�s���?9C8;�}�NhH���&S>�U��o]AU���b�=�Nŭ�3q붿�����6��p����:��o�5�O:٘��F�f��V���O�ֆQmn>+�Ҡ_֪	�饀5�-XU�J1�q�Q�ş�sQ����F���UڻnO��F�h��4eCp=�^̠��_$Qs�sϓ;u�]����縲��͞|�{`��iٛm+x�~���:��a�,��?J�����aDs�f(ah'���)^	l��DY�h�*,� �#c����2�9Lv�(Kó�K'���BiQ~ʁ�[[GyIݩ ���F�#`"/ 'w�Խ�j���2�m��)	RF��|�*Ul���t7d�
�g��-s��%e�\ߓ*��N�&*����N�~��miHz��Tz�O*i�D��>�.�;Ҷ7��y���N�x�K���9�'��ԕ0Q7֕pRje�� =�Px݀�j���4�O�]��0�ܜN��ҫ;F���u��pdW>��!��)�=���݁�[��3��f#���%�� �%�I������� ��yg�#��2K�KC+�
�r�"��{�4j�mS��s��N_��4NYa�#�1����n¢⨑���NOVQt���{�޿{���5�[mg��*�G٬�/׼��̷Ut�ed���\����Y�,�.�A�:hQ���,��0��z�Vf&�ܥ{�
BU��F6�)�\�XS9��z�`�'G_,�9T'_�Zm�����X�ּZ��8S%2�:�o�~� m��H�$0LO�Q/�-�`�!���h;:n��0{Gn�^�Nۇͣ���n{�j��|�:�md�a{�r���߶7O�UH�q<F�3�{k;���8i�q��?��˝����ޥ��������~A�GGnr�^��j/^l�7ov1���;j�?�c����m;�\Gmg� �ھ��}ʲ�y�>��m���w�}�ў?}�^>����=����ƅ�,^��ׄ��]{��]{�n�mf:�?�\��쀍�p;En�y7�<�y4G��?:n{��
���Oa�mנ�G�0�=��#ä1���t�f���D�45�]�;;{)���v��B'N,څPh�N0��v\o&��e��^�E��ص���=�����3i�q#苎�-.�a�-�1h��v�|;C��@���K�0d�;��Ɩ�d�,=�nv�sk��}��mo�oe��a֋_d=��8��9����_\��_����o�6!L���+{o%X�!�E=?7��]ܫ��Y���K-��$�f4Y�`Ȩ� �_\6��z{}�}�ɓ����h�|��a䞶�����߷_��ߵ_���������=�������/�|�=�����FA"��H?*��8p�6�����Q�`�}�l�={3A�[�SE�ե�HE�������
P�Q�m?��+�Ў7��A�_���`�{]��=V�<�w6nCE��_Dè3�B���<�w�lxl��ԃ����~��(���tX�A!���g��K�֨����;��x�9J�?³��@��Ɂt�g8��Q*;�,;g|��@�oS�����6e<j3��Z[jw﮷��Y�O��.����[�M�����l�(����>n��b���؋�|��y�j#����b��2��C�i8T2z��0� ��9�v�΅N!�L��.j�n��F�@���.w�=ਜ
2�o��#��h ��uYF �b���F���1"O[ʒ��,��nży��w��34,����%�rſ�ҫ��Ŀ�Sy����+%�YWW�Ћ�=.��&����u7K"���w(
�mwycpd:���b�"���:e���A��~dyEɂ�b� �
��7�m��7y��W�M?��gȚ/��Og#����_�_��l�W�i�^�D�ٯE���5���Ȭ��l}id���ha-�L�w4�]x����]Q�'���W_�E��«�7�xOGXG#^�e�q?r�l���TȈ|�� �Ft��*b�yow/
��a썷<�l萻����FF�T�䓔��:�i]��R�u��b(�|�C�m��9�ho�F���9���rm�0�J�0Jz��H�o�
Wr����ر�(��;��Nie���g�K2��K�iv�v�l�N�N�0�]�F�mw�. `@�*[���7�ŰλƎ|[��t2��"�巌
���:�X	�U��-���+�)_: ȯ����L��.��B_���"��I�w��D��E�9~�9�̙�����+d/�����^��R�v8���q�����4j��g�`o0HN������[#��s�J�80/G(�[�\;�$rOew[��C�5�n�#�1�9Y�̓�6>��;~�������,7���r��W_���?�G���;(����o��˿l�߿O��G>)�J]Q�֣���<��}���IC�կ~��������O����y���D�fy����|;��̹?��(�v�Q�a{��ؙ*���sN�ՖVֳ���[mw��xn"h���Lv�t<O (�R���� 2}H�$���C�Sc�K�t�����4R�ǆ�"��
����l�{o-�fݺ��3�A���kV�����q��3;kЭ��1����H9g�Z���ui���Ñ���FK�#��Ÿ�/�Ƙ�u'�I�=y�Q6!q�BeG�`���n�.��v����D��Yc���z-;�\Fa8�[8�q��1e��1��4��层�2@/���w���K�Ӱx?:���ʳ�Ņ���T�1�?;F,��Ce���0*,�k�R"G:��fYz�S�1F���G�`���`�p�mb�3���Θ�U ��K��	0�n����Z��Y:0��6׎��0���v�P@޸���_\�(Jl:����K8*G�g�j-� ����D��F�to�hY��g�ݵ��ȣn�:� �O������˫��߷���Y{���s�0�X����X:�2i��?9
uF�1��s5��D#K� a�$_��@B�P�sa��b��v��ӏcd�Z_��W�t5��������_����^�(B���?m�}�F��nM�ֵ���C0��c����7F��X������#kb?D�\�Iĥ�BHcg�S&]�0?w}�����+eX�_B�&N�K�
�Gn��:�LR����j���فA��5�m��f�!04��x�='�#��?��p�XWF�bX�PEH
��*h	��N�! ����@J�:��1�@`�u��,{��0��i昛ǠmSc
P��A�=�.r�n-�������\z-�N����}x��}x��mn}�Xޅi�T������''<�x�̷���i�����ًms�p�q��p��4D�.9$<22���1{)��#�LW�m�Q�����2k�;�f�k*�︆h$��Tš�uT�C�^�qod�?f����
��+�A�g��L��"?����F��7$��s���ĺ���>^��u��� ~�f�Jѫ��ywβ�A>��(�<�3I�fldmo����{�;� �e�O����3Jш|�T\�M�8�^x�w�[Ӌ�����t�P���۞ݱ��Ծ����K�+y�)�*�O�~�~��?O��e�{T�4�A\(�E��O�鋡~8Q���r�Uufݡ���ed�+?�x�~�����ec�� �8������_��MyӇ��, ��˝�&'����rU�mhyZ�Fͼ�z��ЃPwww###��H TB8�FGr�]Yb�n�1����g;f�Y���,
����Ju])��l�#�Ux,�����4h���dʵ$���0�-GI���H�o���Ȳ\��g����GKD�O�o�:�'|�_#�
Pi�����'��,�t^�w�D
[x��M��o�U0�6�4}���C�.�P�e �}4�^1^i����Ż��*.��<�C��2�-7� }2ç�� ��w�β&�������p������ﵩA��({��z(�n8�|T��TŉayN;D�*C��e�$��G(����o*TYS�+:|�.~�Y�M9�1V��A���H�p�Đm��Ҍ��b`�È���5;����v�������Y{p�~��)~O�>�9f�	kop�?�S��G������(������S�n/_�M�.��3p�zC��-,#74����6�s�D���4nT���ǉ63�ؖ�o��r;w����-�m���;�u�����Vѝ8�,^;*6偑�cd��h�92o�Jk5�ڒ���0��ڬ�����y��Z[����4M�:�պ���j�ҥ��MYp>+w#�����ͧ�I�5�2]��Zdk7M��[F]�E��` )��7e�F�k��'�5�2�HOZ��G�"Ҝ�d���OBU|Y�a�10)�D�z����=:/�:ER*�)���,����P���2�hcuy90�;�G�X�2��A�ǰҸ�����v�uT�%Y��cB8"�����i�ē�,�ޮ�p��5M;�=�`v��c�v�\���F���S����>��є&��YϹ����B���X���Y�O$|��Ä�w��<��6+2MـSV�D����������j_}����+�G����0﷡����?ad�#�9F�v�=��0�N�1�H�,FA8:v��H�1�<�HB�3�$�!��?�JY6t+���z��<�2V�G��G��tKǇ��gh��տo�2�Yw����|�>��S���ݕ��<B�2�������<�#Y�;���#Yed�v$�$F�=6n�ݏd] kz���r��[g6o��J?�QY%��˻e�@�Oc�_$^� ǨG6\Z�$�*��f�R��7�!dG�0<Ψ@G�N5��:���4�.Ҙ#<�ꍫr*�Z�y�D�)�46�9��^�/u�a1;�&;�PaQ�l����gi���F�̤sS�*��mn��z��W������[�ޭUf�����\}��C_�����>妁4w���P z��~��ԇ1����-u��}�ڃ���P׍�ݦ�T�v#�e4k��*��� O���ž�
�&�5�w/� �w\Q�Զ3N
��c��R쌬(г�et�ϡ�vT��a�{�HO��/i�3�� L^H�x��ݥM��Y~�#Y�����������p�R��F�	����w��,G7�f5�T�54��ף���mon��=���2��Ȃht7�,�+]��+(21�"NU|y�J�. @e���V�A����O����eA�k�<s�/~����?�O������}�1q�ҋ�`)I?�%.#�9���I�I��0���]�C�˺��:�F�����k��<��J�E��q�nQ�֢ xLB/}��}�؀���F}H����Ҫq��]��f!�[od�_�(߼}o�Kc�Y2����W������x�aC�UHJ���;�De�����;w�^��#1��p����4�I��5�r��4i��6�6�S1�Y���IG'��B<��K�r�T�4��׏JON��!M^Ґ���ftF<��ߍ�l�����s4 _��h�#l�M �4m�	�=��*_( �/ͯ���_�ˇ���U'[m�-�+2� �?}�ճE^�A��'FG{�����X�&L*�*�^}Z�oZ��[�Zv�^���q�I�Ê�L��[�sE�ƻ���#ܥX�/��Y�r��Y�P9
>�(tk��_ڗ�~���r]�R�F7+�N��pE�Y�mu�#G�ܺ�Ό��K���jSSc�<���ɱ2��*8�jd��wG��D�=��kdM�..�|�Ѥ�,$��EeN>�9^^�U��$������t9�иc�k�/�h�����]hWB���1ʫʳ|'�1z1���uA{h�i�E�$��n��Ȋ)���n+���2�:+5pP��! *��P�wm����O�bq&e�>H�7�}XI���C�f�Kck�����?���GM����6;?_�F���h������Ӏ�mc�o��ƨ&oq�ugԋ��tX�I��/��2o;��O424����:�Or>�['� ��'=Fz�t����Tyu�2��=V�:�h�G ��K8�آ��p�']�*����\ʓsp%���F|�_�"+Ȳ(g������3����C\e �4M��s��t�(����C&:��m����
G���(p�v�i�n�b����a}�^� ��Z���9��i��C)Z6��U�x��mΩ���W��v4��X��HV�:����H�*;�M�C�g�M;�"�<��].?}����?�I�����ۗ�<hWǛ��n���?����HFJ�F��4�OB�Xy���։�����k$��!���B�PQ*�
�pMo��`]]YðZ�)�k++���J�w��,���u�����.�O�/���5]p�A{�H#��-�;Kmu����Ù���Ȣ� � ���}���0�����,��n��y?]�B#K,�J����p�*b�����-�4�Rl�杴���_�r��8��v><F��V��W͉2��><N5��Ⱥ��v��*Q#����ͅQ�]�	B��)6���B��8�#AI\~/!���gc�8ai�z#W�eB�T������<C�g(�m
�76|B���9F�y��m��K���{���{���[cXY �!k��?�~�^�~��c��:�+�h�G8��@����i�;��՛����71��m��#�Q��ˉ�nz�s�݁�ؑ�a{�\�(Ө(� �PV=e�� ɕQ�����R�J�ideT������4"�Q�af�$.w�I�V�Ɨ���]z�t�?��^t�c=k��0�qM?u�����U�HZy��%߇������+��)�|Iy2�Țls3
��Ȳ���m�m;4�{{�M��Q�R~�ЊqmF�bd����7�$s�i���# T�ʘ=����>����g?k����]����ݛ�W���Y�7ݶ߾E��9�1N�2�+�u�Uh{���-�!��u-ųgOQ��u
�
v��B�N���H@�q'�4RIsa�^��S���O�|;��������W�j����yRm,S�j�-g�PN��=�O<��+�����Zz�̯oLTZ}���̖����(N����?m[��L>�XI���Up�5*#^*;�u�����}���)�p9���.�)Z6����lo�{��kl�C*:ȧ*�2�*��,K��0qp����P��g���h��s�3�E}[+��N����]%Oe��J���hKO:�nM#�2�P ?�c��_����k���rҙ�\D���'�^���v��`��x��������@}x�Iҡ���WST��^YN>u�1{�5��o�mnn�����/?��rc q���K��q3��m�m��%>���x�S3�U�TrTZ5�,�#��=�81��C[�^���h�.��KC�TH��{�6tw;��߼~��K���,�Z������2#�I'kU�qQ��]>���H���.�E'bd�]Zt��3��G����۷o��9�!�j�:9:>
�ϡ;S�{�{#_'�y`��W���o?����L���4�hA�8��ƹ��c�����Q,��S�02(�$�Z87X��Z]����3mkg�mP�Җӷ��%*3��Վ"��1�C*#mH�;r�B�ď���O�͎��i�gG=	��/yR_;;�G��(�n40FQO�ɭ\wv�u�!��(�eqx����?���ҍ<+�젰-�����Վ�^NE/ ��`m�3�[md�K���\��\�[9����9��H�L{֣��7��G5�k�g������<�z�&0I+���%ϙ�q<�W��8�Sk��TZ-^(XI�gyO�vic�(�b9���Q��29*l�c��G��,Ҙ�x:���u�<�\u���3vJ���V�>bg� �F�ĻF�Ɨ�H��uy�&����Ì �������:��N��J�C_Og��?�\�������I���ß���?���9����p�����/j��m'_H� �0>H,*w�Nt�/�i���XSQVxz�B<-uY i`�(-z�R(Dp��g���{wrx��'&��%Ij���m�?:<&�4�q��R▐�z�(6�ƒ�� 8{A�?�1-���L�.��OE_f�#nݎ��40�h�B��%�_�˫�N��_�wUB>�9W���/?���0�p��T0�w6\ρ3�  �#:�;f�)~�Afyd`��0��ޒf��;�7&"�g���T"���nM�) QF0Vj���#i���|�.ңi���W���g�
���1؀ź0�!��g�����
h���Uc�C3up|�l�����s��$�����C��#4���IƳ�0�28�:�]�|e$���w�}U��{����DsрL��;��8�����P(0�����N�_�_�#��a�4-M�L:���U��{�yUZ7?X�*ݤ�[�ܿ��3.~�{}|�.��Q��iD
h{��U�� n�O(�m(�(�8�鵁��W��Yȥ\�H^U���M]ʃ�@��RIX[[o���F;���X)�%�$|G�N�}i���Y.�*�0
/��F��m��O��?)c�����[�zE�獟�
7�W�	����}��g���?�� d��=��h��(O�E�w�t���������(�kQ���<z�͆ٻu���ѩq��T���+�U���Ic�s�Hg�O��l�5:�����I�<Zӂ-��;U��F8����K�n�\q���\Ca��vΪ">�XӉ�L��!Q�.,W^?vE��Z�~�[�F1
'ևr���B%~������}������r��]���$�V)�P�S��J[��yὤ�����>�8똿���/�(�����@++���7RxH�'��Ǐ�Ym�bZ
���g(���w��j�*��~㬕�/���}��'I�5ԟ�q���s���}����l�}�=y���yL�?j���#ܧ�|��E���~�_�f�aL�ɝh����{����4"�|��~f�|D^���p�z��#O�u$�Q
2���Q)ͦ![G�Zj������������.�<ks�����7�\��h�r~�ɵ������r=Ոm��]��ȅ4�s�K����B���"4�r6�Ƈ��'O;j쨭S�\c㈲�k{v�v�}sk3S}w�N@3�U��N;ʻF��]8�Fm{)�d�E.:�����д=�*ol���2$R�VJk�{^=��c¦������4�W�+7R�_e։��6�!��ͳ��?/�j3��zrj��wZ�����s�:Թ�9�,�]N��;¢������Ⲃ,-��c��n��S%ů[�_D�1m�����v�:Z��av����wu�������d��5Z��a���!�F�F�X��e:eJ����/�`�\v4���t`\��>��e��P�-x1|�,ՙ_��uL���R߂C35�$Q�ťv:�Ô2z8����?E�B���'���R^U瑻z>��M~p桬���Ъ�v��	0h@� ���2W�Zz�lև����gj�<gk�����Q|i�x�C�1��-/.���%������_�z���ox�'3�L.�s: ��XȬ�,Z��P�ӛ�E,5�d�<�d���vĉ��J�n��y���9�ݔ�
��]����B���8�&�H�q����5ųV�B�hb�d��kX`�����F�)N#�ww���-�{#�ћ.,����g{~&>���>�7���A�=���8�	���. ��ޙ  l1�����s�&B"[�CL�ՙ~z[|7ip�_�M�*rJOX���Sx^�ĝ��m��O�~S�
c�)�7�2FV�F֥��Ĥ��0{>�n�8s�@�,�T=�Ɯa�se��r��5Q��ջ��1��2JӉ �1` ¹IA�+�g�����X�L��gFmăw�)<�8w��M��/:������������L����5-�/���t�t��w.i�g�7���p	ׇ��]���s�w��C��o��Kᯄ`�
����'S�0<�J7����B\�$J�X?�pRʧX��/��	��J0G�d����ԗ'����� ����(��Q����:���7�����۷��`S~��=k5Z\0�H�SGn�kD|��io�#o1ؔq5W�FGP�����V0-{Msjѝ�wbtx֎���x����A)�&~p���k��{~��}��1(�^wrj���Ý�\�y�w/w����|C���E�c���
�#"*���ũ���<����#đ�>j��TE{��4�#��i�e荗��T��U2L��D���iP�J�oGǇ|W��ϝbV��=/�'/��MŸ��:��v�J�W9g�,��f?��ӯ�4Ck}m�G�۹����J�<��H"�V�Q�>Ao��2���u��?�H��/1��P�ݲ\�07K�bd����x`�'���!r<���8==~;/0��+ʩ���^ه�����j�}�$Ӄwc�yV���~�Ϲm�k�],�ʷ;�^{��]�~��K�����r�����jF?q>&Ku�۷V���_~�	4�qרG;N��mh���e,��)�y�It��R���v7��v��J��۟���v��b��<:����ll!np�U%;dD4!��u"��ÐO���:�ΰ|*�KK��Ҋ|L�S�2�#�v �w�SvH_�a:�����v�{2�w��9:�a ]����=t��0I�v���(u�Z�e����E���N?�	ڴh1���b�ql;���2��f"�C��Wn���{'G�/��8��H_d�b��ɉ0�O����e, N-��Q�tF�O��VX[9l;����y'c���O~��.���t��@������И������3L�1�S��^�Yw}��o�c��·N|����W�����R�C+��i� �4h� $/GZ���w|�]����~�OC&������/��/N	cw�ݲgs5��h8>hXil�ͺ�G�C��y�Xq4T�Oö6�pj����k�F�š�W�b�J1������Zi�I��y���蔖M�p�>��:۳N�zu���N�c�L=�h���I��j���<lG��8���B�A�'���?����/^���Ȃ)�1�Pp{#ˊK:�(A+��k�0�Ȅs]��TXS!�Տd��@��iO�ʈ�V��Ѳ��<)sM�F����PB���tfr����}y�n�c��j�B�C�Yn�yp0��:<q$놑�m�U�E�=��$]���g����Sf�󮇕�ӧ���ߺ0n����7�gRȿu���R����U�0�7�`�P��\� �؈3A�H�إ�����3\`�XK����^g��H$��,8�^Z{���rq���zf5 ���GE����N\|{z��,i�0�(���4�<W���f���<�o��C1�v0�\�{
�hd���v��ĳ���d����Q��5JCC���/�u$R7Ћx�Iv�������_��ͺ\U`.�z/��;H�~�H��ӧק���q�a+^����ş�����=]$��ܺ�?����8�=������Y����SJ�tJS{V�)���4$�$��&����M��>U�(���\��� ��#}#vJ��n������&g�<ko^���N`v8���x�tL�ڼT��b�|�ѣ�r��:����7mssEh/
J複��+�g��3My�z�iN�]�4H����������F���޽�>z��-,w�q��G��}�3a��r��k�5(�U�2��֬?��k��(����#	:�e��p�HVh$x �G����դ+��TA��+N��'�9�ȓ���ࡡ���idy���S��x�`esDT��w6$z�h�g啛<eӦNi˴ 噊"qc�\%2���FΝ;���������0�Pλ��0�fZ�wo2��uX��Kd\����u/YG�_��8��	F���Յ����=���67��Ӎh��Yck��RF'ő�#b��~�W'.x/�ؾ{���}��������O?y��4��,��9�XU�WI�cd���C�G������
�,b���^|���z�9�\��tN�������b���o?���k��G��2�ܾy�ml~h�Ч� ���?���Q�j��R��c\c h��Όc쭵��x�~����p.=�NO��q�����.�Q5j9z��v��=���*�e:�0HgWY^�467��?F�m�0�����9�5�y^XN�k�K��C��Z��K]j�q .���sD�((NK�����{Y��,���ed�X�~ζ�"�6��b��+%Q�Se��Ve\�u�5Sų�W��{��#S�(o��_i ;�o�w�
͍2�n�NG�}���@g��)Y���pyF�N}�rq����2Wu���;�9'\��઻|�����CaDؤ	�.q�+i�4��Y.�:�J#�,�a�<0��H�e`(�����$L:�`�g�|E����b�� ��W�M�j@��ah:��Q|�Rfu�
u��s�뢟eV�Ằ�!P�x��74h��t�������`$�P�	��tFE�{�B��b�aJ��^�ݎ�P�Ƙ�%������9�����;��D�HS7T���*�l��3�9iY�aK_v/#w��Z�[�����:��_��_�y�H�^�Z9���J�� �"I�ѵ����6xQ��X`J�I�U���޸l� �[# d#�N%Ɨ�D���4�C�+2���F�����7���W�Zxۓ�W�I�WGE�ds��"�Y�GG��du�-F��X*�*!�蝤l�D��)'���O�^eӅ}��ׂ�߹W��.�˳�^��O\�H���9�1��8�N/b�Xt������cf���x$bqkY-Z塑U�F1t������.aLp�D��
����Y�
Q�+�)����[s��/�L�,��z�81��Sy�X�@r�ݝc`�Oc<��ge���!}v�Ȓ�(!.�͐/#���~5*�[f�����P�7��c�S/UGQ��E�(q���)��?�	��߿p�c���uN��y�x&b��'��D������iyu�U�¾^����Ž�/i��n�
+��=d��z8�����L��ɑ6�O����T�Y��Hc�F�J$uqg�+9Y/���
���=�t�y�9�uW�q�ȭ[���Q��N|��eF���s�Ɓ�˂��b����&�$?x�=��Q���&��S[(B�V�ƥP*����GZ�˼L;=���R+�*h���C�t�ӆ667����������_|�>�������;w�����7.,�+moofTK��2f�O�[�+�P�0J���ᨁ*�<�+J<w�^��eAq����G��YG�L뜶��K��wtd�t�=h�����PAp#�9}f����7g�${�X$2�DH ��*]եZ�;wfw��]#�_���,iF�"mf��w"��-�K��\��եEj�	-3�<?��Yݷ�,�Gĉ����=$B����w,�d��9��B!?�=�3�$��X��wxX��5���e���3R�/�'�9}�-��ws8�
�
��|F��Ke�Ux����_.lO�
l�:��u������o�������=e�������� �v��8X15=I�P�fm
!}ҕ#(<ԕ�Z*�*X�6�sV�������[���(X�}�)�y��˒ܸ�`B�e��\+ ��3S�H��&�a�אs�KJH9aк>H]� `��̵�����ѣ���ö�b??7�>x������^�=�p���z��*<}�$��m�p�$�D��6�I\��RD'3��.�����.�Gg
=m:u�z��m{�['x���DZ���ߢr!���e,���]�RFс`P�����7�v�L�8����L)����R�U,R��mo��Q��e�Q�Ia��W�}�A����5�Uˮ�P�t����/:t9����!��Pw�H؇��U�K�����\PpdK���]ɣ#���|j6�K�Rq���iͰ4�,�nZޫ�aZ#�ܒ{����L���=�rf�ȃ8�uPJo"'��I;��ŹyJ=�s([�8��w�#^�Y���z��.�W?A)�ޙ��o��<گ��T�w�Yt��V)�����Iʳ�-��̷�̓<VZ�t���^�~���<�K2P���DY6�r��7`��J���s��U��w5��wռ�%�*��d�vyw��囖1� e`�G޳�b��`
�{�)����x�	��8�lW�"K�*�I3f��)��#�Uvp��{jU���/Ϝ>���'�d����������Q��/��d��y��PV�Y��KɂD��(Yh�"�Ġ�f-�*�ȿ� ���t$�v�Ւ�����h���$����J��r�>}q9�3a�����ر92gӄ�aU�d=��R�ʞ�M��&����;�(V�z%��VY31�=��'�nJH�H{x�}����7��Y;�����~t*sx�\
�	�
����jڄ4q![E��F���7�J��g�3�kJqǢ��ϼ�E$d<����A@V��c�=�ۤl��0A���D��8[%˓�r�a�T��6.�v��Z�3���o?�ի\B\3Y�1�s˥�P�s����x���Q���剒e��X�,O2�qc#���?�3�u>Իn��ԇG�o���x��G��vn7|�҇qH����a����T������}������B��G.��Tj�%��R|�/��:b��fMZ�5�f絵я�����dh(�
XKY���G�Gjv��ɎԎ�Jb�FQ���ה'��rG�Ϝ=�._����Y���#�	��}Oz��僎K���H�

H��*,���[�D�q���'���1g�\vCAO�O��S4��Q� �s��<�Dk.KǼ�`�B5o��@�̔��KUl>��s��ۥ����c�"'�"x׆y���j�����t���l'i]�'���w��6��Sk<Q������}��/�?�r8���}��	*�5���˕/��V�y���^���:ra��N�w�N @�{��q��b)�P'҆{S�9�D�(��A��k�9 �q���/�u�_q}�2�������>�l�K�܇�b���|����ݻ��u�-.8h�`H�*;��j
�m�ą3}*9��Y�8�����$�J������d�q?W	/ҳ^��)����q��R��	��Κ�ߺ�v�8��S'���s�Vq���b�x MG���{���N�^�j�#�r9���o���S�Ch�XY^oW�ڮ��C�{�&�b)�n>��}gﴓ'��6މ�Y�U��y{�H�!���g}�h$���: %wvv
�8��}��P��&^�moMD!w�����%S �l!.���LL�U%H'��3�]C�I� ��1-�e��B��d���2s�L���������]Qr��=Y΄>�@��<~�(~�qy���O���؃P�!0$�h�WH�����L����U����u��Й���#*�>�:�픒WK+Uvj)�� ؞l+�l~�Ua��>!n��X� ^��Y,�C؍(t��F���Y)z���<�X���G��J��4r��+��'M��m�i��eo�
���Ǜo�dF�0|������d�V^�*t������LZ��� �1?Ɠ4���
���&o͡�7y+
/���,��/�����9��������N9��@*���<X�釼��<�-g�?��U��S�HGFa������-q(�o8(@����̪���%ܼ�x4(��9Εp␷q�����2;�錗�x��9��sp&��`�DrX�ȸ����¿ռvƥ�ϟΉ�'�ηC㴽}���������'�ړg�ma�Nt�!��'��W�� �h��� 4��H8�K*�'�?�~��6FG��h �&�p�e'��f��`�L��C���ܳ1�@p
a�T;��87?�pP�LA<�I�V����H_��[�Q����`q�-��h�  6Ϻ����t�_����8b��`%ֳ�M���0�_�qIU�K�(��S�*�Xy�#y0���o[=
�ˈ�Ӝ9��{���4�'!$׌NBk.�d�CQN���+B��c�����q��0Tde�,H�)�0�_�)� 1LQ�6�m��M�� ��t4���m{����c�4
�t�:6N9Lcw9�0˷�~�8^�a&/�7ڋE:(L��u78���$Q���0e�Nv
���IzI�|�O��R�AtQ�2�d?�u�P���]��� �)�e3֎@��'��b���{��	�O���V�t��(=> ?��y�4e��痸��t���f�ZT˒)D�'����o٪��G��h$�>%-�;���X��Ў��e����~2^����G����a�O�\X�$�XKt��Z:�WkЇ��%}���Rr�o���ݿ���~�Sv��'��IA�9�Ճ�w���
�]�5B)��Ѧ30f�����P�.]�@|Wڹ���a� #����z[Y|�^>ܖ^>��6 ێ4FG
��r���_�s�u��,ۙ3��� q��I�p;�W��#��'iK�Ϝn�)��G�왳m��:{�B����,.����>j�֖^.��~U�3I��'\���I+=�!8�^�c�3��ϙ��O��Ǐ�(�^���G����y��/��饩u��Km�>��Ν��֭k����������/���s�ަ�t����=vTZ���<�E��%3
L�(4�U�mK+eO��/�wK1�w� #���y�;t� f�`�Qy�0���y�r����J�/r��ѣ��R��U���!y!' ޼y���!X��y��9r�������0��߼�>��;����v�$J(��
�esm��-!��7�ʱ��>V��M��U�`�u/Ħw����65������۱#sm�»�hu	e|�E���M>�����*8�v9V5yt��u��7���I�.�7ͥ��;4�y$�����붲� �2�ۄ<ܬ-�������l_���(Y߶Ǵ���U����/~�q{��K��TX���Q�Vr��˗�P�A/�.�;�/���>_�mg0��QW�~����_��CM�P�u���?��j��e�}�z[A�q��8�es��Bh3�pB�ٔ�H�iG&K���Ѝ����9�0=����ڴC@��|� �P���������gO������B�'�(X(\�'��N�{�ه|�/�ϲ]�q5���rۖ�Ll'N�m'O_hS�G�1'�u�ryI��l P�,ɲ�����l�T��Y�Dр譫��25��nH/G׿Vqݡ���>y��9~);0:;��\�u�@��	��!�}��~�z�Q<����ۆ�l�2��.�"V�=;���)�B^�O�9�d �/*��՞��>y���`���'�Oy�gx���=X�x��?q����R�N��k(�7�H��wRee��>AX�X��\ 8�*�.�/��Ea���UJk�G҂6)�O)F�K�_�ޣ4W8(�DF�"��"7��K7�_M ;@{*3����>Z��e�
��R��(u��CX=�P^�B�N�zY:����j�|x]��-�-x~��]Elb�P�Pn�!*eu �x�5�Oq�̳��
f(@�M�'�i2cƻ}=��6a��a=.�>{�D���L'm�_���6_<z�e�#�!"
���U�����KԚj������%d��4}���O�u"�Y�E��k%��:�u���,u����C3��17����8d�M� =܎�N i[h+�7�w�����,��邮ϔy� (����n��gч��2yHj�S���{|�h�e�?����&���=�~�ɂ��k4�����m�ؠ!	A����p=n�G������w�w��4{6�,�We�~�NC���;�+����{T��w�^(Z�ZdV�t�
�+�T�\�����#
0�m}sEz�-.�`��/.m�r�ut�mO
$,͕�Pφ�Q����I�g�J��8�����k-���=O��閌 �y2�tK��֍I�Q��_�㻮ɤN�+��/q4����˼��ߍ��^�n����V���}�]O?�Wn��-t,���j|�}0]�,�����/gI�������.&�&>mt$
5�������܊�
��(qxs�Q?q�yA�,U�<�u�=�/��.E�-:tG��[k)Bvی�\��s⸇h�ޘ��_��e�AJ���1%�Kb�b�w>��%FG�k�1岿�0s8�u�ٽ�{��$�v���K�'3%�vOYF{��J�#�w���E˷ny,�����zFן<N�ͷ�۶�W��4j� ������%g��0��Τ�\�=Y���m�����D>X�{�N�~�Z���Xv���
�Ϟ�Q����l[�.Gk��w$�^!g[,�K⤃��dc� �v�b�ɣ�G���ts��,�/��\/���e�ҭt��ɃB��۷sw�J�x��{�����H�*�.����E�q��}�UO�\R(�\���S.U���K���2�08Ea�y,�7k<X#�5 @����,��ӧN�+�.e�ީ�����%��@��B^�6��r������l���y�tJs���/ql�.§��_�v�}��ڗ_~Eb��hޡ螰��B����(9��2�*gv�V\��<�~�%@�)��=�KF=�^�ʥ��o��8�|��ܻ�_ͽRɇ���%OO�V�!�fX�śm���+����>����1�N\9Z��D UxW1	�I�^t��%�*�\�l���.�\Z�DA�3:�5�GJ\�1�(���:��Uj�Iaߺ/~�#����a<�O��]Y�Nk���jK��>�Y�8D�l�2�H�,�쀃J��_�+mg�A�*3�����P�����F����N�6�3�/V����@�_~!E���'C']b ��H�<'�k�����ӵ�y���"P�����0��E����͸H����rx8Y�||K�P����]bZ3�������C�J�4f�K�2����Th=�V�
{p���ǟ�@�O�c!6�l�5�6�+g�����Pu��z2>��wە�k��O�x��&Cx�uD|5;Ez���GLF��Y���|ۀo��;�����B~�'�� x�G?֧3o�r� 떾��y����'�+�b�?}���?�綗���?�o��_�{�=|���*Y��tG%+�����E�5%i��Ւ`�a���.Q���%2㑘e۟QX���%st>�����,֑#GӱMN��N��X?��%:L�H?+ي��ڕ�%��������+O!�
rmo=�7�ŉm�y
Vv�H�\��k��M������mh÷01�O�n%Cq夏�g�f�)���k]���� ����pAE�f7���򥱓�������O╏�Ҋ�$�u��[��yu&7�M\�����%~�`�{i�斍�3���[��ci�u��ō,���T��������;@f�p˨�ʖ��.�������;��`��<rϻ��7��Q�����>;���x
cFQ`|�{7^b�f�����I�݇F��-aF.�ĭi}�}�u+��E0d��K�-�J�'��_jd:��
�kk��r����ҍt%�1����Js�n�Wɪ�>��gl�yM~��.<z�Df���Zt9�x�E�*!��'��d��Egۙ�)Ќ�{��̷9����:��Qe2������=xx/K���@:4z�§����� �S��Q�>`^����^{��n������n,J�S�~�lϟ>F����y��D�z�B��RGC{�#�(Zvl9�[�����[6>ӎ<p�����0-� ��O��z����W�lл�l����Ig���W	{��'}��^x�%ɥa�Ϊ!�~�b��[�*�u:��I*4.�[F�o�9�������)��-imM�V����<��u���.���ӏ����#�
<K�V�#�D���딋2�d�H{�\N�v���NM氌�?������9!p~�EtQ��}М{�\6�*�=h�C��e��=V�Է�R�5�N{طk4��^!ۛʨ��[�vz���i�P�ϣ@�;{|J�J�v[YZiϞ<�Rt��-������D3��T��O�8q��I�~w)�~o���~��������[�V8������(���Y6��W����@��Q����e���וJ7Yʐ�϶h٬?��y��) OOTH�_,����ݼu�]��S��)4yeM��Z���(Y�
��*�&u�Ll͔ �����^1�e�2�t�����[���~F�%�gC��(�U�)�y��w7ݦ���^{�@��_�@� �{\\��o�&M����8�'=Iq|x��|�i�Sfd%ڡJ�ǲ�~)ۘh�_�/�_�����ހݾ�fT��|�m�U�ӈ�a�B@STп<��2�R(l?�xǯ~��z�~��~�TB�Q�/��'�)�;�=/�R�ec)��P�(�>cJy�g��s��e�4l��̯yx��(��_��S+&T�<yR�Sq7-Ö<�{��Rw�6�Ǵte�;����օ��J��5�B����H>�vO�4y�G�|I�=��).����3Dp�闟}'o.�N�A~ķ9Ȏ���P�(
���f���wZ2��;��ж�!V;�@�}�Ka�'�
 É��m�6,=Gn酫���~d�M.�/O^�]h��[�1*Y�3�ml�cg����_�}�=z��2�%˙��v0���J�Kx`F��L�:�.*���.�%�܈}�)5W78��8{��Y��9Cm䕑x��̴��x�c����L�FD��EshP�Й�U�,��µ�U�<_8ӡ����$���~01_�7|)Kl��k������;q�V��[�[��_�;3Oz�mܘJ����_JU1�Ҽ]��	DB�����W	"���y���a��S5���a��)��<6�AyJ���n��V�Q�r���gy�&v"4h�8k��5�K������ٺ<bA�J@�^曳X[ێ{\��cg����َu��,��p��7<ûN�z�����o���(�DwM?��'��D귻�@\%�|�1��$�I�1�S��L�X����N�4��]���i���g]ů����1����#l����@���5�X%k�}��)����^�2��W�*�5�$�>�î�m=`C��5-���D�QC)PXQPqɂ�h�����¤�)��Q�"W�V��xC���6�ó�(n.u����P�L��G��ܸ�B>(Ax5O��d�~�'�Ӂ'��~,�p�8�
�*9�n_�,��ܹ���/4ޠ��^�u��-��kٓ��у��R�Q�* �޸�������N�=]�F�C����L�oW���Y�.^��.z�����e���Y>U��A���#��@8����~�=�����1��@ݒ�<n8a�CT4T��޹KynG��f��rn�y��@�=�#�h?��2I��~�_|�~���s���S�)
�T�r�ϙ��o���}��W��S���Y��|���CA9��ԉ������do���\<0���͙���ٍk7���۝[w۝�w���(�+�/�Y.���mr���۾$S�z|��w���������\�x|�+�'����OPn�_�������o�j��m����f�SZ����\�� �{�j����Q���c�C�8S�޿֒�����=����Y��y�"x��6V�(�K¹'���*m�
S�W��Q
�)���: ��dMR0���{�6�����tۧJ�3�Q.��?'_"�6��c�4Iٖr�&���A�N���OLσY�����P�O8�;���<���Q�;������{���gO��0��NW�d{��\�|���a8'Q�=����WG"OM������G)�!��`8c&�bûSfqI��	�7.�SIQJh8*��5C: f��]��W���]�)'V�/k�މo4K�i;4^sCȤ�{�n�G�i�)GQ$M�/Ţ~�dz����qu�\2(X��'}B�d1ͫ�ȉC���9�2q߇Y�a�O{�,�E�"�V�.t
e�c��7�!�3����R���(�nS����P�S��-}K�o���x���!|,d ��4�.������?�捴��Q���^2�dA=��	�;p�A?t���>N�=�U��2��|D�u ��;ʻ�:WwxM�+��8XDZ5`��_�%���
�Ű��PUvq	X���O*z�*�rx��3Y��O�'�dec�������������4�E�dQa�}�7An�J�Q(��E�� 4�VbEP���e�!��Qr����(px����
�����G|&䲋�O&��b>r�3l���0��m��u�@�3[A��d��{��>�-`���J�:HV�u��pZ
@����(�At���9o���{}ޭ�"�d6��p	;Tj^}ׂ7s7PR�+���Q���%���������؋ibIX<c�qK̕~܆���t*o��q�Q����o2X����W~�/��8�@���<3XcmcyE%�N�\�\\t	h)YKK*]ֵoݫ`с�`9���ڇ��Y.�R�Q�{���>)���^^��<�黼�����MRr��"g�>�ݟ�̲���x�_f�����z��L��{�Ȑ����+��Vn���K�������=a|�!xn��	@���,��R�e���#�
?��Zv��|,�K!�,��qɌ'Oը����V������6n��T�:<�	��~$�̎���D�hpep�7#�H�Q,���xp���8>��5������
;*(�~T��!�M�>�n;��H�$�&����d��w���@<{x�MM�;Y^w�ް��Z��,��#|�3�`r��مkWD��ʣ��
b)~��aW sمxS)P��]�d��=/AU��zեW(k4H��^	����gf&��D��Voݾ�Y�����d?	?˭PP��٤���,M��
7�Б�0���~�)B�K�2�M�5�  ��TZ-�qaqi�^�x��j��Q���~��l���g���٥J���")��/����������^1,�"n�IǄ�:�?�0=3��8y�:u������!��ɧ��d����}�M%�.
V=��S�v>o/<��)�^�`��#�g���Y�.�}UQSV��,�mo�lgP�U$=��%��Ab�{(�?|�e�]���o�<y
�ʣ�R�}	CylS�K��}�V�7�(uQ���m��#��PXϝ?��Eɘ�2��.�ٞ������������p�B�E]�*��#N�]�9";��S�QR:{�8�vdNe�)�����z���e�u��$9�L��{C�==ҏ4∼��P���,3i��~���5��Ǐ�˴�w�}����{ЏG�_�*����FxHN�/]l��x���	��;�f�~�~�p�8� /8�p�7�{8Μ�Jj��3�Wޭ6��l���K(X�s� �%����! |]e+���^�=ئ�}�`�ԥg��n㰁a�ْ.��3�-�K-���(�v�$�YK~�c~H��'9�C�6�Y�P^���K�0��X�;�RI*�e�3��Q�I��̣De|��]��+�����H�Z}�~��V&d:|�RͮR%͹�?iG�6>�{����\)�%�x�O����/uvK�U�Q���Gf��c�����i�3확þ�����j�N�w�r���D>É�,�Y,Kg!l�*>Q���cZrdF}A���L�-3���.gmU�,�H�B���k�����4�L�X�7q1�'v�`��[��;(�L���G���'�Yy7}���t�
%������=z�(����q��;d�V��tTW��,7�)=#q&z2Xy
��z���,+��Q<�
�V���>�� �+���2�u�͌� �5�x����T���F$Wg+�.]VVJ��Z�J������p<��F����>!m1�
X˃��>�I���?���UY	{5�J���/��(����я�&�_K�����!4�gzy�	E:�h
XAf���_K���`7����K�]��P�%���n�����x\��,V�������ke��z��:\v�g�"X�Ձ(Vk�+~�Q�<�+
Vf��~��R�͋��y��#ʄz{�ɇ]xEW�z�?w�պ�}�$`,�)8��v����Ć)��vic�7�F΋��oeK섉b/EC�Ƀr�u��z�;�U�����[��w��o��w��Q�v~!_���>{���E�����̅(��G�`t���
�L���v:ָ݆L�x�x�A�*;��aU!�R[g���d��63=�Ia��}9���3��{�d֖�x�k���7��{{��	g/>~�xf���W�x��af��=�ig4�va��z�㌀h�Qy��&+��
��*ϟ?A��Ѯ�4=�8
�#ޞ|w���ٺ�J�k�|��O����U��;�&n���$�~�`�.sfE�L��捛Y:v���v�ǥ?��w��wG���dN�������[7nD)���������a��S?v���9!V�S�vV�q���̊3b���"ߤq�  >š����:���=@OX����_���"(����׿�e���O��o_A���	-n��{w������w(X?�ݿ���zX��۩� bb���/:��������.�{�l!8v���5���D�~������{!�:�X��}Z�Q��={�|ml��ό�?}\Xd�8��=DA��oQ�o�'o���y���ʕK�B58�bF%D�׏UW��ɿ��[�W���}���9�������ܷ������9��̚��g?�m�r[~i���r�d����(�Ҋ{#��/�/�w��G�v	�*�@� ����Y�B�p�r��޽�>� E�W)�!#�+�lw���೜h�9����.�i?�&����wX�:|�f�]�IQ_��f�����c�����8J�����J�E/wF�:s�l�ʈYp�i��ۦ�]�%ʙ��^}�����~N�:�ȝ�rf�Y+�#.�q�E��9�p*<��?�P�����K�a� _m�\A���:�M�\YU"��fl��,,�K+���3\�+ዦ�[���M��P�-i�������$��}�U)k�+���Ѝv3�(͕�>�_�B�fC,�e���j,���Yb�	��MzCyRꉟ�-{����P{���6�>�S]��ݞ��K�	�r+>��V��Yz����8�(]>�1���A�Rڌ�|%^�r�ʮ������!���O��R�6�<
(m���F�˾���t�hm%I�5m��2]��Ym�I"�r[�QfEN�͞^.Ͼ�t���KLk��qeN��L(o�NyŃ�G�4t3��7�d�⠄���s�3��Ç��A�������Jփ�(Y98�=/f�վ�\�
��N�-+hP��q#!��s4f�,�?�x�
֡��`�od�7��:�	s#MOV�;���a�n��:���m���J�G3Y Ĭخl]C�Z^ߗ�:�
��.;�B� >|��d:8�,������C[�O\�T�aԻ�O��=a|5�X�)N{n��f�%�{�n��1�N��J�kL!�]d�0u�?�le��:������E1a��,�w��i���@� ������R�BԒE���ۤC�[��h�<��j��rF�%���Tmnz�a8j�`�!�)���/���M�Y����v{l�h�ZvaB�����wQ�zL��������phC�W�)f�71��<���_"�Sԕ˶�i��[���e�ko�ʣ�
7��x!�aث�/�?n����Q�����%���[V��#�2��𢌜^��t�mҳ3� >� �����C�n���*8�ɛ�P�N�:�N�<� t�yw��:ꮰ����R�VW��;��J�S6�G^]����~q���ctTb�������k9$�����x%��Sa�?r,ˇ."|�=w��Iמoe����\��Q�*9.3z���(���%k��Ir�K�\�5,稽O
<.�B��b=�O�}\�_DpFN�������\�� j�]"�%�}�����ٕ:�ɋzK)�q�y$#�����oJN>��s�Q���`��w�ܷ��A	xˑ�ڠ,��V�,2t�p�JH�a�E���$��6B��~]ʄ
��cs�k��'�QX���������7훯�'�Q�k�����Wx�o:k[�N�;K?�����K��{(�����Qfo%ޚ	� *< .M�`.-��g��l����)|ۙ�����y�v�F�����km�G��}f�ߺ%I��k�͓ˎ�Cqy���o~���_�3��I.gVU��"�O�x�k	��Π:�#��/���%�΂�@H��cIyE�D�^r��
�k(��'(YK�*4������و�2hq�'B=2���N��ﵷߺ؎�M�i��竡�����/�c�Bp�/J}��˸�Qg�]~�/�F��A��m�*eE��ˡO�8�٬#�#�=?q2�.GQ��K�Mۉ�{H\&����?g���<�3���~��:��9ܼ7�po�U��{S�_���L�����G�ס�,)Y��\j��;��$�� �= _�vmG��G�K�<6��ãz�I[y��Ct��2\!�U��<"ڸ �2ͤ��Q�ʿ2�p��p�!���>҄$7�Siv6M�~�N�{嶒Y��q%݄3o
��8�_�'xĭR�p�7�U��#�Gb nx���f�~�iZL�o���SN��/~�����8}*���d��?��)����C��z�~�����J�h�3�$�et鶇��������	į��[d^����>�'-�`VyVZW����xp��\�P���*��y��ɤ�q$ʐ���|���4���,�`;ql>3��d��i�S�L^maam#ę�����s��$ <C�*ҝzT����T#�^��~3�w:ܾs�}����w�������}����tXW �L�J��>��!�Ϟ?��z̝Y�:��Ϟ�]��5|�I��Ǳ�F�=�6D�+%�B���0��r��E}�;|F����=M���$2:�1�%�v�f ���K�g���|��!�̶���m��y�9��Y��� q�� �z����$�
�:�v@���7�4����"_����Fk/�����v{��ݞ-l��/���AI�i��j�x�C��������	��v�-��2�0P�^إ�P0�م�w=��ݟ�'u��������Lǎ��V�F�Mod'_����s1������,��7ؓ~b�� !��W�O�>����3�{�ѡ�arCǗR���ϱ$_e��	�W&��
�n��iZV��Z%,��#�Jk�n�/��F+}�Rk��2��_�؁�l������)�}�O�=��f��Ēokxd�	a�D���G�ʌ`<�V�̻�f���3�,��X$&��4d���g�]�7��(�)pyהy-a�N���X��2�q087��~��ʯ�����y��(�U\��`�j��p��L,�l�L��l�vg�Y'�=EGw�2�8��{���=Q��SaOٳ�v҆5m��YЏ����ˆ���w7o���P�)�
��E��b��v�hS<�@�u��$C�߼�E�to��˗��k��\D���l���3�ŗ��������kWo��G	��]H�7:sO�s�C�Tl��zѾ������;���o���m_|�u���P���hx���IK'����(���#�7v������tig��ff�0<�[����"� Qʈ�c�8�N�F�m���1���J��������_������Kh�r�Yգ�ԩ#�ĉ#��E�:��}������_�����+�/~�v��9�	�@�*ڼu.-�\��s* �sH�|@w/��'ϟ�'/��EO.�������d�[ɡ�Z����@z9&Z�ᙩvR��g�ċ�=}Й�&�h�ꬺ��6��)�:�mrΆg�&q��sx�0��x;v�M�sawT�z��2�H;wt� a���i����U=�f�0����i� ����.*��d��G�W�V9s��3��sG����;��>:yF�t�O��R6�N�`�?�����˽�v�=��e�,җ9�E�hH���]���|p�
C���Sʖ�j������~
$gÔA�+����Q=Y��#+Y�Ȩ(�?<ǆ�F_%O�<P>(h'^�Z��L<�Ŏ�w��e�ivU�ꔁx���|Ԍa�����#�i���-���m��Ϟz��f���>�a�j~_�>����(��-?��?�B��T�������>-�uJ�!+�t"�������Ly�n�Ï��uO��O
τ�_��d���ψp��|��� �:~5-Od�4_)W��'}�}r��xi��#O������I, �Md@v�3O8�6��0��2���Qȯ����=
�ߡh}��W�;F<�Ƚ)�q�2X���^' ��
�+`����W��a��N�QH�[w�=��[���V&����N�Â�#?=�|�'i�Ê��O��`���H�� �Hf�T����Ql�P���(��0M<�V���]�B��:�	�l��|��p��l�D	#L��S�0�I;�0wa|r*�1s˾~U�\8NP�^�;�Ƀ-�Wk�jiy�-��n�u[�����m�\��լ��l��)D�Ș����������g(AI�s���ۊ�ۺ���k ���t�O-�'a��k��F�<F։@chԁД3���<��覔��*z�[��$�{�z�h�<|��9�������V��khg<E��,������b�Uv�G�]��r������%B�e/ތ�P: ��$O��̼V�����K{T�5v�D��w�o���J���2]�H�H���Y�Y�6G�MCԚ~�l��_1�q��)+�=w�e������L�p��K��=i�Y���<���\����t��{�ϙ�\Ψ2 ��6
�8S'X�ި�T�&޽�p�w��"�QN��9�%
�u��]7�Q��z,~W�:���'���1����G�7�6Q0pKQ�{�����a�U���.xdv��8�R�s?�BY�W�]>4g�=@��W'Nk3�ĉ�N�O--G���ru������p��M�G�����]9��8�R��_;c/c��}ii�������������}�ۏ�{(ɽ���ټ���B�~�v�l�����)����ę��̅�(<�b�<�#6E�[[����y��x�H����r����ז8��=����3�O?����a�t�<4L_!�A�r۠H�'��9�h���/����7������蟷��{����f���{}�S���s�\w&m-���z^^]n�P�Q�W�ۆ�74��%4���]���{כ��!����h�PzI��c'�W�Ee��Df������@,۔#���/����Uh�7G�W"�O8��5'��DљOې?�A2^� ���ܘ���5����ݎ��t�#w��LA��?��.��*/���#T�\2,�Uhm��p��Ye�TFAYJ�A#*�ڊm��7�����������?�̲?�\�X�JE>�2�ϙN�E�͖����<��{J1���$A��'�/:�#�\֙�g�@�����'�(;N���Tکx�y��Rg��_{�IG?�ҏ
X�����2�+�1��-�����7�!�4���'��qi�m S���,��.r�ni3q#O�5�t�=�*����F��})�T�d�K7ІA%<iW6�>�J��K@�՞&`wTru���Ĕ��O��B��,��	k$�	(��_�U��~ހݴ��Ζ��{��y��N,�m���d-h;QZ�Ql{�J�?�e�f�)B���� P�鬬D3h(�2�v���֟�?vf�Fu���,]p]�M�I?{FlA�;�yN����N~O���`�[�B��Vnه
߭����O�Խ�����SX��`a�M�0�h��#n0�ė|`v�b��7!`!{�ͯq� %<;i��U�@FF��h�Dpf��8y��J�M���3[��b5�Y �>�_`��m ?�~SY����cz���Y�~�d��on!!m��o��������9v�J��B��=`����SJUWnp�n��zz�`���D�h���~v��;�Ô9�W�)ŧ3��n=���_�K�n���
z|=��~J����ӊR*����|��L{����fP�e��$�B��ҶtY�3o�!�/�v�B��2a�M;l��s���(��B�f���[P��b���}PԆ��t�f-7�H^��)t�\�P�Z�� �JyOGa�
���2���'�)���(;���ȋB��9zm��P�h�'��j��j�o
>�����⡢ �U��e
�}�k7us��S�^.�̱�����'�μ8���o��w)��u�C(V�4���`P���̷E�z,�S�g}s�y��K���WU�~�-@Z
L�O�B�v���͏Jd\�UH໠��L��4��W	`uxG?�-��8rT/²}�3�.�R�&�f�שX.���ǟ�����nݺC�V���|pzf.��*Q�&�j�|S�q���Ż�<=}��ݹs�ݼu7��?���&�~�|�Di��e2#�<��ޝ!={�l{����{~�N�9�#�-�t$���:�:���Y��Ne���Z�-��&������Q�����ӧO���ٔD!F�t�h'zﴜCas���'�G]�Ɍ.5��B�{U�\�;d|ԠC�p��F�b	�]D�ZE�P`����t�z�F�I�Jh0"�ù�T$��َ��"�Qz8��s9+��Ӝ����8�Ʉ nے���਄Ey�|���H��0���IO�N���I[�ʥGW��uګ<��b^.�L����Zʌ�˗�����u�W,P�S,{�~��B?�U�T��g���I8P������.{x�m�S@��=rOx�m��fJ�	���屠\�j�I���)_�G��<bۺs��=��(%��-�]�5>�����m�'�1@{�-C��lf@��䕖� @⿸S_�!��dWS:0��6&؆G OJZ~w�q��G3��R`d7΢�!�(tЯq�]7�˻��'��C �?�1���9���R�}/~j�U�O�R?�=����TX�m�w�0q�M~/�WځK���F��/�U�-�	�$O#:ѯ2���Y�(����?̞7͡�M��!��5���F���Rkd�la�� �OYT�\��D�h�v�M �*���������>kO��8W6ڪZ&D����3yp4�!���x�v��rDKRٗ� �ps�B�*�䈮��T��8��ĸB78�r,%�����:�>~�kj�MOxZ	��tPP�.���X��ޝ��W0���ve����Z��^�G�S�݇ !�c�3�f�ʾ�&�� !��(��"F3"6�j�0�u�=S��턷	�mԙ�g�Q�0z*�h��W�u���ӱ4��R�/�q����|�f�,1�/qmc2�����1�����0Z:�A0��7;�(F�K�bό�v��?�{ �R�����6���,Yt4x��ڋe܎'�RN�����.��=W��:pd+ߠY�uG6]R�咄?5�%SCC%��CS�3�I�E���ţ��!��J�a����n�9~^���Έ;���O������e 5�W��(<�k��H	���s�ʬ[��߉[�W�4�op�v��e~��W`���mx�6��	�W�mL�[c��PM#�:�#q�[ #��pE{�OP��n���j
�+���
|�
aoFd��)�a=���+�������f�w[!�4����7�,��L�I=�	M�Az���y�.G��E���G����ۃ���e�GG��s)*��;A�v��v��Y�cIC!�G=���ֽ�ʑkis��v����2oˡ0䬕��s��h묊{�܏3N�qO���<��Ν�m�����.\n��]@��O�l�m׮_�)xf)�����"|ɋ�W���x����4Hk����>BE����y��M ,%�'��'����O{~՞<Yh?�t��b�@ۅ#O�7P�"��]� �#h'�5��u�q͞�K"��|���F
�Y�	�@X�N��\f�c�(So�P�2�w�����"i�ʉ�gϜG��Ц�ͧ��]{�=������u��/�����_�w</˦��}���J�8QȲ�E��B��D\f���(���
�}"B?�ʛJY�R�=���m�y����[�_�տh}�q�	�!�,��	/}��~�������������w�������:9��V���,�q�����-�����u���4�q7N�T��`�yj���V[Z�]�6�')�J���D;v�p���Y�Z%�[А�leu�]��?hO/�7�l]Ӟ
`�O���#h�6x�ĩv��=O�h�N�lG�GgP��)K���ŵv���v��#����j�RQ�ڗ�-�K���m�]l'��}� ��e�?.W?�"���ﷷ/]i�N����о<�l�}n�T9���<���i�ʸ�T����躵"�QLR�󊃍ug��)B�3�t���򑧸BOS�|S>�~�U/=���.��N��۝�x��q��kdy��K�3Ét
���O�j��#�bc�j�����/���� �ρ�Aچw���b�&1� �pWA<D��K�����5m�����A[L�.x��nQ>��x Q���y�ȓ�<��z	-A��`�]9��{�Y����3�~�+������үf��rTx�m�0�>�Ez-%�x�hF���'yX�ˌ�򡛼D%0�f��I?���y �ˁ���w��g�(9��0ʋt>ԋ�(�
�����v��Op&c�=��k���W;n���z:*p���vh���(y�q���k. �U���3������E���ɸv��kշXF�I�8�Y��nw���d$�x���d;���G���3�~���L��)p	��S"#��K�F��h��Z���װA����a�����A�[�o.w����c'	@A�w�r*�Q'���(�$y��/*�J�
�l����d	�v,��&�+H[�+��C���w���;/y/�E���w������ppמr7@^�����������[�V܌ ���#(J�6Z��Q�װǪ��)0)LL8��v��>|��Ax�e��������\�r���^�Wl�C{�E�"��LW^#"�5UJ��|C1�h,x�P
�Px*�D��i��
��˯׿&u�����,�t ��0���PgמǴ��;|3�n\IOz0͑]���(?��c�#P�Ը��?���I�1Ņ��6�q"���=�Π Nf��Dᚤ�c�R:�+|H��Y��#>��V���lٰ�!���#����93����D/r���zr�}Sy���#��pɗ�1\~�Ye/^�����Q�ZE�qt�x���t$z~�fyȏ�xjp��u@���v���M�4��q
=���a��"����G��?~��=����lZ
Y22�'� W��~�e��s���JޝEqt|4�E���J>=�{1b�|Ѯ�jt~uu��,5�嬺uT��V�U���B�:P���m
Q����4`��M�S�*��ԭK�$�w`(�n�C����
�9�^g���kye������v���v���v��m��g�vr����HţN"���)O�o�J�Uiw�3�(Z��}A
B�Cƥ�`yr�>t�
��O�P\��V�r��v�����F )�ŅU�����A1�����s�i�l ��"�%>"��2�!B�X_՞>_i��h7n?n�o��wQ���~��n�}�2m��I����������/�>����a�S.x���g�s�Ҙ�,��Ki?
5�H�u�^z;��@G�^�Wo҇��ϟ�l�z2������ΐ����5�Ryw�����%�.iA�?(��h�(~��M��xf]"h�9��!%�<x�=x��v�(���cr�wϑ�j��0�W�%헶⬔�Ҷi���Y��xy���Q~�)s��̠�j6ݣ�;� �Ɲ<q������ӏ?n~�Q�t�r�qF+˪�g�m%�%ګY`��n�G���Cg7��ĺ�q��ݨ[�<�g�\J�	�lR�I^��п2���3��>A�Z8@�,�[f��,���9(PGok~7ny�x�,ɘ@�q�{ ���k�7�$ ��_�!��t���!^�|�N^F�LQԺB6ę�
��: O�y7�2�q�K�e�r�ڻ?�^�I�' ��0� ��?�$���O�f�eHs�����	����,r��)�_��M�ػ�?*���{Cx��I;���]ARiu�(L9��*�o�_�ѿ��{�e�} ���HE)z�YQt��ϐ������X�ȷ2{�0!����B�3��+7��R�
�(;l;��hO^{��������` В�I��@��2����T�a��Nk)��U�\��&�I�Fn�+��=|�∛��{��p���n�˾j�CYb&�J�{�c}@蘊^��՛�@�Iz�hǑ�{�f�����|�48B�����>�f92ٚ':�Q�be���AGRs�ǰ��}XƔW�,:_b���[w���{�>��{�ud� ��L����c�ײ���`��0	1
��^ ��_e'�ʡ� �n��?�O�a�nq��!�b�0�|� ���Fi5.Î:蘎CE+e౎��I6B��[���m����*�=�����"<���x�'vh��N��A�.�y��q�q�F��;w� �,��%d
X�)K�i�C��^!Yw�m�@`��֧p�<~���	t�X�NA�)�4���4��]�2O*h�KƽU��o���^T��]N�0�S����dh
^@�R*�Z<��i�IDW��{�\��x*���D�i�r�hgN��ۼFɢܹ�Ve�<������T�S0�X3K����F`^�+�a�5ʋx#���N#�`�'~���^��P��:4pTXe��(��,oe����(X����D��t$�t��#g6�����VVi�t}W �rM�c緎8+�+Ļ�����%KY	)�-��!�S'P�.�`��N?�0;��:�i�<m_~�m�w����o��v�֭����ﾂ>���ӈ��I��w�O��k��E���������l�_��������E����۽���
J�ֲ�'��w�m���/�'����:s2u�������Xr��|-,.���%?�WuE�����.�Yφ��Wxo�{z�A�g�⋞/���-��[iK�(��ߤ3�A���%3��Lу%�w�0�d���)z�|�������?��C����׏9._��6�Ld
���H�ҭ{��Cp`CE�m�k�}̏�3�3Q9�=�?�J�Aq����/rł<��S'O�\]�E��?t�|8Qڼy
����?A\^�x�;�8�X��ON�'T���OB��v���ȿ�]F�<QN0��١��u�R��<���_d���ٞ��euP�a���b��R���?u�Aؽ�=�.������L5Ph����w��4�4|mdH?��ۏ�B�ڿ'oo�0hs'nev;���Vi�P`���5�x����L����3ēv	�|wߒ���0�t��wM�o��qv��`��n?g~ę��ք��@�Z��f�Z�7��3ƥܖ�5{�Y��粛��e��cP
F�=v#��q�x|�]#�EPe�
�~����d����<�j#_�V��2f�Lc����ŏ��Y:K�R�iՓ"�J05Z�����*�R�,��0�(^�u�G'AI�"�hZ���^�F��=ӭ̡�J��������;�������[�FaH�4{L�?t�v YR�R%Jծ)�.;�F�����|�C�_����C�i',P
��r^�\���[Ձ�hm�(���@������A'6`�ey�U�E��*)	���� �؍��7���u7��P���!�G�PzͿ7>ŵ�'��8��Щ���.0�}׭�+��$�4����I�\v�3.�ف���S�U��&�-��T���)i�K¨��0kR����F�*�:��{ap�c�s�eF�IG�*a�_�Q��3���3���+�4;O��ʔ�IaW>g$*�5#挄B�T�AX��!�<}�,�֪le���y�"UJV��:4�À�����0�e�%�Ǵ�Oe��B��WC,��6$��C�P'>�bx� �v-'a ��G�;��X�.��+��ʞG�����$nq-.	��3O*�|J�}�������xQæ %J�U�@2�`��ŃiU8���wM��e��͵�YO�<��<�י���z9��vE����/��O�?�S;��,����� ��^ޢq�.� ]��� �g#�zX��Q������Ց�����Ï>h~�A��z:�xY_{��ӥv�Σ��?�?|�u���P��oV0�kk��f�KX��[~���W(k(+/����kw�W_��r�U������������}����j_|�m�v�&4�l�3F5`�L��8�������ˉ���L�d=y�e �j�%q��q  �9��4M��rZi�IW�C�Z���+$WE����F��(n�*OĹ�Ay^��������ʊXXE#*y�[� �qɮ3��J�Ҕʏ�����ޢ��moOP�T��G����ﳤ���[��Z@����8���=�ovV��0�9?��?�ƫ��U��9�r?Ҏ��Tlq8<@��N<0cyi9
�;�w/�~��1��xށ���I�@L|0˯,'v,eJ%��4����0��܇w���v���F9=�J�2�v�����K�k?�$i(gȻ��ʅ������
�}DܪI��!� �H3�	�����s؄H��������|�xh���G�k��q'�������w�i����k����	���F��e�>BY�d�:0z'��)�ߊ7%l��nk��пʇ��7ݩ��Mt+��������4z��}\��@�f�<�����Ǵ�~�!�/�K�@H��\�o�r�#Q�$n��tބ!�x�Y�K�U�R�}���2w#I���M�������DZip�A�*(ƨ+ê)m���N�oN�~�J�!S�d��h�k�m_&k:�({�	��U���Ά�N�Hh�vf�����Pn)s�x;vͲ�.�H�w��y�0OQ�b����L����O�)��=e���q�/��*:m@�H�����U�]o["K�4�b��G�Q��0��=���f���(UQ�T�����DL��n>��r�����:�:��w���v~�z��-���F�qo�r����~걮m��y4{�i��/�n~����������i���������x~��`��C���=� ��t�' ��}��T�2�I���M|�[�o��3�]�_-g(F����]���M���_l��=��4J��Ie��n(�/�/�/��e<v��_x|-���J�3��Z�5�N?�N�<�S�.d�.�q_��I9���C
�<X�@+7߼�mXB4l0������L���D�:
�J��F� �V]֢��C+`H��*�>��� � ����U�_Pv\�g�*zK�����&�����C����(VF9�ҡC��<�f�IS���kQ ��aF[(2*Q�p��쥥��gI �J̢��=8�/�3D������v4s�J�ѣ'$ϵ'O5Ot�n����P��ً�P* �$����b�U���Ż�\�P�f�����i�L#e��*���6�c�8�&��D���c����i�����տ�g��N�:E=O��x��f{�d��>i7�ߋ���b���B���e_��� ]�Q�|ãݟ���"��C��k��/�o_}�C������ͷװc~}�}���R�k�����u���(2O�t��\�|�p;u�T;r�hh`�����Kj]���n����fa��e{��T읝]�ֱ�R�N� ?����>>�@��R�l�ݻ��r=h/^�b']Y7��'}�7����(0.���۱m\<Ef	�Ԍ����ǧ��ݻws���;�Q�d���p���"�P�#NBc���J���c��v��:}��<q*'!;����;u��?w�]8!w���R���p��RT.�ޤ�_�h=m�<l�ߏ�u��m�w�=|p��x�����?p�\Ar�Ţ�9-����(X�h����%�^�|%k�|8�
m��Jz��:D���2*v�4�-�tTr�L&�G�ь�6Fl	�/G��!���7 n��Z��>�WΡ��^��Ⱦ�wd�����y1΂�CS��΁ �0 2����q+;a���O���@�Ye�{/s#���w�)4=�?c�����R��{������	��8�ݟ�](�$��|���Ώv�A����)?�aZY��#yM��?�L>�/����?=������=�Tږ��,�T<�0����������`��>ՙ	�B�@F�3Ed�8%�������t�%���e�$#=a�O�'H6t���YYH���A/� qO�> ���y�+l:m�{\�H���בM<��� i�Vq��Fe��	Ĕ9r�{����>���l=ͤ!�"S��HF��eʗ���증w�DJXd��{�sxO]nԩ�rx�h���_���q�w��g�T�2��t���*�*~�c���x,���������� �L���;���(#�m<��RPv�S�H��Bs���vR��p1��×�N���4m����c�8�Ƙ#�] @@Z�,4�N1��Y "����3H��Ҋ�Q�$�k`���Ifg�`�Ly���G0�S&(���.�,1�7�O"N�J��yh��'�����=!����.�QQ�.�*O���u����TB&�(B�K��1㲬���;�s^$:�K��o�#e�#GֽJ�0Z �Rˮ?�C*
z�%s	M�S�h
W�w�JEL�J�Q���$���ómҽ8(�֝m��̪�N���ŎSڭ���4?��M��@���=|�BR�Z���w�es"X%o|L�����z�>
a�W P�TB�'o�i��Xv�#�Q��6}��T��������� ��f{��&���픋�mmAO�ħ��m�Om�G��t��:
�R���ˡ.ԧ'���iğ�����_!�i������3�~&TYo�o��ﲏ��ЖK�>����[���?k��\�����Q�<�����w�������myŻ����(V;���J{���������n_w�}���v���v���v������o��������������?��7�m�~{�ݺ���#�ݻO�-8�b=x����{�~��z��_������Qf���t�ԡ��.!�]Y�.��p���!�Ʀi��g��2s�������Uv���Y�rEt��;��_<�N�=�=S���/Q �Ǐ�6O�T93^���u;�B�����厰O>��]�p>��l��|j/ʃK�ȗ�!��.�V֖�������((*E��=Z��Ss9�F^a��j9�r(xR�a�a�K�K�l�;�2c�~������A��ߌW	�ߌ����!.��^��O�۷oQGwړ'��Ң�l[9��G�*���Bۡ�6�9�ڙ�g��PO���V�wGfH�#��*�.�t=&�<��K�r9g�+���E�(]]�-�t���B2���������Ю*����Z�(���`����80o�	:.ē���K���=0�1�[e��=�q+�����x	�
*�1)� �Ue�/q�R��'R����0�?~;����99�M��a���׀i����z��%����+?� y�N��;��J�~7?��nZ��i�J9*anX�w���/Tp��#��:ؓR��,b<�2Τ���^R�����K��;���n��A-Q�̤���t�6(��;�m�$���L��_�R��&'&k�����:����Ξ::��h��N�@w��3~/s����^{��i%��3(�D�ݸ�7���r��%��?�+�=�n�pV"F����iT'�o�%+?�	=�� �W"��e�{�d�] ����~�5G��m��M����NNa��[k���P�wÔ�x�2 �O�*�ho�+܁��g��'@��0z��)N�/��S��M5D!�]7�u�Z�ȇ�r�u%�!�ݰo@�e�[wH��tw��R�ڥ���O�xP�)�p#�t�4�ЄvpSI���&Nx�2�B}�Sߞz4�ݓ�<1�S�G���-
�B։�yD�, {�_�7О���Z�� ����gaF �w�!��ȓj��=*\%�B����]˃jy�3%
o�e��m��]|gF^��qτK���r� ���͛��2�i�
G*s(~��K��ᢨ�dWu�~+eBA�y0��ʌ��4�b�:���wx;`]`�ʔx� �&�x�/�]�P�P!�d����I��(z�#�
���4���\���r���ʶ}�]��榇)���f7
�7y.I��K���)��RН!/�#�vμ�筶��,l���}����e�(�
�Y��i�_	Uҕ��e�h����S����v��i����ԛ��Ba�6���}fj�ռ�Z�<������;���s��D�"����*J����7߷/��U���۳�D,΢p�C����~�m��'�_~����Ͽo������~�e����w�]m_�d�����e�޼u'qm�8gy��\���6���ŵv�����?|K�ߠ��m�(�VV����b�� �e�%MF�P~!J he*J��aOt�u��ע���Y ���%
�&0~p��ε3�N���q��+g^���k�a[�Ez?��"��������_}�"���/�����ߎB!n@6�v]� ��((�����4m~�y��sgQJN� ��=y��#"�_3��|���{�l��*@���
B/�S5K�rL�;r���l�\y�䧟|�>|���S��}���g����r������#�IB�t�
�����zY���r�G����`u8h�k���u-�מThO(�cАe2��=-;|���k�����N
ec�����#��_H�r�3?z���kbPf����U�v����{�e�1�B\� e��|#��κ�n��9���HF�տ`�?��]�7����7�5����� a��8{C������*��+H<�!T{���m�W2i�,i�L�G���Tڲ�J<��ȵ��,���}˾1��?�zL��� _�O|��h�|������C^��q3\A	gء��x@%�#0R0�3;�괻���oZ�q�h�C���1z|�'�8��R��3 �@#Kȋ���7� ��������w�ۉ����|�A(/V8v��=����w��&���oA�t"ޓF�ͼ�4*Ϩ|��=O0���ü���7��|t��D@7���X��</��OCL�
ON� u�s �C��W�6~:Vb�8b��P�W����p^0�_?�&��^ʩi���}/��I�û�i���[��7�y��3��=&`{)�����7�џ�����_`�^��,CǕv�@N��)���`�{!���aϻ߉?�	]ws��'J���� �"�.�X�L<��(X�Kޣx�7އ�I�ա@/���Xw���#O���붍��=N.��u�]�+yP,�ǐ���d})`G�ϲ0g� �v!���|:�(��S��ŋ���5�	w ����'�3g1����UJ�;��`*h33ӡ���B.$��-e�1N;�����l�w�lY&;$�b��B�qJTp�8UZ���e�H��JeR3�?
���P!RLt���T^�W�?�e�S�)��I*�*�x��%�^'���H�文�tᎢ$έ&f=���8x�}M�Dr�YO֥K7[��Z]BhO0�F�>�ߙ RB	SyT��U�L��{�\h�ڧI�5�D��)���&�/�w�m<o4�;��3�δ+o�UG�c��sh�ayy3Ko޸Ӿ�����ڵk׳l���-x&��M�ء��o~h��������ߵ�����b�?�$}��u����������s�E��+G�]^Y'łSy�������Ki��9Jk�K/۳gR�
�5q/��d9r_�'Ν�����=6y��Q�깴U�+> ΢��ڌ` %k��l��#�(Xp%D�ؖ���Ժ-D��Y�lfv
e�h�|�|{��+���|�]���p*�*�ҧ������-ۤY�.�Q�Tt��u��z;��.]�����e;�t)� �.:�w��Ј�	�&�K�uPm_��Dg=w�3f.5<w�\{�w�g�~�>��3����4��/��y:w0[�C�r�;��;�(�,z��0�9��9�De�.�Ď�['�G�:��/il�I��-�6���^��C���`g�;��{}&z_R�n���y���_�i�)�Q�~�1�w%OSa'�����:�u������=P��է����K���W��7���_2�ɗ0C��'����i�/�*]���x�<��v ��`~�·U��la��V�a "a�;�{����%e4>�|ׯm�x�y.>���Un×���;^#��������@�y��G3��"�g*������@��*����C��,��m2����C�vy�0�h
/*Z

&��r�c9�|e�Ub�u�2աZ��n�;=�{��Ћ����x��N�G�0û�<��;�/��
��������I0o
�2� 2��ih��i�1�
�Ʒ[��CA���p�ﯱ�C���7���+��N��a�o׽~�L�������dt�;j7�Wy����-�f|�L�R֢3�����w7���`��6u����;H~`7h*�rILڻ[�W�63�I�k�u�(���7A��^nD{�Ð�l��y/��Rq'~��Q��?i�oU�o��jJ�r6�N��t���JD�� �0@`�8`+xFu�� jCT����E3
l/�eIxڅKgR6�(�xD���\jfZQ�6�T�8|轟�Qj��5��0�/=G��3��Bˣ�uV���w�ލ��P��LZ�k,��
������yO;Ζ�����0�h�>/Os/�T��A u)�mͲ�T��#!/m�zt�34*xVHǵ<��O���Z*P
�~ρ��̊u�A�@|eOT���N��R`]:���f��+]���.�Q�D�ՙ#5 ��}�.v�/��·�J�=�]�j(S���"��xz�J�R[Z����䛬�ó��6���2���l��hͼbtR�ch���pn~�t�q���G�X
�u�Dgu�`�D��}����ʕ+9�"�յ�}F�o���_~�^��~��Xx�83�~/���&M���Ä�߼�������o���}��w�˯�AI��ݹ� {�Ro��|���S�M���_��yQ>��*0�P���:�N�u�m�p6��+V��FT��q�n.�	u�U�Zd*�4��
��!�,M�L��i�F�e01>y�����:T�Fy����QfO�:�Μ9N{;J��v��\f���6A�E�(Y�㬷ǚ��A�'���ѧ��O>�8�s��g��x��H��*[�ӑ������Q�z�����O.؞�S	=���%W)w?v<{�T�>x�}�+Q���O�sJ%m8�J�%���}Bf�i+�+y }��C�eɂG�+Wx����8(bX'������]^]Π��|�SV�%�	��^���!3W)9iY~�E��Y�Gq�i�!o����o����>l��`v��7u�^30��L�e*����m���}P����CKC��.(��|G7*.I�]w-�M�2�Q��!�v�$�t���zO��3��I�X�d�0ţ���Q_��0h��/�����C�$��D�{���ߞ��!��=}v�I�#{e*������}�)�C����`4vj>.�I���}���8���4���8rU_P��E�6]�T4o!�n�x1_
硕�a�xL�����Nv3{ �'5G�����NƼ�W�״�ҥL�d��5��'��c̡�G��:�"w(ek�;~��:���o�v����N�)�M��"��� �7~�vթ�����?@��7n�M�vt����!R�C=��A��v~�Ž�*h��F��a�k���|�|�4��q�~�M⨇o���o���6��tt롍n~O<q���o�o�ߑ}�۞�ާ�:��\Gt�F�S
>� 3.��dw�_����8,'�˝�[$hL�t�/��cQ��r�o4�0ۄ/����PEQ2%�.��.x[&�;G�rd�ĸ6������~��P���̉�ئ��Gf=�f�B*�'k��Y}O�z����CP~;Ky�G:~���E!B�r��e?�._i/\�贊���
.O�<ɩe��e�� ��g�Y&	�Q�w��aW�2�fĻI��9� I�(g������wȈǥN����>����J�d�:����Ε%���P��@y��b��$�q�o?}XE��c�|��I^�z䈳
��1�����G�U?$�JV�p1�i:=��I��o����R��mu}%եz-3*�t���,���쑸�C ��6�{�8�R�c��Me"���z�ql����E�
����Q��b���h�Mx�4��y�&���������~�E޽�̴�9�g̒3N^����BY��y'������ɳv�^]���3���������/yo*�SN�����I9u�l;v�(�G�K��3qK{x��[�=�>�(�@�/h3nʟ���=A�(���?b.t�ezl���}��
���<�N��N7���u�����~hs�_h�z��cm����\�M��oܞt�r̓ԉ��>�Y��l��m�ȼ�޻(�5OS<w�\��'��>ZK����9<�[�;L�d���)HW�f�8�]g_��#x)�Gќ�.�P�~NL��.Av9�p8;>A�����yP��zx���(gy��\�<ޥz�f�ܨhѴh�E�k�.�Eɂ'�L3�Dm������n?PP}B�σ]e�o��wQn�����pv�uPQ�Di*w�W Hct+{�=�߈�g�I4|�J��}�;���0���Oށ�C�L2f�u�&q��m��{���ԝ8JyR�������Cw�%~t/��zv��y�O��4m��(��?Fʝ_�����.��;��#?���*5��0���H[������*�|��t�$�&�V�>�BwD����m�U��W!�i%6����̀�1�U��F�r��6>'^gTp&q f��Nt|�8&7۫�����!��>�I�S�<�{sM�MV)�����&�&y�v���J�L��}�|�߶i��n�}�)~܃�:�1���a.�˱��:N���0���|���{%����-Y���Բ���a���r�<ID�e�vo�V�W�گ���ܺ�������7�@�^�q
*� �!Ա� a�`�H� ��L��C���M�6&"r����1����[����q���v2H��'3l�ٙ`/�FNGM�j����t�T��ד�0ELt쯁W ��%g4p�o��/�7��`*ݍ�i�@p
.�PLp�{��UQت�\WA��0����p��{��T\�J��K�q�����ٗ4)����{�%�2��s?e�g�S?�M�m���^&�oӎ��O]rA�Q?�xȁ�0����W��V�W&5ME�S��R�H{Z2���p�����<�5� <��ש����84<n���(E㑑�~PV�8��$�uy��l���ew*>���[k缿��v�a��6�������Ѷ��rt��fp�
j�S�����/�#����F[APx��	��"�|	�@����JH����f�ˬO��l"8xB���3/��������v���v�������ҕ���p؍��O!��R@�}���>7׷�SQs(�޾�>�������S��B���>i_��=%��<l�o\o�n�Dp]"|՝Kж��{T�ӶI��}Cy�P9A��7��6	��:8֦��]����X�.֨w�D<��i <��_�e�����~���x�r͐�mA�����c*"����e�ޝ�9�̽ ��=F���Q��n�I�W�%42�����a��;6�ViO�H�df^O�=�=;��,c� ��	�CzT�.�}�"�=|H��Wg�<$#ˠ��$�˝|�%;�6�S:Vᙝ=��{�����~��v�ܕ�ۯ_������A��Cڶ�KiD�c\.*���X��5�#�CGY6�f�lc���sgڻo]h�/Ϸ�'��mkǏ�x�|�]�z��ዯ��_}��?�ߖW�{���C�H~&P~<`�M�[�eus�-#�nPn�&:��,�|lЮV���Fl��W�cx�8���g��j�^ZESC�����MS�ơ�#����6=G�'�'���Ĺ��wpM�*|�K[����
�a+U��v��v�⥜H8;?C���m��}m���.n��֗hC���z{����٧��޺���CC�z�xm߂�thn�M�җ��֡.�d�fjj�d�?9ێ�8mɒ\���h�;�f�t������������3�w��2�r3M;8@A �����'OҌ�]@��@��`�{����q�d�o�}�+d�B�y������Ǖ����v^���h7�ߞ>}����8�����Q�'i_�q����=@e}My-��O��1+�c��ޑ��w<��0=?S�4�J��)ڮ��F>��ϋ(���ۆ��Oߡ\�!��_~� ��l���jiqG�£�_y�������� N�
�Vg�i*m��?���"���S
���O�!��w�_	)m���jHP����4�JL~T-C�XS��|�6�]MF����x��e�绲�^�1���Ol� ���O�$Pe�}����e��2�E�tC"��)����~����#��@qd ZB�a��/��jp8_YZ�6y2�l@�O(���x��	��R%3aS�Y�Kt�� �6neM^gd��w�p�q��h��=��X�܆��2��N��mp��݌(�[�L�4ꌠ�$��nm��
C0����F#������)o�f4�C� u��P��$�Zr���[�%�K�*?3*������w���T^��Q�.Q !@޿*v�Q,��z�~��q�7��uԵ*N�������@.��'�
�`�=�)�n�H���3 t�@�1�QZU7�3a�ګ���B�N{���.a#�"�+p�/D���e��V�t/0�rK:I�
�O��,�H����o��:$�n� 锽����w �1�O�e&���+~�=��w���^u0��J��;`]��ǐ�*�E�Ug�f��o7�(��E<�ҷay-"�w�V�\�^I�S��|{��\���
��x�]���Nx��ޞ�� �C���d��}8���؞@�������L�a�my�[z�v�Mۖ#��gg�lWB��tf;(��Y9��6�z&]��%��U�害B��_�v-�^�~=���#��N9��ҡ3��d���gQ�<��X�n�p�b{�w�G��}��g���9��28Kv�����՟���G�����)�[� ����TYK�m���N(��[��>�%�F�����H��d����i�x?��s������?m��?���_���={�zP�nI˲��l.ut��x=�)¨��*DΚٱ)�(8�o4g��Lp���8U�)w���w�i��������c��Ge9Va�?ʧ�$�����尬��l����?�Gg
�c���^<_h�K��T��D����>m����(����t�.�\ݓ� �3#�;�R���Nڛ`�ձ�w7l+t�4���v��9��C��q{��w)��зeYY�i���k?��c�����U��{ݜ���Ӗ�04�i3}4�`B�|��Yۍ{w�}y�=������[�>6�w�W�K/T�,p�efVE��P�l���8��*%����a��<o�_,�U�{����g��Y����~����(�����=z�rhr��<~:��~��Oۯ~��v��9�g�l�ֳ3�;ԥ�)��~g��yā���g|�ɣa���N�!|��h\ҳ���i�33Sy�u�����m��K`1�'�;m��΍%pݩL�����{(�CC�&may�%<`�������z��{�6���Z��Ç�sO�7�|Ӿ����ӏ?�79/ﳞ$�dJg��҅K2�e�U����Kl7�S���hf���l���4a|���,�<iDJ=֏`�o��/L���K�@	�����޸�.+΂r�]{���cT�K*Ƙ̇e�_�6��A�ƫ�lӃ�|�R�0���׼ǉ�YF^ﻼ�M0\��� =�<{>�(��y���8��?��Y폾+�F��3z�=����2x��f٫����O�x�o����>�C�gx�o��'8̗�<Y����#3��俊���]��Ĺ���o��_�{�=|��^,��u�<���	,�X�������8\,s0�}� -FHSA \^�S���ݎf������ W��]� r���v���v���v�X��P��X�4\U%l��6�8q�-��	F+��0�Wm���c��^�I�&�(�i�����H����������RXf��/� d���¤�@;�R����o)(ƫoҫL��~�SH�
����B�ݸʍ�ߍ�<����'�{>���+����^{�V��\�~�N�܀{ ��3�ݴ�~���00��9���n��7��8��F��z1��i����ͼT|��0���~*������ˤ��.����� $w_e7=/ �@&V����y3����K�3��mP؍+���;�X5���v�{f�F�`/ba�6?�M�i��C��t,OaZa6K��O|� �~�	��,�}�[�����cS���S`��d��a��Ky|W�p��ĉ�(��Y7�=r$���?�;e>z�^.�-�����Wک��)�ʛ��w<mp��F)��U�� g��g�M�e�Æ���4����Q�i�ҥ�mfz.q���������([��/K�B���o.R�;���a*�*^.�\�b�'���g�*���lއ�}W8r�{Y\y�I��W.�?��[g
ފ����r��\¨"����"�Վ�8�:R�{A^��p." �@E؄V.3�	��}�t�bJ�Yd|*u� .\���47GƢ������ٱR�}�%!u�;�g�n��ޠO�0�K�;
ݡ�	��ʛt5���cs��R�O�>��+�5��栁K�ܷf��o�y���d���m .��2�Ai�{��	p�v�쳏�/>� ���F0�|��Q���o��_�~��j{p�8Uq��h��G����
ޑ`�ַ��8���o_i��V;s�T��� �
�mZ�/:��{����B��G�=��z�q^��g�q�x�%`�ݿ��ݹ�={�D��n=����i˚��:k�&.�t��3�V��m����c���o��.>��%��O5y���A�Yo��=�^�o�kO���I2�S��I��6x��1��P��M��@fz��I�p_�xuU��N���65��:}�P�iy��u_��M��B��������J��tV%���r<�����.�P�t���o8=U�e�ڣ��#��{�n޸�nܼ����>B�y�]/�����w��=y����K����uE}dN�#�����mzf��:y<�8��"|�*3�Y�|�A��5�/�re˘KB�Ļ�H���4^�Gk9���6�G�<(��
���}!�!��h�S3�/_��f�Zq����*�����x�w,#�[܇�R����~+��3\��>a_�(����>���|��8FL�=�o�V�޸����a7-���Ob��3HX�w|a���u>|+{�gߋ[b5���0��88�=~���WPq�/ȯxT�H��g�Q�~�ߦ����o�?27�N�8�Ξ:ގ=����m�������݇�v�,�\��r�R�2�0.iW�A;�%+Ģ��Y �ҁ3O��A��5s��&JL��[!Ŏ8'F���P�Bu�ıv&��6h�N>,���bu�B�J�&J���k�wT�C�Q�`��[
"2�!��ݮ�!�ש �͟��C������123�G�"���}���4�6��n��`�(�Q2��9�Gy�fi��A���V]�x�i5��?f)A]�a�GBy�@�0�Î^<tsH/��;de��s�O�:ÌB�)��=i����Y���<�H�s�L���y�R��0�iP)6���-��0�$����O�/���ӧXmٌ"��?�F�[O3���D�x����K,q��_�
��z5.3\�f�S�J^?u�~�c>Wu�/f��s�*���l��5�O6�!��Mcz�(
�!x�̡�g?����(�P&��ٳE�N�Y�3��9�5y��xh��|E�Q�r�����Q�Uq��
�����Oڽ�w��x���=�F��;���2��w��aXe�2�7b��8a
�������q�|�;!'��<u�L�'���u��{�����
a�F�=��ZS�"}�Y�hY�3gϦ��W�kޤ��OU���|��+���e�b�#�]�t�]�|%ʕ�9'Nz$�!�����у�e���"u�?�}���R����/��@ ����ٶ}K�\>�".n=<�6�|z���u���}י�������8���9��Pጲ�8�ag�:�"�6�/Mk��ZN����*Z�i������h���NU�S�����(Y��*�����d�)�^�s�no�T�d��6�.^�Ǐ�>|�}�ه(X�K��#������r������w�?��<�>�	K?��(X�`�h����(n�a�����g���O>��m�0*1ɫ�-��x����2����v�I�*��{�]�t.���'����1���ݸ���(
�a?ʾ��8{<�ջ�����q�{
�A�ϊ���z��J�����������>���u�4�1
�y_Y�h�<kׯ�m�}w�]��F���.1ևeA�:��v�J���57q9b��"�<E���g�qP�}Z�P�����Uق=Q���D�'�҉��e�*G��5k��{�{5����˄��� *P5p�B}/g�ʁ�+�z�� �z���������^���,�Gt��[�?���<��������={�B{���P��'\(&���mR?�(kgϝξ5�<�м9�*�|���b�b���d����2\f	�Kd�'�Rr�)���ӷ�a<��^�x.�=xڻ�3���wQ 1�="��g<C|��w�V@�U�������.�ߐ��נ I����[N;� ���
S��q`p�U`��]0��f�=O�1��+�LC{O�<��G�P���47�)�e��"�^OT&���_d$+Cs@h��䡊�D����JɪA]WD�ͺspRoտ�S���@��7�d�9u��86�!�������������O�ç/ۋ��R�\��
N�3T�'����VFT��r&���g���LR ;�*�_	3V�rĥ`��^���Yz��G�i��;�{��	������ѫ����|QfS���T�ྸ;���������:�(Y[m%�۶��K��ku�Y��2�:ũ**�ĎwM��z��@=���(�d�S��ɠ��:k�S�.K+���Ž��|�3������o���`h�!�$�ᦿ�ծ�n��+ T��r��aI�F�+xi0�(��#T�*S��%��cʞ2��^�!��0�R�_��e��R��ۘ�K��k8�9��G�7�*�,�^��e�ғu7�K')WL��r�W�A��UO�@xBe=n�p ��5����ػ[���x�O�-�(�p B7���a��|7|W8��|G(�[�Ǆ)���f��H4�ψ��(Tҡ$�K(S�r�q4������՞�;��S��&���Ħ��۹�g���ۙ�'�g^�[A��)�(g�T\<�O%�2
�n�;#�B�r������}C�n݌а̻������,�m>d¦��J�-Z�&�1sH���].ݺ�&�珴c(x�Q$N�g�p���#���r�WV�<���/��`�C�(Gǥ�X����U���Q�Ӯ��e�,.D(�xm
����G�ϱ��y�p�و��|�x�b��q��2��s��}��{����K��u�6zY�ʖv�}A�}M.CS�VYqT��yM�XY�]3�.�<�ru���a_x���Q<''�7��ʧK�AW�SɊ�	~�8Kᥬ��43����D��R��Џ:\��l�W��i�Q�)�����N�U�ө�nm��挎����Z�EI?١-�����$�=G�����~��O�8\�p�Qalm}u'�C����?�����_�{�}����� �+O<$�V������mU�w������g��%��	�Ñy���UOĵ�4𱶺J���`����#(W�Ϟ�R���(§�GirY�`�6u�]�z�=}�|�~�G�0��+~rj��i2�j�_�e��=�~Q�p��)��?B!�X�h{��̐��>�P:ڷ�\m��_�?|�M�z�f{��m��"�A����T�:{�,�ө��쓋�uZG�z�Rm�/��d!x�LM�����p����]��K]a�d��b��˗y���
�~����(�GQf�]��(zB.=��z��Ax��e˙�Eں��Q���n��r�������ť�����v���v����Ue.<���m��j6���S�ڹ�dy��3��A^Y�R�/���ۉ)�*%K��s��m�!H��Z��|�єq$�����E�ݾ&.�$�j�	Q��G�ݝ 	���Է|�� y��V=�}�}��r<��w�q+����G�E������û�gx���6��'Q���g�[=#�?��Oi��I�gd�fw.��� �.s���Xq�񻟌K���b����q������ȫIO,�k8He,����n4�?y�H;��u��� R�����տ�뻎X<��.���M�c̑�QI�Do'#�0?N]g�/H��Q)|�J��dx3f'��ú��f�\?M�O;�Hc+/�T�rY�&O�q٠G��!`��<XEώM�sSk)Yn|��hmem���\�����(W��HP���A����ur�[�T����'�B�t@�0��pv*�w�nu�e*P?Ɲ�_̓�2�
��Ox޳�5��+@cV�P�2n�4B��?$�*��{����x'J�7�R6	���n#+�����������,̧zO�q����{�L[��v5��{OC�;(��@����{��{���ޓh qZ>̚Q����^�\U�(��ow����v&��(�-߆r���%sI^H7f�{�/ܪHE���Y�ҭ�/nU�=��;�?=L��aP�Rf�<�6�7�T����@��<�m�ƅ��¡@��޳�x7�U�U����슴%�����y��S
�.]�7�hթ|�Ξ�R�>"O�;��u��%����P	A�Q���\z�]>�ݸ~��eX�G!�fRFx��*�휲�k�d�V<��y�|�~�WJe���9��l��0JeK�t8��&�2C��0�<��o�`=~�8���%)�IL_C>�3I\�Y!
��L�݂�GP&QV�n.�W!���/��;���{��J]�l��w���K�έ;��@��gG�8ሹK#]��a/m��`GJ�'
@��̒����E%X�����G����S�,VW7�=��~�ھ�����ի����iY�?mP�QQ؃,m�ࣀe���2�=$���J��jw9�Y�j~޺m�Ay �!���{�VQHd<��:���ɶI�d�<`���-�K͎�Q_�x����~��Oۇ���}<ʎm���B�ķn�,\��Zh��'C�^��ʓ�P���O,��&B���Z8�D�c�/���\�rt��>�h���G�4��,[Z^���e��(t�ё�<����{;J��E<ua�iy�~��:�|�=}����fP��*cX�	p�C� -YT
�yr�Y�H�@��0�K��%�Sm� <�"*',,,��?�n�7_��}�m�����ZY^��`�;V�qp�vJ���r��6GU�����/����d=*%�r��N�f�Q�Y/�Ea�Omm:C����!;O��x �v��-�haJk*Y��\	O���~|��r�ʺ��`�����#�B�l!ˀ���������1iN�(�<�Rf�N�'N�g/�=�t����G�%���9�80S3�������,�<{�6z���e��^k��y:䗋��ey�!�$�/l����6���d�m��dk��z�w�گ�=v������_��aj�
�[�_��5���ݬ��Bb~Pp��߄�;�3}'�=������-�(~�K��>���޼�[����<ũr:z�睧����^y���WFbO!R`Ͳ'f���~��>��"��3�`H/�t���~*��Ğp�я��i���O}�R~\�� uy�����]S���1�өv��|�xf����].�������G���%�ā���=Y���Ͱ'�%�޶��X�?Wɲ���n����M2"�T��r>+2��	7�*Hx�E)Y�&g��1:h��
���d�6R�0�R�L��/��k�VQ��\�ȜHB�>"R�&G3c:ZPGJ[���1HEXP�����~�$l�K�i�Tu������վ->:ZJX;t:)o���ݽl�S�	��zw)��`"DSE�q����i%O�=Lf�d~x'z
PE	/���z$iA@�/r�=�λi�ȿ�������H��Z���7��_���ၤ]y @�!��40�r�I�")��>�+���u�~��w��C����U~��w-|.%eG���42ԉ��Xm>�^i����bO`�+bK��{�5̀9BS�Q3�gR�~ �wp�b���ɏ�%�R��58|/3��I붻����uS
U-1�YA�'}�Q8pψ���T��p���W��*����l6GY�nzfP&�?�٬�O"�����.s�Rރ� Ð�ďЌ�����M���w�dI��Q�&|2�����7�v��h�2�.�Vys$�%>vn.�sY���{~
/��#�U�\/�ri�ݽ{�}����{�+��~�p�"�"*~���^ �&�
��ˀ
���\�73������&^Tl�wɃ6\��e�*��U;}����(>�RQsf��{s�~�m���~�n���
O*��������%���!S(�.����p��ԽʆJ�iZ���(�$q����֕�P�.�3g<
�X�i�=�����9��͛����ν�����R=�#M�V7���q�o�'u��S՝�].�@��)m9C�L��d���ޯ�Y�>��������U�#�X�:�.j[ѽi8𸾹�������S�a����PoA����J�x����{���w�+�c-��Gg{\*���=eGQ�=}���>(��eӴmy��3��O8{9׎ 4���D\ui��t5m߅gsrߙ3�h�ҞlShg���+��[�^io����p|xb�'	{��Rs��U���s�m?�hW�=������yL����tV�� ��̤\�r�]�t���ܷ��:���������o�M���~}��,�F�ٿ:�nr��K9�?t�,95u���8�8�r��U䥧�Pbg&�ْ���PhS(Z'��gt�(�����S�x���9+�]eJp�T�X]��)ʖ��TV��r�ji��0J��7�U����F]j(�r&,3W
J �Y��>^m�uG��?r<<��p��v��
]Bo�<L}�]��\�(Fy<}�4�j����IҠ�H߽�κ�@.��9��r�Emڇ����ٖ̜-U/�\��=����6�ǴȀ��Lk��9�|�O�����D$�ov��wdv;q�w������Q�ǟ�e�����2��w0�s��#J��ӓ��d~��{��`���S����aO����'�Cd&��LS���wh }j��Va;�Ry~J�|��m�ۘ����)e��)?����A�~V}C��ϜW?���jʳ�Y�(Y��S��v�4z˱�65�B�ɺ7ړ�rA8��f�Q\�GH��Fs���W�f�G���#P v ɘ
����^^�7tnG���
_vLnH<����	�"�8�������EgEX���>�zW�6Q��,���:��6�9�bǐ�p����P�c0��q܅��"�h���1�^�
S��;�`F!1�/S��Q%ܝ�B���)L�.�s�v��1�9�7R�H�U�����O5��{��D�##Q�Fy+.�+7�K��n$B�ԓ����Nq���	���9��#����R���Dy(K>�?�'>��<��oډ��a7�x��}���S�kbi��%}�o<�{�G��ɿ�i�>����G�Q�z�IK��Y�0I6�t7\��h#7����(�0z��W��aV��^��Uyح���M��Vfa�[�^��{ 
����/��x�c�K�&��pW�MZ�)�2s���4bg=�	�Y�C��x��m�\o�s�˲����U.%�VFІ%c������s�9bM!Gah)�z\��l��N��X�����������i����}��x��±wg��b�|��
���:��#������`�믿i�|�us	г����ViO�~޴j���,m�96�MeK�i��e��s�T��e��2����Lj>
�»����Mަ"����(7_C޾���a[�ҏ˹,��T!|��E��B�l�3X�@O��5�8חt:{�L��]"9z4K&U�ŗ]��xɮ#�?�t5
֝۷����CA^��K�/�5�>y/��o�рn�l&�ڲ?�}Z�(�Kշ��D;Jg{��ցCwp)�˅U�Ut���[/�:<��稇�(X|�~���_d�C��5�~Ӗ��W��Ӷ'�zٳ{^^5��=v�:;�YYg�ٽp�<��9�u����5�i��_|y��$iY'3ч�o��C(Z�f� uv����ͣ�=��zrfϙ.3/̾�rxE�����u�d�Y���������B��i���n��T�Uְ��P�+gw=t�-hT��;H���/C�'��ǥ�c(���e�z���k��_�}n�A�JMQ�S�a��Ӯg����B~<�b��#��G&�v����v{F�޻���v�rC�� �f
�8}�X;w�d;q�8;��^�k���O�D�FaR!��A������\r�=U�G�~�RJx��YYJ��љ+��zȅ3���	�.'�,�:VY���ٿr��,T��@!wf�{�nݹ�n�6��mu!��鸟�~F޼����'P�ϟ?�.BW��2�M��h}icf~W63�m�������"O�˭L�#�Կ�ms��0������sP|�`�W����В�z<y*T*�[���������R}q�O��L�W��	_΁^���F�%"��2 ���;�6�{)�䧿w���6����
�t��<��E��o��z/����'��X��* &P��Wю�~�@�%�d�{O���-�����P�)dʲ���զ#HG�����Odfg����P��ǜ�P����5J��G�ۣ�(YK4�~�E�g�MBT��#h.��Dɢ�ڈ�ɪb�G��x��J��T�)D@f�|E�!v��/�����LjX:�{	��-�o�k��r�M��E�r�{�b!��<
�;�]�+"�襋��>�[4x׏���3������5U�r�k ?t�e2�I~��H�6��Ȭ�D���&n;�?X�V�/^QT-?Q�����zѣ��$�VMx�7�de��πՑp�Ks�"#��:ȯ�XDX3E�{�*w�=~	?E���c��:1�0<j���r��v~�T��hL�n��C�ȸq������[bK�z�QY����^���{�k��J���˪Ŵ��Ѭ�(��0�9vʜvRI%��/��n~���Sy䯘�
����(��/~���\�8�:�ި3��)`WAf���2��~8KpP�4{�QD��{�[taZ�SPpP`t?�J��갱[�ǁOӎr���6P�<����<����a@!��4%�JT�eYn/^,d/�����C-�q���ϞD�Q�r�Y6p#�;��~�y/W���
��ݍ'V�n�(�g�;7���iʎ�V�W�2��$ۍ�7W�^m_~�B�U��4������?iTj�g��{�s�2�5�J]A�69�hq��|��	�=�������7�p�K˜r��N����wߵ�ׯgF+����*����t#��7>��y(���������ʗ����8�Re~ff< �eF��H���8Uܜݻ~���E�)u�)k�Kj@���ށ��0w鿻�hi�a��xy��+͚�ֆK�\F��xd�����I��8���;��C�Ϩ��$U�	��1���.�|�����﷏>�����ۙ�q/r��� �'��w�5��S�~���j��S.�=y!�|f�<���[W�:��n9�	c?�>.G�P o�������Y�З�e���8�x�%-O!t��
���\f]��ȋW.��9���o�:H���?�p�����v���������J�jZ<�@Z�*1
6Ό�6<�Σ��3�9���(�'N�f��>ys��{�F���k��v���,_s@��8q)�`�F�����#_C�kQގ�͑�'OΖ�����§�_R��۽����� ?o����Ȟ;�NK�(7.u���A�R6ڥ���U�2�Dyu׮��z���y�Q)��F�g�t�h�u|�ʚK8�
(Jҙr��>=��ҥ�����x;���o���(��P�oSG�0�����~8+0>g�Ϝ>�e��(���}���[x)߄�³l����l�G���;�&�/�q�>�n_��^� ���+>���7�_$P�啴\M�(���U���gc�ϟ���o��ߞp%�T������O=l��2����0;�[�������p���}/Ƚ�_����}d�%)i������}���;���C�����7�×6`�/�2L�Њ�L�S�~�S�q�I:�`��&�~�p�G��t�	'�;�#�*����v�ӇN�#��9���j��k�P�z�����%"R`�W��v*���;C;�,k�!zQ��N��?;L��P�(�>��IfS�Y䩐��2��������E��K
f:� T�`�Ƒ��j=w_x��#u(^���U!$B�3Aө�9U8�Z9z��'��
�A��:E��|� +��������T����$M�L�,/���Ly�L��{���Ф���PѠP\f�k�2R6+?8���wA]"�U���-	S����M�A|�t0�C�|�%��
0��|3�SH)�:M퐮u�^6X�6�y��p�kf6�đ�B��YqT�����=�� ~�W���?�>�٠����i�?��:�u3�G��wq<h�؝�.lM�X��a"�f��jg�|'����r3�Ą=y�b�8�\��JV1���ed�u��6�C'I��Y�4���� C��*�6J�
Vu����/s�@)I*L��8���PhE��X���O����,�q����s:z��<|���a��~s��͛�r2�]��5������ɓ�����B^A�ӽ�TR�ߒ��U�t�ûe�Y����l��N���Ic�[���p�0Fh��Gp�DP|��<ܸ���72:��2f�� ���D2 a�QWҎ'���[.����)�iW�r����i��+�pO�c�Žql�W\
q*��S��˯��=`�ZA0��|e�e�$Yѡ�as�,���3�S��r-g��m�ڀ쌼���e}�.|V��LG���������Y6�>�Foz����z���.|z}��'��ʹYM�L�n?X�*��H�s8��VW׳L����9.�;����S�hE��rQg�>�����+W��(8���-|�T�U����i�.?�.�����+�w����[o_�2���ɓ�T1w?���@�i�]W�8S��5��e�b��k�@�2˘�Q����X�UG����h�=|��˼nn:����'�,��o�3�N�4ytz� �3<)���Đ^�����:��%v**�s�|v�>�>մ�"2��8ܿ��}������]#���+�Q����襶��i�^��cm��e��P��uϟE�<ю�O�dN���W���v�0�G����6��r������ʥ��4
�a��j����T)��V�GMiºt	����&�;H$>�]U9kɨ<c#�-z���Y=��0�/�ص��(�q��C?4�R@� �m�� z�y�~�s�a{��ef�<�b�O]�����Y*x��ɜ�:77C~PQ ]����u������aO���*��X91��ч����ه�]�W�߸��}�GR�H��W~S ����S�!6�F���p���wO$���-y@�x�D�=`|���$s�?%�`"�4���i����f���0��Ra�ɛ?���=O�՟���!��������{��}�[�S�T?Zv��M�z�ң�[:ȯ�F&�n���O�|E�$���M�p��� �	;�"�J����;u<�θ2mm�_����_�{��/��d��17����#��6J`6���U '�@��5 �h<a�(?����^!GP]�25	��D�bn���Y<v ���3�2��U��~7	�.B	���*~�_#��T_�4o�_ZDP[q���"a�мfP�).�k�-��k̶�� ��{������n�tj��@��m��Qt�E�-��d�B0���J�>`���}<&��f����*iM9c51�&���.��ԑ}m;.]42��t�}��7���&�o�q	���O �8����4,��
С$͜j����kAE�w�M$O�QGF�ﺊeB��Zp��P�(����[�"�N�<A8�s�x��qG���&B�~�"��*C��c�9K�0]�y q�W� �!i�ka?i�q�%���?a����c���cϥ�B�B�	S~��t��mc���Q��Dc~�Gwgm5�&H���x/
��s:&:�I���hw2Z:�����%4Y�*>d
��2�$�F@��蒮aE��0e$��m���E����C�5�S�b���@Յu�L�4�(x�/�[G~k��B<�x	����U1~�5y��2m���m{s���m��8�����G���'���O��0U���()�mw��l���@��� �ߧ���P�L=QI{����ٓg�y��yF�U4�jJf�:��X�����������Dq�N 7����^dy��$x=����{m~�����w� �_�	b���/�@A�t�!w�H�,8�"^�GI#�ܰ��Qә���WV�ڋ�_g.�Q1}a�����B�S�{�^N6�T��?]��j�͏��r@�[��w��V�p��S��XQ,���VW<�|x>^��'���G+/ϟ/�O��m���������߶���ݺq�0ҍmJE�%��  }�t���P�G#��!�0
R�HmD	�^]b>��k���9�uv"u�W˱�I�/�(W�Y�DϞ=lt_���:��┙ڢ��b�O?o�{%�x��;Hߦb�Aq�k�_u�������ٞ�r��iO�<s��?���l;yb�?�B�@)<�Hrf�P�b�D��εP+(�=ӯ)�g������c��;+����gИq��N�#G�4Nt�Y|��������~���ؾ��t�i.��O�7{ҽyu�RV��>rq?J�+3�|���E�|�=Y Ƀ(�.;u9۾ܑ�E;X]ބ�_�^\^���4z�I�<��0J�4�~EeYŒ>	��28��)ʶyg�<�Y��<v��:�rat�,K;s
�Z]s�}\�w�}�����w�BY��rϔ�r�h#�#ؤR<Y�A�~���R�j6Z���),n*Y�?^���:ϑ�p��+_T������
���	�Y䫱��Cy���;c~�n�q�^{ \\��I'�t�{���f~��L7D��(w���k��2u�H,���ǲW�.��'�Ki�=l�����G��@wڢL�~�6�)�J'��j�
�"(	؆���=�n{��]���G%W\�$��72��.��$�7���<+���F�W��7���	�5��ӡ_+��ɢ�x�§�{���x#�)�a���k ڱ�x��s�� �;��v\��|�:����Vo  ĴIDAT��81��
����T���W��H̖� �p��WL�A�����t�ᇴ�e3<PuG��IVYMϙ����K[���k������Ə�CN���峧Om'�ε�䉶��?����z���tAc'�jػ��R���6�itg�ҩ�P}H�i�f��a]�'�yҗ����=�i���ˆ�؊iW''Q��e������fl"�������E:c�����A\����A%�LMe��7"�,��-7���<;�t��Mn	�P$q��Q��K����� �\ɽ���
cX"*?�t�n�0��=<dܡDQ�3Ssi�wl�+���~���I���pO:I�o`)�HNk�����3�^�����I)!�B	�*\�|��P9��!�!4V@GqP���/g��t�e	��S��=B8񍡘d�μ�^�>×���7�;rlC���Xt���\��8N�hd�1������2x��?����V)F�N�t����Ow߆�$\�g���w�frp���2f�uz�|��&�i�4��N�������V�c{r&���uf�wE�n��\n�?���a���m�i�Z��l�N3v�O|��Y��Y���"Ĩ��hq���g���q�Љ�^��p��{͇���A�Q|x�B��WKKG�yC瞁�@,"��}ˋY��l��<2C#��DHfn\z� #qy�M���������W>�0��3JW"�G%�Qi�:8z�2������rq+B��t8 eGb��a�|����˿��`���1~�,���pxj��;wr���[��-Ҽ}��Ӷ�,��n�n~~��'�ֻY~�ި��)3F�[�@>�S��ג#��I�.𭏗ԑ�ڝ�(�����1yP _L]��Ӌ�M��������ŉ�Lڅ��s��͌�`=��
� �?�P��g�_�q�.�Q���P�O-.-&�?|�c����s
�
�xs6 JC4�N�̋�^�|���vd~6����o�C�+��i�\Xo/�/��p��l2=�%�.�(ȫ@ll��ӭm���J3gN���7iց<�e��	]�M8sI�C�:ۨ4q�� �SE�%}.w5,܇�*��"�[& $@ۿ�^ܫ��,֭���+�(�of�t��>��HW�{ۙU�v�N:ӭgєK\ƻ�esk���(s�����о���,[��������
0�ٛMG&�x��ǐ+�8�w�d�؜9u2����(z���w�f������ٿsgO��޹�._>�f��m�d>��V�?�~��;�X�-_)vbXv���7ͣ��%�������ʷ'�j��ҁ����"��tXA� }�t�U
+k�=�x�}���[Fyw�K�|�~��ɢ.	� �З�����w2k��U��R{_X�����tv?��c"��ɯy���PF�Qmq�M~���R�_�
Wv�ѯ!E\x⡇�����n�)'��n�Q�j�7yL��ޡǳ�|������Փf��7x����4����O=?�/N����S�!Ϻ�W~�Wn�V_���y؍�?IW�.O�xU݇�e�o-��h�G?֛m0^���e=��BB�OÃ��:Ǐ���{g{��|;w�X;u�H����2�����������ŏwڵ�/ڋ��0�6	�t�i[9��y�����((�/`�K���Ȁ v�a2BA�#D��� x{4�a������m��4a��9Ҩ`�KaNS0�g�mjf��z�~`(�h��`��`���@��c0l;�5/�1�;R��8���I�� �eZ�0=+�N�NSSw�"ah�uV���QMAF��g?�٠�U���$yFU-��ܢ�ԯ�g2���9�wH��a�fo���W(�b�gH�p��A+\�ǝVˁ���Wi�
q82���"�+�!�סE{tn��2��~��&��}L��d�U΄'GM�S+��xJ�������I��xU��>XN�ոM����,�F�K�T~�����5�\e-o4�ġ���@b����|2£ɻ�%
"���|M���v��hG�U�ܟ�}4*�~�w|�'<u���sJ ��vZ!�H���(� �*����X��w�e|������=~0�V�K�ON��3Jn�(��Rn���q<�\m�-B�/���M�y��M��2>��ZYz��V��:|d�)<:��������m�-·@!=�g?�Nϫ��"\m�<E��݉�zU����8��������`Ғ�����P/��x��Ġ��eW���+�Ԟ4�(aܽ$&��ym�O�'���G87=����|���[.e>����r_�N��썋�!���ˡ`�iv��`yZ�JZ�g�&-���Ꮤ�64��x�C����Ig'��ʲg�4SW�}`�>� A�Д{��@Q�<MPS��:�poI�#�=��>R?U�g����)fF�[ ���+���ȇ�ɀ�4C��7Rҷ������>H�?�jG�m��#��6ys82��#T�m+.����Oۯ~�^N��ɍh1h�Fp+~��9[t��K�Q=�}1�A�������0��0n��`_��=x��]�q�]�v5�ڻ��[�Ҏ8���Ի�?��޻���N�t����I�*
��P�=J�a��Ν������7ߡ|��NgY��MiD��.2�@����>p�Z��Q��O����ގ#+���<��t�=�;��Ls	�̭cc���[!�KfD���ω(y.�t���&��+W.P�������?hǡ��{����/�n_~�m�v�n���eʲӎӞ>x�J���y���w	3�z�n������ȟ��e=K��qL��S�Q�*���y@���Q����0��e�
���������c<*�қe=q�t;z�d;��9u���������ﯷ7�/���9�o\������ydn�]8{�����v�vhB�mf������������my�>yj�|��d��U��3�?���{���gm�Y
�I�'8�~�����~O�����^r[�x��_^�[=���������{�,�_���=r��h���V�ݝ�$�����^~���7����'e��o)I��<��n��>{��e��i����l�B�Ѓ�x��F��Iچ�&䣴}s2/���ޓ�x�n�e7u�=g
sm�dp�輒azr�]8s�}�����O�k�{����Ӷ���?��w]ɺ����=_V�B�o�¸���Y�,�z���@��r��>(X���tT�%:�F�z�F���D�Z��~��I��xll6�+P8*����t��s�0��Y��>,GgM{��7��T�@�̗���a��T���W�:Lal�c(^�9qhs��
r9�4����6����H�,t���4i6qÄKX����J\�����N�T��A��,���c���{���߹w��u�'��QVG#��f��Qa�8�b��k���ҿ��ba$$��q�Ybf��c�O���t8����Y&*�ӫ����x͔����-3Qx-��@�i*�\f	�.H�v���0I�+Y��M:�#,�g�(k�O�ݺ�f�z~z����]�8�S0�LA��Q7�K�:�6�Q���w��nO5�6̀�n<~{M�y9#cݫTd�2
V	ĥd��bQh�4)���������|�$�~���r����њ�ִ�+\9���z�=>���\��S�s���duz�l4��+�͍,��Ō�Z~4���Y0���x��㶂����#>�}�&U�q�A+/�:����c��CTBбh��+́�(Y�q��QJ����+�O�<K�3_,rϬ}��nl4�!y�!)������V�Lҕ��|�#3�̤7zqMw��+@,���ꪬ��3+������OfUWcL��Ȉ������~�H�:O0�CF��A��X��x��V�%S�e��d�)��,=�A���"��XO����S�dN6Y8��ixf��q��fÖ[Gчp�
��s#�Ǧ���a���96R\Y:��oY�Chj�~6v��0>9�I���pyQ /��d��tD�`��K�Ve�q��]��E���;���n�����U�rQ��14����!rʉ��.��T�����N2���U8%j�1��dC�I!���'ԧ��<s��m�mZ�<#�m���|�B�S���rb^{���ߔ�uAr�(|����Z�]!�D���8k�C_z�oZ=+��[���O��em�5�����q�����=9,\m��ggn����?�/;�ꫣh2�K���ŗ^�.\���^x�o��\=��Io�ݿ�q��m�3>��9����|J6�'t�eɀ��Wh�G�:��G���|�뙛���*�{���]?�����Y�C�r��8W+l��hi��W�x�>�y@�P�^�-�Y����w�9~�_}o���o���ؔ]���'��`��_���Ɵȑ�T{�M;�|Y{��}��ַ�>������-�+��3�x��
֖_ �|���q��O���O�pU�z�K�{y�'�z�X\�|�3�0�Ǳe�d'Urb�|s�,oE��Hc�!�c�B��i��$�֋{r?�sw���_�k����q�����Ɉ�HH������]��V�K�?3�|����W_��=�;<�y��x�W�_����+�����4o�׷|����0�<����<Ϙ�%eN�*2�PR�6�>TE�I
�rH��X���t	�Ăq���ѥ��w^��u}���B����,�m-��<Q0U<ў���Y����}9	3z�>N��6��0���tt�QY��yѲ<�7�먙�'�0�@�*%ض+���q̺�k����Ӽm�<Ny���X���W�7W�+/?;���k�Goc�������8Y��?����,'�︒���qgG��e��MMJ1'���r��d-����W{>G|�����,�_1�̀���e��Z@.ʨ�Pm���~�[�"g�s�V��ǻ�C�ׯ�
���<��q(���T���c%GZ<�_��fmpBx~�!g�93��`d��<h+__ݐa��(c�I�b��X$���&ys+�ĳ`c� �:�ona$mG˛I��yཉsW3h2�88u8E�,�݋���J�<$��ld������s��'<r��o�A�Ph-&���M6vj�΂� ��%O��O|�o�����y66� �+,`�nB�dT:8��<|���^��㍸d@�d�no�:�C�j�6�0�#�:%ʙ<���c&"?��I�Q��F���4N~��C-;o�UD��8pzLzCc����ڰa����WE#�fy_'�C�m��x8�����1/{1e�5ϼ o\'߹˕'X,Y�M�V?Չ���0�����oO��%8o�\"�ZzA��?���ĉo��q�-]Q��q�x������ʦlk��P�?�|�.�j6�`WN֝�n���w''K��oS��[��\q5�P���J^�`���	�)x���Bg�D#�8<X��۫,}t�T�Ҝ�	�c&=�c2M�b3����RXG�$�W�x�m�nb
Z\�-�@�}]���%�ǜ��%���!�⍙q��A�E6D���%��
�6N�uUeЊ�@籍�rk�o��-@J,����%�J�J��l1'ø���KX0�s��*g�H3Fl��9WïǈX�*c}�86�9�3��9�D�N�W���ģG�j'8o޹=��>k�+2��-Rd��gn��,W
p�\�3<~v�H��-1�}c�g����~������ݻw��{w�����/ə��|gjߎN�!p���o���Π#<�e��3gQ���?��9P���׻��t�3�q��^��!g�,��Av�g���=Ș�n��!�!�˪\r�'[a�z�q��\��`C�1a|�lަ'�q�A9+�5��qR���לaC�ȸpR[}6M��W̵���->���`���`��_��6c|��G�o��oǟ���w�0�������s�;˭�7�]/�pSNȵq������8H� 7��J2W��/�����/�A�1u�>rX�vӏ?�<q�x��f���g�R�{��W������'o�+�[��� �om�ۺ(]]�썏n����c�w�l=�>���I2^�$�r����Dr�4>|d�������k��8K���so[�ڇ㗿~_��a{�[Jk�̞h�H��43�y&K��s��)����O�Y�2?5�-�X�E�-��	�#���-B�|�?��ǀ��\�>d�+_�|��	��6�}0�l`�j������% s����\�X�5�������DD��b�K�tBd
�6�Ӱ\�����)$�T�z�4�},��/R�v�L�̚c�o;N.�`�x&�5���K�xy�v��aV[�=��1(rR�������x�kύ�����������_��e�������]�z��!�$'��Lp{�D��C^,���s�.�pr�9�N=X,W�0~(�
�kA�26��`��f1��ھ{W^ ߸ѦGD�}�Bƭ.�a�z���&���{�6Z�e�E|�b�͆�#����2t�u	Iܽ��7�Ψ��U��1U�L86��]���M����-
9O�l�9�;��A�������Y
?Oa���r�2��T`$���4�,���@�m�քae���bx�k�u��0��R ����؛)����ʭQDգ��������f� x�_̫d�F�#�����ݫg	1J&#9��p����A?����SX���x��V���6}H��r|o���3n��o��h�gBorR�I#��_;YW��"�٧���U�!��۷;�W������ly>�M��d-�9�d��j�7�HJy[振6"�1a0:�<���x!$�qKL��(ZN)cl��1�"?�]��I;Y1*��2�訆���o6h�)W�|�:�Ng��vGtK;ތu �j�����
���يl6#��a��՝۟���z�AR��z�;�d#v��-�{�����/��k%r�y�.�qD݋��d�'t�M���R����`�iS�t��8��fi���$%ܲ��[���8�l��͓�����1���O`�o��G/�S�r `ː%��?��1�Y9v�1�^tD'z�:6�<�6O�=�/��rP���4�S�MP���,�����3Z��1��g��:⇰ݿ�	�>�������=*;I9j8��'�)�s��ܡa�"OFש�j�\�>�F{�s��ڠ�)�9vcS�l�}�ƠǄ�c�2!ߐsƳU� ~�>'%�[���e��q���b���ig[4��//��^^�8����op��Ø��<�6��'j��f]f֛/�'@7����/���5��W�>��];q�s ��uz��2H�$��M>�̳zr�5����dbڲ�Z��C���c��/����Ǹ��H�c�A����1gZ�:N�p��Y�wĭȲ�W�l��_xf����h���3���7�K/�T����������t��?����y������rx���ǵK㦜���>^}�%9]ύ�����~p"�g.��w�'}4lo��W�xc����Gr�x*�%�,n�e� �<_y��U_�j��+��V��W_�Q�_�H�އ���'�]����v�Y9�����n���������pg��fƣ������W��؈�������y��x�/�o���W��GG�"p_N��}2~%'�W|8>��=�����g�y��Ԃ��I#�Y��oZ���X�\�8`����j��1dl+�=52��$��`<C�p����wN8��c/2��SIcG��`K|zN࡝��u�$����Z���˂���~I`B��q�l��\`�S��Ά.3�⯩gl36���O�4)�����������41_�0����j/A��g�ȝ��X�=�1K�r��]�����x���o��⸼r�+Yv���g�������8Y��$<le�p>�w���������pr�'�+Y�)���F���-J��J�Í��jóX�t�E��9o�+�S٨q5�"gʹ���h�sVeG8֢�c�1�����l��|s�L��|x��/]�a�%�n�EW�m��s�8miqBt�����y��3x��%��p�'?
��c��(X����1� D�͆���㿩&g�y^6����js�[�(Sc��
l��P~u�q+��E�_����y�4�~��8Ŏ(�t����%�ci�S#�;�
����'u�G�ha85�q�pZ5.�Iu�-8H�B�w�'����S�1����SXY�Og̓�$RI'��Q��`�zcǜp7U=�F��͙҄}6Z��'�㶔v�$�W�q�y�M.r��B ��^?i�e`��{6�	񊌈����<��J��[��=�\I %��-�2%u����y�Q��0h�_z �l�9'K��T9X�>�q���7��]��X�y(9�&��1'y#�%�r����� pf�vi���������{c�o�̎/���6lR٠�!����0:�@�@������K�郝cE��fy�0����@[���E��M�������r�)��c��`#E����pK8�ɧ�>���n�2�-�lrDD3Ϥ����I`��N:"�ܼD��ӤJ���MNz���a��<��dN`�c��pƞ�d1�#�dq�ou��QD��	�y���s��p+Yqe&t4����w�]���n����i�M��oMe�.=��i&;�m
/�~���|���F��Y?��Q����Z\�?�T���5B�'�Þ�!��W����́T'ݕcJt�����>
�b¤���(�"x�I�JN#�!'>γ7v�Ԃ�l��vBmx�>'
Z�bC�D��Bg}�o�i��8 �����G��p��2��?t�7��799��5��� k� '��,�`;f;�����9�W�$='��w������;����x�ŋ�]�{c���?��O�t�����8�V��3%'�/���[�Ǹ��j��o�6~�������/��.�����?xߟ��-��q��0��4�n}�����!N�_�7ރIf\�ř��w�^�(���+r�؇���_����v�.l]�x�[��W��}���������o������ϳ�xY2�J���3�s�9ߐ}����7����uQ�63�}g�h|��m;Y?��I9ye�����4��$��A��Q���<����SA]��?Et��<�b��L��tX���hJ�����yjp��Q��:D;xm�3�(�>���	�V�����|�@�h������D�L&������"g�>DN�����Ewi[E���IJ�ؓ)p�(:G嶛B�ڍ��.;n�g|q��)�r����e�,prrpr�TȘ�ɺ�1�x��������ʋ���va���.8w���HYV��xC�Ncԟ�d��g�Pd���R�6VT�������W�l&����5~6c(1_gXe�mT�wyu}����,���?)/'���EE�Pɑ�1�&�#z(�{��z�rmGI�����9�/��/�}�	��W�AaÆ��I`aBD�뇵}�[��u�P(��3J���'<�����B%��l�h�F\(��?�-Š�7�|W�����[�sL�B�,��c-�8Ɓ�'/�dQU���h�?-��]�:�tu��J<[�Ǝ�U����x>	.�jX�w[Qb'�^����h����2�۸�K�I��!L�Y�þ��<����g,8�
dE�A4�(di��"o�L�d��K��dƆ��n4~]�1�X�����q�J��/��I���5�L�#����4�-x���T�`~(�#Ԙ���W���^�+��(��։�r�d�v*��u8��k�c�<D���f�o��1�l$��3śÐ��"�R�6�߿3��|l߻=>�sk<ؾ-���o
�D?�?%3F��T��=�?�I9�φ[���H[o��s��l���A��)>�����t���f9:����܃��|Sۖ�
�lB	������w�1�{��W����v�^����♑w�3���uA�\:N��`S/�/�\Ǌٌ�/�W/ؠ�yD��+��+'��'t\����gɉ�N�-}oۙW���ņ��%�n���C�ܯ�x6��_�$�	�|;��x�c��E��:�Z�ӱ�3��+�c��8Y�8��8YP��	�TS������3Z�8�s6���u��C�q����:n�S�-�^���~�M�ñAVq��N��׸��!F�~Δy_��ZH���MA��Z��\2��6�J�^��]먢�!���Ȇy�k��	:��S`�͜,�窚�_8�?Ą��$Ƃ9Ɖ��w�ď$\�~i��G������o}{|�+�ޜˇ����������?���7��sl?�WvoI�sz���d\��>���K�������v�._��>,����ƻ�xw��?�>��'�x�)r�#r�y*ߜ"�7A��Ň�y��?�f"G����VD^�j�#�_�_�b���W�\���5���ۚ㽏n�������w���w�`-i�%����R��C1~�P*}��5��[㕯�4��η�[���(��@����[�����{�r�>��ָ'�|�1[o�Z/9x��dѸ2����"���Q?�)Tv��)�ƙ��i�!̓��\���u�����s��E���I9�y -ژ	��|r��s&L�UFI�Yx��}���I�6���o�Z����3�É]�Y�y�>�l8&�;$�a�|��?wj�{�r�T�*�/��R���{h�ƕg[y���S����Wޱ�q���Ut���.]?��/o��zi��{r�������؍��_�d���������]	teKNo�3ڲ���vAM��7lx� /�8��4����i��X)h�N���,������HZ�eyEv�7�  ���
ޔ�֑6b|/�C�Ω{��������
.�ŗ��(Rv��o���-q%�'��8�ϕ6�Ŕ���<�d���(v�4��g�a� ��ԉ����B�B�EM�I(��J����ucR��R=Ox���+6ꋯ� 'N�B3�������3/�1Dp�d�o���J���M9�v�b�˽�.�?�g>h�H(~�~i�4�?�>~/��.mI��V��h�^��:����v]A~q���G�7~�N�&lo�hg�%�g�|��a�BW�	�U�l��ϲ����T֤�-����%z�h�W�2���9	�N�o��.��e��ڦ��y>Uqu�<�z�C������Ju�O{M�9��j%�Eʘ���Q����cm���dqK��qж6�o4�����,W�_�;:�~:n�d�w?�T�gr�������'�W��a$`,�o���r"�8�O��
��U�3f�e���"`�*���uL�m���~)R��l�UI��.��I���{�a��9C;T��v/��x<)סK�'���Yo~���1tXp�߾� ���<�-|��� <�b��[hF}���7��v�	����=v.�C�e�M_s�&��t!c�s�@h�~M�7(��\l`ih�����j�8���������^���t�\=�4%pD'���cNrHz�A��%<rb�s�֒'6Ѭ
90_�ܲdA[� n��؈O-|7>��_�=�؀��26���$;��"���=��N/�2�MW���uO1���F�Ð�l�rN/��X�D��3��D��ʐ�/�����gҌ�"��!i{U��<'^���|���}N������
�7 &�����xê�Oȟ���f���C���/���;ߓC�[���}k��կ�����;Y��/�b������ǲ��_�μ��8>ܕ��}K�w�����?���_����{V�7�L�;���'~�+^�K6���M���}g����m?�����(�����l]��<�������+^���M�ʶ{)]��C�<�������?����K�֝�����Wr�>������q�{M�a]����a���z�~.���_{�����;���w�d��� ;�Oo������ͭO�]^⥹��/�ʢ�@�m�����{���%0o�?����L���Y@�a�9�<���*+4�:��ʃ�o��E�RҴ&�+� '�h�?�s�O��~��GJCF�J�6T�s���h�?��,�,��7�ӌ~پ:NfA�eq�ɪ��#�8�����"0�F�3L��|2/{�Oc��lx�B�Ʊ�O.��Vq{3W~�a�x��t�����g�,P�fY�Z�C�rU�����k\�z�W�����r�v4{�d�?��?�����}0~����d���a��MM�˗0\8Y4������~o���J{]�����/,p'՞��X�(�0��j;J��l�d��9�r�#�f��*_��=����8X<���P@�+WVJm\y�ƪ���B���X���z�� g���� !�3O6h�#��O���KHz"ΐr����R��� ؄��"�r�'jI͙M)�F�E��\�Kɣ7ɾ$za%��,q�2��Nn��F"�&�麪��Qw6 ��
27:�����e	�	~ƚF�����b3 n�K9m5� #p1��Q��y���$}U�|?hE��hƹ7^�S�6���l��?!#τ���c�N�"*�s�=�,�v2�O6 |6�g�S��o�n�}��Xf�A�`���o�O��Qz�f@��g޸ʶ�<8���"d���%n��������@�1z��"u�5n��K68Y��ŝ�q"+XQk"�E�[9�bp�8�ĭ$\�~d�3)8p�6�q�℧�#9Yw�΃<�u���q_�֎�,��!W�oW�a�~H�70�L��K���9�	���t�z.�_e;p(�ˀ�̇ ��\�})'S����Y��U�>�g<������;���,vz���7�O:+\�_'$��r�8g�G�Fv�/��`�>�)WUT�P����#;x�;d<=W�ek'�P釪��}3O:F;	�_����� 1}&�?RxA� ���q�88��ͷp�����$�a��g�
�e��]?�X���Y�ʹ���鏝c<���'�j?�%}
o�/s��g�8a�1�ȉM������F2�|m�9�Q��O��#�jLX�q2�'��m��[j��C27��ȇ��rg̠�[����g�Va�����<�Ov��<��&���Vzp�S�X�.�|��5��n�u��M���+�q��ߓ��I�N�N?�y�S�ȱ��,�8�rQռ�y�[OZ�ON�p�A��Z�{�;��[�o�=^�Y�]y8~��_���˿.G�'rP66�]3�ғ�=�.���>������5���`\�|Y�[��;��x�!�_���r�x���l���'\�����w��G>�Ҳ���kr�.��Ꮚ�qE�c�/�f�_:��{�����������;?��q�򸳭��������c^!/{|��,oH��7�K����h)yoɾ���K������=9Y[�7/T9v�'�ޑ���x���'wn�{8��U?�Bcb�3p/�[��4��`����E~�<9�o8���2�� �)[9R�����Sp�-�H>l����Se�_�M���DhC����i�s��� �����+9R��@k��[�w�C�/��b�&X��B0�e��&A>X�8P8��!�sX�=�(Z6r��Vt�'�;Ȓ+��^�t�
&�=�����&���Õ�V�o'K�+E��%\'���ﵓ�+����������l��O>��h{����l��g�$W�r�Υ-m��H��8����n��%|Cm�$�G��U����J���A&�12�N0�dZyX�Q�R\�-�x���Pm9�N�l X��A���� ��/�������#�6�����Qx򼘂�l6��`�l����J���?�B�ء�@;G�٘) C�Y�#�>m���ތ�G���d��"/X���X�	�)旳46��6�*̲���8���LưC�`�%����gI����iA}3�E��P2m��W�:T,`|f����9��e*Y���}�hH�|˗`��e�IZN���z�UI���an�Ks�MgVu�> ����8�/�*h/��l=hyL�@3�]�&)����#������r*����`��r��6�,%���x�\�����Hs��Ù�C�=n���n���p|��>F.ȍ�R7y�\_�s?���cW�l��}?��g�Ti�c#��sG��D����4]7��]���Ϻ�<��1��w�l���t��9�0m��+4�Y�u��-�2%3�� �`g�L�+!�}x9��2l�T m���)��ɱ���crp;�OUe�ӏ�&W���~̓Ɔ����|o,u�12�B3��]���zuVn�`:J��|J
E7�������`�H�?`�)�3��]�	O�L�}���s�?�蟥P��BLS �˙S懐�િ���e���)q�q�����@��:dtĸ]����=���c�+�E�#� �q��$�o��ķ�J*�8o���8Ҝg�m������++���|c����������x�����~������������?���h���Er�*o8����㙛W�w����G����_����D���θu���ӟ��W��������d��W��������J�iO���t��e�,ۆs��|�oi!N�ᄢS8e��mpRA�}����[��;��3N�6ǭ;�����}pk�����g�팇�Z�i�mIv<>"������>�Aqkce|���o	�o���ȋ��[|�������?����q��Eyk���'_�.�0�+���G��ҭa�\/��h�ט�L �_(�0��pa�(��ƆFfN�Ǯ��X���{����Ӽ��{"
N`�=CL���[�>�tgC�w�4p����2!k���ԟ4ʘ8��r�)���Pi�����o{�{�_���)Pƕr4��i�mr�i<xfS��ѱ]�@����x)o�d�����f�������I��r��b� �0����\�0��ڋ���~m������<��~�eF��?��ON���,'�C�,�Y�8�N�(	�7q�͇p/mic�F��<d~WN�CM�]3��z�0q8���MB����	e3��A
�W�W#�[�Jpث.����,�ތ
�y�@ra�%��4/����!��<q5�<Af�b#��*ܫ͞:ȶ�m5d&|��\!�[	{�>��F̔c,�<	_��eR�L|L��vF}��=Q��d"x���i�4�#�g9J�E�1����"=)4!~IH�l��d@(�Z���C�h�B_-�4ɕ�sȞ��?�	����U&`EI���%�+\���c�i��Xz�8ۑRD�"��Be�S3��0�\rƨ�ACw��J6<;Z@XNL���<t�c;�p����!ݗi�F��R�F H͑4Y���g���F�ls� W��[�����8��b>��Ƃ�v���#��pL�S�^��}�c�r��#g�WT�l��6���3w����4�m��.�(mT��1R��g�ěKdCȇ��'e��RC�v�(���(g���q�)��������7�o�����ס�G�Pg;�@9:%���qE�K��rl]�� ��N|�׿9�Ʃ �L�Ƨ:�N��z��7,s���[\�5WG����Y�E�6����m螙3����s.m�l-������!��
�V�#�:s6�?N��P0�
�v:�N)NS��DhdO�g+,��Sd�r����6W�p��p)� �jh�K'[r�֘�F�"�-���8�ǎ������{����ƛ_�z���x������Q��ߏ�������}�!'Z�9�,2�����;�ys�ɟ�������'��ŋcI{��w?�x��?�q�����Gչ괷�]|Rf�N��#Z/���gIp���{w?�?�5>�{�N�o[W?{��/�9��.���/�4~��p����흃��{����O>�'��ָ}{o�x<����"W����\}eZ���������+_o�{����`����(����������*?Җ���7~�P�FR���Fc!�MJ=�)����*c��B��C�+���V$�b�Z3C�jO��)̮��#R6����[��!�8�ޗ�b��
��1t���@?G�3�A�^�������,,x��xc�8vR�B2nK̥E�j}E��Z�4��rP�FG^ɔg�RJB�>�	 %�,��V;^�G!�.��M��,���P����SQ~.Vٻ�X�&{�̩���*��.z�����׿����7�d}�u_պ��4�����w���O�[��{4��gXZY�^�_3�憷q3�6>ǚ,\v�
���N�|��?���ܕ��30�\�BAc�3uv^A��d�f��V�N ��g(t��?(�FT���_ymk}K����k��?�h����=��꿎y��PA�
}6�J�m�D�v$]�-�ܺ���<Q��C0�?�6���ӆ���y�W[�"C8�-��?}$b@�Wm����w�j�XS�sh]�ܰ�i��7��O�:~jdA}G�WYG����Jg���R&#�M"yމ���N���7>̇t�S"�jJ�v�c͑#-�G�㫔��yݮ뎎���9^^H�����x�b��r����W=��G;�¯xLzH^t�?�c>��<�j�+�j��\uJ�r�=�y; W����9�}��]�݇۾m��|>���x�}wܿ�� ��)����{>�}p���w��P$=��;�iR��F��~��}�]m&8��Y\�L�Y(6_���$M-z(��<V.sL�"Rc�0�5����s���1�Pi���ܹv)�����98��p��t�r�E�E42��/'-�u���u^9�Tm	UN����ǘ��ei�:R�R6�F��3���l�F�rh%g[�R�
'�r���#���N�i���)-7�z�&�_�a�ݤd���k��iW�S����Ut>NDʂϼ�D�-����;����*'D�:��B�c�b��3I�0?~rtS�TL1|�e�>Ǧ�އڤ�\]�)��c�B.i�=��w�N���7��׿��x�����^�:67Y�W�ݻ�ǭ[��'�|:>� +@Կ���Ƞ�n��8�u�����k��W�:^{�U�	�e��~���~��9���eOwl?y�*χk`>��(��Q|���G���g�*�]扷�m�+W�������o�g^xa�����n�˩�����/���@g�������c��?��x����s�<+�rݷb�/�?�\x�*v{<�]��#䶢�%�Q���XR�ž��WI�v���Č��.w��GT"8u<���{J*8��u�� ����'����zUO��}Q���Ix)�<��/�����0x`%��
m��hX��2N�T��C��E��||H��U^Y���,;����Ѡ�8���)��3�a�E�/3��Cn�>��ۉ��T[��?�R�7DÏ��������l�s�\7��C��z��������[����~p��%B��I�R)����5q��|b�4���Yx֑K������-�͸���ۑ���Nc
	x��V��+�M�,;f��߯(F �H;2~e��&2�ja�G�|+��
�p��Dg����P�(�����gM�����^��Ue�p����[��z��z^X����������L�W�pQ�H+2�2(�:*P_��٥mצ<Η┊Y�8.O�(��*5z�����q	�-i�,��]�p���m�)x����I�d��!��j#��ʪ<|H�����E�Ѱ'��㊜�t:9cj�0q�䡨X��R�S�(-�K�U�2�si�4E��o���Iy#�p8�B�s�Qh���%mF�Sћ�w��p��U.�L�#9]8h8_�y;b���sV�YI�#m6p�p���ړ��w��v������p�t�C�3u��~d��g}��?�p�ә<�-�VC���X����`/�ͪ�����;(O���:��_�l� s�"��ؼ�ӛx�JS�q�a+
�y՟ȅh�.��J9)����W�y�3�����"�:�]�;�P��S�Bo�d�H˟qW�:��V�V�:&Bc~�2�
��˨+\���{o��k���4�:�ł�����c�\��s�����`vꓒ��HI?Ƃ[�Yo���(A
��*���׆5<����,�W�aҮ/�3��U\�W��~~L;�:?����y�_�.c _ȴp�f]�#�
�ٕ܀�@|ś+Y8e���W�eS�y��x�o�����x��KڿȬ��ݻ� ��-�~���@x�G7_�����W�y���������۟�[~0>��C���}��ʕxnu���q���.���l�)}7 g�y`�o{l?#���:$��uq\�vc<��K�7�16.]�~~o|����}��g�����ng�,�������@9Y��@�7o��k�9���\�s�����l��Wɛ�Z�� �7�^� �������֡�1�ʐ΢�~~l�P�ˢa�MC��ׄ*���뢏�ӟ`��ʒדb;Y�	�cXc����ĩ��$�']̝��x����+McO��%�n?�)���'%��"��6��s6s�<9O��}������/�����_��}}���D¶�ƴmk9�M��rqK���x���㺜��u�i����r�>�����d1��neM�,IwD����r|%�����ɽ��@�Z�l�c�I168h�}�׍��x�.Q��Ò��$�Ac�Ž���^[��F���@�4���Pq�
��g]�b��sJ�jG���D.�Ҟ�A�Q��8@b�gbxU� �޼�6�⏾l^زc���TW�C^DW��'�&�,�3�1��=���>h��/"y>R|Q�pSm�)r�]q~��`'�9�$i����)�$�#Iô�`U�YI^4P����hG��8WU_Qrp�w�#t*�m��F��a'e����s��0��2E;rn�\��wE����vғ��0�K
N���<+|�F�E����:�-<�E����rťB���i�C-�+��X�<p.xݶ�p���U��8��&��ǲ�;;G��Q�Ô�w�2ƕ;_ɣ�+l�㘶�~�b��K�Z��fR�c6rl�Pk�R�lf\�-����}#s� χɠ�B���M\��$a:e��q���X�t,��&:�~:&?�i�?��ʫ]b��6��<��t��<�a�X����eѷ^�b�NJG�c>Ň�o6ݧ��ߔ�C����>dM`A�,2_��?�G߶�_e�/=��f�M}�m���.Wt��~�BW)�xp9�g�Qk��W��C�ځ,:��r�߷�?%�� c�|6�u\t��$t���"�Pj�*�`�[�;��Lmt0ј��-�ٱ����t�����_�<.p�Ob�Uu|ں*�b��N������&9��f�l�VY��h�2�K/�0���o�J֍��^��]9%�}zg|�ٝq[N�����:��ۦEwS���_x~�*'������|\����'r�x��%���]햳�����CE�wqG���T;|���G�I�Nu�g��~�%�1ٺtu\�~s\��̸��s�H�8W��a���{*��?��5���C�Kƭ}k��r�K��oYT�._��������fo��~�ݾ7>�����-��O��{^u��S���w��Y�&��8����8Eۏ�b�(�{�	qE�1X�
g�(5�_�>L�u�1�tG��H(�E?�8֢���h��i$I^)]��L�=���'�'� ?�_�S���j|��?3����ձWvW!��)�r�#���;�U,l��8�s�W��nb}F��dT�ޝ�U^�C���nz��
�uٖ�7��k8Y�ƍ�ߋg?��o�W��r��J�&���#F���>c�Ȱ���IRg�ŦvĀ`�0���=W_068M�P��^�8��ɧ^�i:������Ç�y�bO\F��ǯb���M����{��W;o9��J�3��M��&��
B���X!D��9N��W�r;#o-��S m�if�S;�g���3�A�����i�N$|`���c�<��d��=t���yj�F&<Ȇ��Oi�MY�P�N0��v���/������?â<�69�@�t�<�cDߌ�a�8������4��P���.�ב����d���Y$ox�3vb�B�4�v<
?u:�[����������Ù2�q@#�M�N�_�-�9��E�b^�|nkL;ә��OE����j��U��'��6J��j�c�N�#ǌwh���A����H7�ƥ?��#�J�9��W�H�9K����oKK��?����bx����[�1�".�̛7��fqZ88�杘�da+|ؕ���e)w4OIS�x{�&��`�qPzC�x�E�Mf�8M�;��j�����N��q�š�,�nu6��c���>�Z�(�᳣6�s"�u�W�"R���۹r�ĕUmX96o�ڤM�(q���q�����7^�cZ�������Y��7m�W_�}�.������8;^�
�/�q�\w&��>��N��zx��Y��C��V�GܮF*�:f<�w�+������ [r�^o���񕯾4.]ٴ�r�����\m��w���ܦ�ǒ1������즜��{^����������y��w�]>�,���/'k�P�k?{�-�������켍O�9]XCNC�@4�����t��˾Z��qA{"N4k/��	�+���+7���kc��%���@���DW[�����p�d<��̀�!�O����U,��~���k�<g�ɭ��/]���A��<˫�?�W�����=S������cBTl^c'm�L��R�Me��R��_Ŵ@cg�m�4V��K(3��ʪܑPy��_x�����|lb��i�<t��`��i,��W.E�+<&G?c���_�����~#�.�Z�uZ���0<a��|!{pʒ�<'%S�v������7)e�%��?�{��.NN��o�C���yA�p�S�Y����u%�g���r�.��?N������>�#'���~��]p��Q�:�#d0�7$�$s�W.�l�����ߊF
#�v�xX]���r6>��NWH�<�����U�8=��j�\'�����=g�1�j��I�T�3$v�����I8DM
�v�d�<^�A#�zd�����w�2I��A���dÈs��ӜY�,�y�Gں�y�	���;��1�V�ř��ZG{hE�E;��d�7���)C�͟Zgq�������u�ꗲy��bh��<���vS��M'���S�&������-��י�8n���U]����5���8Z���L����"8��<�GxH�'P5�%͂q����/�w�m'�<���رyZ�8�9����q{�S�y1}H?�"ƹ�_q�&ٸL��I�Q�Ҷt�b�XtՆ��З��z�b�u$L�;x��#�:�n��B��l���|�?��|�P~���b���p���w���5h��7�[D�*�y|ڹN�q�jQ��/�E<�Z�%16f��0�rljl/6.rQգ:�����r9 �tڐ�q%�"���(���y�Y�u�mn�u3J��7�0`�<|��WڃG0�3���Y�'���0���Ь��IQ6?Nì�"Kt����,2,�9_�N��A������	�)��Y]>+3��:��|���In_iO�l:ڹT
��.��}�K�8c��Ǖ!�yI{��M�k��!����=��9.ƫ�~m���k�矗ӳ�7�����?�}zo|�����;�kM?G�rL�Q��I�6T�F���t��Ҹ���q���q��{c��?q{Ҳ��#�4Y�ѥ�7��+�(m��i��7�]ϫ�ƺ�����H~}�#߾��±��>�����cCp+j$Cʕ+m�#>�s�:�w�ƃ����}^�~��oH�'�l��8Y��l!��\��u��u�&h��pogܻ_�j�ƞ����n�܇���ۉɸz�!��)uެ+%�f��x��3�0J��D_Ф=y�A{N���ʈ�#����p.�>(q��S��R� �m�'�O������F`�����_�s������w[�5m�M?��BdI42���'U��s6꿒�;��u��ylVթ��:%�o^��8�r����i��:N��r�$��d���.{N ��.�+�.�gn^/<w}<{Csm���d�/�w��%�q_���O���q��Ir�Ea��A6K<3��q��� $����,P4�L���+RJq��>�1��2�\����զ8>83\��w;�����١_�$�f��o-;���@=����3�<�o�r=�iq�Ou��b
���k[iý��XX�a��^\Tt4���W�^��:AC������nޔr&�Es��)�]��2���������@B�|����W�/z]�Y���e���a��5�Sc��q��?D�S(�8S�����_�9ж�e�l�V������ܩ&�<rΦ@��KE���?�/AS�jчÂוU׿�8�꼉����F��󳲂K[A���$�
�M�>6&Ĕ6J�����_�r����qsLQ0}ˈ�-Ʌ�\��ڻ	��&ѷM�����,��-�>It.�2��_�����t0�:��#Q��G�/�K3�/��:P�)p�e>!���l
NL�%�=/:�,Y8�|��\�ˍX`s�3'%Ԋq��-h�aR	�f�H*�\�Ne���1�wƈ�㠔@}`:�ʢ/�~S��Ѿں̠3y�@�'�AU	%7B�q"�h�s��~a�Ya�qLQ㥌���:�n� �7"U��8��)2�3e���}\���x��Y���DQV�ٶO�otʹ�-��� ���o��s?z�z&�6�krX�V�da����3M+��ߦvJ/���xᅯ��7n�x�o <�^�����>����g�V@ru��v���.��[�4���r��ޕ�u�פsg��D'<����)8Q[������E�6�OZ��sx�>��Z^�k�Ɩ�7`�P��_���h�N��_�|]N��q��u�]k���;��(|'C�:^�Ӈ�ŕ�ñϛ�%�%�n*#b)j^�v���/ظ~���)��yϴs� ����F{�Yh'�͟��/�� ��l]R�2�O��Xp�S�ǉ�G���"'!H'{	>yh�K�Ug>9.��7��_R���h��#�6[O���~Lx*��;��/��!m�c5M��*��rSp��Om;��;�|ɬ��|ް�|"�����t���=b����e�7�>����N��]�'wV�f�_��d����^�) n�iN�q���+���\/>��o��i�7�7�d}��9YG�h����iC1D:��n�)<O�_�A�Y	�q���8�!f�q;x���4�`q[�#��"�.��\�C��>��
u|��x%��
��8+�!×3�Y�p �Pd��ߩ�����-�8�^E�B�&����[(���ge �@[��
<J�ӖM�� �>s�14q��Ně�ƕ�\Ii>z�q[D�ڻ�qx*&J���	����҃�oj��q���:(#�2�ɉ	L"ʻ�x8���bp�C��q�Ć� у��9��z�9N�S�E�"�L����,Iո�'���-=ݦ�<f�L'1�h�f�����f }�c�}<4��hByڠgԇ:�{��ϱu�ʽ��9��'�"?�g� O���ɃG��vD�s������x]U���Ŭ�-i>�8Ƭ���i�<��c��)��!Y�x�M��V>�]����[�?�+�X�~�x_�㟶?v6i�e)벘K�缃` T�S�rJ|�a�?��EYs"���,T��[zzb�m�o��Ġǰ�:�\�Bꊮ�+�̙c��ү�q{EW�4�Mj8�"熤=y�V��U��0I�aB��*p�j��g�v�|Cy��0��@;/Z�@�\R��"yW��DA�|PTQ�&	W	�T7��3Ǆ\i~<L=�]�x�h����=��uSze����+(��|s �TQ��y�w���.�K���"�����k󒜫��g��}�fMľ�"�r��޿�����-?��w�����\�V`l��9X��n�Ϲ��}<x���F�^��w��*U9TK�|xE��1��OƮ���;��]����Y<7/���-<�6��]�Q��@���Nߦ�[���틧}h�1��X{'~d��L������d��� �,$��y��3r���y��0$0�w������d�8���8nZ,h�MÁ�1NN\����E�܆�0c?�&��<��D�@�`�����z�S�0��I䘺�:�8��=�����"p�M�r��,_ǿY���yjˠV�z�o�IS߲v^�����5ߦ����٫��L兿�z��8}>��&�4/\��8]M+�n�����k�/��E�G:f��M����W=Z �&)/��~��x��n�go^Q�q2V����+'������x���v9Y||N���_��Aӂ��y�6�~1�����#�i�͋��*�"�D�?B@������b�8;���Q�.6ikt&���7$��Țr�v<,�+Q��kV�sx�ӓ�^jl���Ɨ�팁�ʨ���sū��@��"�J0fM}��:ޔ��f��V}hq�2D��J4����&�yE�`ӸTR
/S�R�Q�nꬤn.V}GÀT�ɸ��)�T0v���?����HV� O����ܖq->������˺/a;��Y���tbߚ�f� �
��c��gB�(��T��D���.7�����eg���,?�i������U.2������h��:P\s�?�dD��G�t�S�@j�h��� ih�`�E["�x�6�J��7����	��ױ��O��[����k�%�����r��1I9�V�)g�8�/2��d��"4���<���͘P���9�	�*��,lw��嬷FHc}�$'�:����g�M�J�7��1�z��o�:N�Y豢�6�"5)`��2va#0��J|�<�%d�O���o���n�L��S~�+2����~�~N|9���@�ᄁT2�����\�&���S�^�Ge���$@I�i�/���A�bo��+?;���TC�+X8X,����!��A�c��YVm�����q�*�?��m]��:�U�%9Y���r����,��8��ǘ���݇{c�������m>�.'K��������}�Ev�U�7�������rXv��.�*�xB9f|�W^�ڎ�rL�9e�l�绸:F�/:8O;{8Q���Pq��!�:��E�g���s����X2C%V�L<���5IJ����֖�Лr�nz��>���p����{�s$1/$�����!{B�*��g��NSI�u��D�;���c#ud]�����A��9.P�iꦴ�IÓ���h�w�Q�\Ĵ�E~g����]NY
���e���Ƞ��8y�U]S���SG:�a>&5nD���	�������pMx:Vy�J{E�W�����Wo��<~��Č�۾p%����U{����d�a��|���r���:.�i���,����O����t�����Ƿw���8Y�'�W4)�,B"��-�,t�o�����+G�&�$�2���"���a�4Õ.om��W�	c'�q�\�����l	�GF��;G�1ΐ��Z����o������ܴ3�t�H�,�G�Rʨ��"�����/��[ҟ:&�J ah�2�2+0c���v����M<�2L6+�8߄j��7$r�#����P��b�
.3.Q(�%��"�� J�R����]�����Gd��J-o��O�V�c5�\X��Nїt��(X�yd
�&���]�0��s܆2u���gA�N�4)xʴ! h�M!gk�@���d�S��p����4��`���w�w8�����q�"t܍e{�ܭ9NY��A�_��vq��mV
݇%�3�컩N��O�#����|�@���ei�<s� �SP�ǝ*�Ê��4�*���,j�:&��9?T�J�,`��1m��ץ��/�_�d�_w����Y�$�GY��*w3`ט��ukj]�����y�\�v�<�.P���x֧d2�?vz�AM��z�q^>.��av�Y�]��0����2���ՕR涴R���FP�Sp5PT��N��%���g��|�	�!kCZ�^���D��+M&|�a�o����`{5�%yb@﻾q}p{S>/���^��s�<;�xt|0���u�Ɍ���x�m�D!Ĭ����=�c/�/9�����\o������x�o��_z��`_Nʻ?������{��g��+9@�����ߨ��e���I�>}��T�8��O+޴f������رgI��ƈ��#�T�{�:F�,e��h�9�99r,U�]�p��cOsuWΑ�EH���}ߺ_H��GR��.n��.�����͛�7�o~�[���~��@x�<�}����~���?x����timS�-�0�M��я��ny=0������gC䒚\Rd��NC[�c��¥\�dNJyo��"m-��$���R�C�|�Y��.s9U�r;�KY�,�j�:l�*�|��� _��Z.����WiX��ǎ��/���`�������*ؖ�,��4�pP@��JC��$�� Sxt��S������Q�x9�v��	�04�WD4�W�kz��`\�G���ώ�������_��������XU�ʿ�w����Ƿ����p�D� $�V�$ZM~�Mw�X䪍2rX�&s&��H���,[q���,Q0��|)$1�ШY S��a՞��(���
]^9� ����=l%u�R�(y  5t���� 댂�-��ƫ@�?>R�φ�n��+z�K����W������p�5q'�d`b`�lG"�2��F�\�AV�`n~8����v�:/��10��s(;���L��c�{Z�CM�Q4Uny���͋�������y\L��w޴�y[D�Fp�>�mH#�E_R>ɴe_JZn��'OG�}�o&G�sOe.�6�g~�l����A�se�{Ӗ�fE/�B�1�/�#��'}e�/I)3��N�zn�_U �Q�W~
��s1� '���[�C��n+xEڧ����δ	3�+v�|�5�.VX�#6� ��d�~�SJ6i�_}>Ï �~(�]�%1�nK��7��筮������t�:�g�F�~^ޱ�����F�
՟��`f�Rn���4�ɘ&��+ɧ<2��Tb�u�6��^�_�g��7tE�	�Y��.��n�X�l�R�d�w�g�N�k���[4+����S`������8��^y���30�S*�~�����Z_\_崩c��r%*��e��N)�L3|dC����3C���X]W��nl��_zn���W�׾�Ҹ~���<���f��������g�����nmx}���|��z��ߖ��2�	�9�X�3 {�~*'+k|[��]�s��U?�=�3.���tx�cXK�&��G���y�0�.�qL{�+��?0^�K��Kg����0.*^�xi\ں8����(���`� Y\�ta<������ύu���%]�ap�޽���k���I^�!��!��i[��k	��L���(��>j�E�T��kY��<%P���|�!X�M��GƂu���i ����M8��:�*&�u���R�Y�'���6�
�+�+�:g���o���L�U[���С�k��\���94��o:W^�&ڳ�.;�_��t�:��>���}��c+��=��.����V˸t����ѿ�a�9� ��7$o����W/���6�����̍+c��CK������O��'�'��l|t{<<�S[�p��.�d=�� �P��K�|�x���GJ��%�T"��3g�UM<΀JY8����3�Rh9��7�	�׬f"`%�C}�M5�c�����\]��C>��vn)��r���%
��HВ��Ư~!�� J��_��y]5g�08(�ԛ��^/"ŷ�1��?��9�E0����S��x�Q0>��M�~.�mO ��P�5ȗ�[�/���$�Wa����U��>�s�tfe�|IV�>��Lْ��I���tN5� S����r����W���KNK@
g�)��nG:����ժa�#D��}���	�v�VY�Tm'�Nܼx�?;�.���՟���~t�L�u@���ӊ�)
���&����V[_�(�&|���l�XJ��'�y�	�I��ւO������������W0c��%���ᰒ����VO��</���Ο���@x�7/n������e��4���w� t��%�ll� �y ��y�	<����[[���y�}����C�YxIJ8ߖ@=�z}�1v����=��v8՛|cH�&�n�9��Ō�4na����������8��wl8V��,�S8?^��́R�E��hH#�hZg���w_����+�Ú��9i	&ڠo�v\���$���Y¾P,�T׏���d��w����W/�w~����?���w�;��q�]���O��������x�������������B�9j�r>�������/���v���LV�~�4�ֱn�풜��/���Ȃoimo�w����xr�����2���-G䆃���ф��Mˉ�Jw��l?ؑ�v�� XN�l�Y�#G���5�r�x�aw�����HV�����x����կ}m�����¥���8�l��~4~����O>��d=Z���,�0x,��)�E��q��>=����A�r��jۤ��z�,*T�?�u�n�0��zk�JȤ��� ��/~&L�'�� �&���ڠH��G2���5�N:�Ƅ��ph��� ���2	��a�y��g:�ӯQ��qҴ;�ȟ��Ep��ߢ��m}�1u��0�,)�zd��5�D����ӕ�Ib�v�+�k��[�P����q�����W���֫��}}|�ǵ�G������O�ǿ������;{r��tYN��OΖ��j���揎ʉ��r�gCe�����k��`9�N�ϊ�VA& f��z���%��c��K��r�Q 󒆔��E�B'h^1�����ЄFxAb;g����d`3��y��h~Ń���	F���D�)�rW��ړK�����?�B��W�J��S���b������T�z�3=6�0�$�DBpѧ:�4����ݜH;�����64����8���x�<?�s	���`a���)'��b�~U�S�8sL�����I����O����j�q��鋿�5)1�i��u>h*�e���&���x�b4����7�dq����"$��su	�ש�r;�7�O
FR�H��Kvq���XҒ?�F�{�	+�h�o��w"4��Z��8h�L�g�g�8�;t~ކ�m9J��Xp���'�.��00����꧅�je�flR�fA6x��q���	{ز���oل�!6�wT�y�</mL�z0K�?/�J��r����N�6��T�6�-i�!8A��D�Ҝ<�f�Q�ƌ����}��֡��S��鹤�ՠa�Jְ,2.�Ԇ� ��S��n�1<�GE��|�_�^����p��M>}\:�����|"�1(~��m�*��������'�z(p�&ѳҸ\G�i�r2Tq��j���u�+g�Ѹq���� '���;�k<��E񠽕����[�xK���ag簾	�8��ձ%kkK΋�<������;�u�:�|����J�8H�.]��dў��c��ѹ'�osݗ������i����lh>�9IE����������4x���(yi���憜A�%9V����Z�c��>�;�����`W<.�k[��Ƶ���͛���u��?������d������ؖ�w�NV�e��ǉ���.Vd&$��ӂ��I�2���?v�(C�(���`=h50Lڷ>ц��XZJäm���h�����`�U��^�R���9.W��m
�������ǆ��;� ]�����>��s6���|�ڀ3Z17syp���E���)/�*�J�\��
����8�ha����,���)�i���@~N����s�]�^o�����~:V�,����'���??~��������PH�/���gƱ�c+&W���(n���D�Ï\����UL7w*gk���5�o���9��YLa���� ��k�*���A�&������TQӱyPF�q8PX�\)�%���4���p�*GFv�2�VV�隠�	a��IQ&�ӁSI�`	�&�YGa@]%<�ПT����	R�ΓN�Z����R)|�Q���u�T���3��;���T�Z<�Q��w��/��
_21�
�>�f��CF^��7O���+Y��ߓ�pLhʙ-ޝ&ÿ)բ�|��*d�`Z6��|?-t��s�`ն[��c��5�;��6��~�!�؛wGMe^Β�l0�^T�AE��p�` 
Z���|�����yȼK޺R��O)]�]��yY,�$�D�a�w��Np�s�_�]�ɌF|�,��b�ua�|R��}�q#��Y��eay�1�fD��,�p��!9����� ��6��3p|����=S�����"h^斾�A�:��E�����R���X��Q�_�n�O8�※0�=�s=�2of���;oJN�x�;�擂93jd��BIp�:fy�n^��}X��)u.�g�K��Q4���Ē*ɷ�9�H7\Grb1 �D�K�Ӟ�����v��Q�F
>)I{�LΓ?u�g̹�;u��ܶ漜��e9!\��S~�g��>~�����o���[�g����f������#9+�Q���P�Y����������exӞI��-�@��4G|ƅ+sq�p�p�p��^�0��(�~��q5���EPm;�1���c����������} ��y!Gi.�j��"+��o�>U�=_�;�y|���qq��w���4�f�_��}4~���`}_�ት��q"��5������#�%_ډ���7PY�*��-���ᬙ�+�E0���n�s��r��9�1��T�c_9Kl��2.��+O��n�_�T�C�p �y�m\��
j�6�Q Ge;�[�χ9��kJS�xT��o��E�a��sMSѿ"�2��P�#�G��)~���p3AuI����r�ێӞ���<lr�[k?����v�5���<;���W�d�6�|5W�xnk������r�>�|w���ZZ���z�N��� ��,,1aG�\)bF��:����J��, ;���7�X t�����,�
t�"��.I��q�=��r	���%��
�g���Ф̡`:����" :$ �/&0b��1f�Y�&by)����-�=u�2�N>�Y�?���ɫ�,sH94jVF��>��:����І�؆�N�x�����O���nB�*�\84���H��-T���QB�N�O����R'�B��/�n|,,-�Ç�2�3�j}9K�I��/�U[~jj�$c����ڌ��҂q��EL�>v�S�x��Z��eF _�l\��8�3���}�<���0�-Hΰs���cڳH��P4��� �,�Ei���#�*�?��\\�t�Ϯ�f]���k|8Yѭ����ŏ�$�O
�+[�fi� o�S����ҼЈvӱC^�p>�9~签(,����\��8TfEylL�X�_�SF�teB�Ŗ�$��co	����"'�sޑ��}}�?��7@��}D�OA�U-�܈�� 8c ���5/}(�E�H3!�M7��:�-	^�M��͂�:� �p��JH݉�����g�k]"L��VkA#�i��ȭU��:�8�oo��r�sۮ�?��#s�k�?�_�@g�?��8��or��g(2��*p5�I���Y���٧}9+���\}o������^���9('�`�R!Om�xC1o�;�i?�ŭ{p5��P�?��Z����se�6��|�!|^�m�~��7��1�x�#p�������(�8�8nȁor�����}9W8��ŧ/|�^�}����X����#Ϛ���u���͊8X�G�����͡�s"�@���9tD�Ï>�����;��Ԩ-���*�� 42�o�d�m��c�w�?�-8(�`ֽ'���RyX���uv,g,ㄞ�S��y# &:|ȱ���@�|�_��B�J��6(]ßch�@{����g	�"�3dυ�y&�?l��vfe��vm�s�mB���d:�]�oR��OL�G����K"�|�=�4G4L���lh����6<kG�L�I�S�����`/&=?���6�ƫ/>3�����;��J���-�/.F�_�d�������O�㕱�vq�+".'KʳY�7��a�+n��L����Q����1�Գ��:�y�|C��de����S��pX)svC��N�����럅�&զ�����5,����f�<�wy�ɤ1n��F�E��;��&[Ǔ�����uB��g��pz=��xz3 ���lb����ma,&j�&����6��A^Ԟ`��I4=�T���z��d� �YtL^?�h�p�(h2�eZ�u�	T��r�P̗�O563�օ�`#ڡ����q�Xw֨�7�BwF[��1i�_�0m�+͘S���z��~+�-�)o�b�Vc��� �@ӏ>&=���I�*�/(��8�?p9�,61�g���UI��}.�����"�QX
ɻ.�:߸�{�+�B���p��J��o���k�Y��]������9o-�N�d9[t���ِU�I5n�@�D��[h[�f����x��kوA3W
b?�!�m$P�}��#h��n5?�tXY��l�!����=�ѣѴ�<m�� �4�X��Am&{�*St{�9������fcΊG�b��޲�L�ڡ�:P����馋`8@��J�6;O��6;�ڐ!��	��/�~�sA��'���a=���w��>�mk�R�Zx���݆d�h��y��n�<6n���bK�.�����ñ�iMA;�(<c�(�Ӿ�Fb�J���-�K��o|}���������_�S�����K��d������|ȉҚ���q��%����\}:::�		���;�a�,�Y,�G幢%�Ģ?Ec�
���y$���r��絶��;��\ܒ�'5@��Hy�g��M��[<��}��꺯�mml�59Y�Y��C�	�q��+l48������i�g���>�@�=T�{�O>�t|$G���ñ_/U;=�x�U��x�Ы\_2�э���_Nxg|cĪA9�#=j6(�*XK])Nk� �̅�N����n� X�c�(Be�K��,��O�q�MY@esq��ϖ��=G.�Pl�f[[��Ͳ9vP��F�Ce*_,(,�p���`l�9\b�����,6� f����y�8��|껦Y��:��s�nl��L�9M�:*E��U�u9Yk\땽:��ue}e�����7�d}[N��/��g���?��O������{'+ce�:yQfɯ���,���@ib�y��|y��6Xl>r[!p��C�
U�\@$Y���c����1��˙�ꨢ�o�*L���lX�(��Br��*��ˠ�,1� a�V:_8�Ҧ���|������Z
�ȫ_9�ę�-Z�=���h��+�EV-��p(@C�����t2�_���
U�)�g�ܼ��N��C?�R��T<d�h�O�JXxj��PL�]���j�h�pQ�>2�4Ѧ̓�&#44l�ou�|Ne��c�̢�%�Z�C��~��L�Z&Ф��,s.���p�1���,��3�:8��z��8+t_����T�'C�����۬觛ў���q�,��`��*��,�e��q��)����+O)���&���Τ`����Ŝ~4�y�I۶$�, ��:G��&}'�qE�:�`�8[4<-x'|q���>��<��1�T�n�dq�J6����ɮ���ݩ<؇�Y�� :U��9������$���
�d�}d���x&[�H]3�<R�i�C��
���9&��Rvn_lHi�F������w6��|��A�k�� ��b�����#o�[���и��/����~��RJ�s�Y�i|{v�8<�4��ۺ�-�u��Ј'�JT%p�~J��6T;Y�?'rOlWi^x����ko�����x��Ab����ʜ��Ϸ��=�e���ڵk㒜,���+�#��9�axQf,��S�����g@_��|�����abADV��ɺ�+���U�܊�k�=.�[����q�����-�����AP�Ct�/�0qb�����};~���NR�A�Ǻ��������{��x��5D>����4���ɂ��P�t�����ֽi��EV�~
�u˺RP�SPc\m��~F!�_R����رZ�b�ȉ'z0T����#�|�R��a�ź����Xh��âl>?�_������	��o��3�ٱ[wm+5��W(�x���K�5�8m�B��n���(�a�K�q��qΞ��}�����"Rdg'_����ԺI�<�=������8�ߓ��:���M����o�6������UY�������������s9Y�+cu��0]�$�Kc*���Y��'�I��M�o&5qb�)�	�V��.�q�,�M��7�RN�[��D�X:�N�g�i�0H�UQxH���@>2��J�x, ٢�A��Ԋt._r6l6�.����(�p�~?��D�T|�B�r}͞'���>��� tx�+F�+l�hac���I;����S��j��5����Ə <��g�X���OƏ&�ar8��\�?S@�}�(��X?��3�=��k�2�TѼ�ld��Zf]��y���r�Ò��U���1n��ٿ�\94�5�l��tI�,�'������ ����^6o��^ ��mY�BA<�[-�#��q��V[�W0�dI�q��l�73g������۷�I���DY��AӬH���Y���'�l>4=�� {��2���%�!)�穊�b�mXl��O����/�pN!������E�+|�S�8��ۥ�$�bAv��?�K�x1,��k�UD$�b����x��@����<�q7���q��GM�)�E�
R&=�gp�@�\U]R���0��V�FhA�o���Mt���v�D;aj羹�
���H�*���u�p?��;`<b�����	Gl-��g��_h��Ww�Q�4�<���]��R�#��B�U��t]9�Xm䴬��}�d���Y�8����x���^׺�한�&�̡������k�'��X�p·�	��>ɛ���~p��W�4�p��_W�^�qaqp�ձ\�y�#E��3��է59iu���8by����"&
�V�P?%��|�¥q��󱦹͉&�"�/�@^����[n)�Ϸi�5>��cU�/K��^���߱��D��Z��rVx����0�9o�����S�w w�u�E5m�?5b]��J<Ԟ�rNئ�!Z[��~m�y��g���z`(\���s�@4O��ʩ\��20! 3k��?�+٠+9�C�i�O�����b'��!��"s�?7�7~��_u�E3����g�%�R�Z=�KK�t���E�Ts��~�KDuTr��P ]�`���a�Q��gR;Y�hU):a�Dr�F`GT��Hi��S͵+�k����z���o�j'뙫�¡������d�ݏ�?��������,����藅"N��2V&6lB�p�&�9dn("k�#�ߜ[(p�xY'ؘ��u"���f�1�*Vd"��J�(MPDq�c2*� 4���dBؖ���\����̸���
�c=)4�]px2) ��|�����H���M���-�~�N1�9c���!<B�G9�L�_>f�$�x�+pV��<�C��1��׶L�u��oU�&iz(Ppk��#/��@g�B<��\��"WI�TnG��?�b���Pc
����������hw0��0w��w�/����1��p���!x��J������eB��̝�i�`���(/Z�9lH#�f+u�&�D��:.^�ݦq�K}�q�*��풂����aI�t\F�Ap�v;؞�̓���xe��1/����_����>� +M���X�OB���C����2��m��(��q��϶Kݖ4�Ŀ�E�US6=x��3�7��)�y���ͅp�2~S�a*p���)/��%/6��dX}�" ������ly�e\l�8���q����E#7�1��-|zs/�V���s�w���v9[�>e�\l&;��W��P�?6��5߉���H��)�U��͏6¶�с�z��ϡx��Wl�uЁ�mv� �T:��¥t�[�Y�E���-�P����k������9���&r�w�]銊eB�ˉ�y:�6!��3���o=����1�2���z�v0����Ɛ����E���� ���u�M*Ư_�L+��]z��ċabY��ƕ������x���͍r�����>�D�)[Ӝ]����Uy
����?l|�qN8A�[���/�`��G��9���؃�|o�H9d��5������5?R ]pB�s�1���ǀ����g�$.�_���.�q[n�?�3�s�7�<�'K;BH�s%�X�Wyջ��v�CsE��Ǽ��[~�U�#��1Y��b0�rzdoJt�	!����Z�3��]C��`�ԮK=�s�u&%�VnF��������g������"7�<�A`:�y�ߝ7~殁5H���8����6��{)�y߅�h�����������P$� �}����	�S랢(����H�q�8.`���f��u�s�Ɵ���J�d/�m��"��c�e_��H;��2�v�����G����5�ln����1���K��xu���W�s�������7�7�����_�?>�uo��=҄X�k�`��U����R&/.(x��M�#���� ��a!ӄđXՄף�185��N�
 �fӂ $T+q"��bL�C����Y�	\�8Szx˙$�C��z�w#E�%X�C�o�6	k���S9C~��R_���t�n?њ�Ù��2y�^@�6#S66�ڸ���mB��MI�67�u���%�\�cx1|��	����+q��m��!�u}B��g��U�@
�2@����&��������t/`��3z�TS�0=N�C��x��C��;�3#C��	�����o��hA��/A����p�g��xbr3qe��e6��/�n�W�)���*t��'�I���V7_��<U\^=�7�s��.��D��?!d
��a�Yass�MЩ���s��Ն�f��$�.dlX�b+̫R�j�u�nL!u	�5p��1�Fʠ�Q,��d�}�vt;4B�2����|�>�l��|�p��و���1��z�kd�2[���'�.��-��HAl:��Ycs�G�)K���}~�A�\B��ܙ%4b��vExS�����q~f�|L{�VK�1B������g��_�BJ�ЖR�����D^a�:�_�i�7O�<<������~�h��D�7e�Mx�-�r�)'��~{#���1��~g��/��n�3��释���;$�ol��$����ĳ�^ѺUo�֥�
Ӹɷ�H{G�B<�c�Y��P��y9_�9}V>�@�a�QRh#��+R��C��|5��W���p,'��ŞH�8���N�Ud<�r"'z��(1�����?�8#�n������#~��oo��v�
.��\��!�],�ϼ"�Ex���q\CwU�*���@w������L�]�_ߔ�m(�aU�z��%�����5�ٕ>��|�0:n�XS�7��#�]� ��[���$����F?�=���(���������?��w���tJt�Kn�S%x�s��H6������τo1>��3�#�y��		�s��?��D���	�ٷ�<vD���|W_�[��8d1M��:�Z��e��t!��o��M��<<��!�x���L��ot���ux��� ���?�)>�pj��`:&|��Z�;�S�����`A'Q�V��.H�1���j�5N2��_\_/ܼ:^�����^/�xs<{ucl�����?�������{���>�7���㥱�h˛3^�cH�0JQ��ґJ1��o�l�M��)�>�%E�[1% /:?��N��F`Q
el��<�x�5�MQ`x��#
��7���az�%�3!�QD·�0��<�&@U���^DTJ�äk���u�O��G����
�0�G�)�Q<���_<�+�R�@�H>t%'�A��|��˾e�/�3)�e�3j����;~O?�O��MF�������/] ж��̏�:��t;��3��7S�d6��Ld�GK�􏤫�G~E�y;E�EV���
@z�6+֟�w�ll���Ɓ��lv��U%
�۰��3�S�a�1'� -c�[/b�}&Q`C ��Շ�����'�q��46mx����!˪ٌ�uP16���x.�Ԯn]�!�ȡI<���λ-�v��q1�=�7��вlZ�u�yD친gQM[@n�cCc��_��*�=E��N�|��i$�18V9��I���ޘDƑ5,�1-ٵ��?���������gr�aL��R¢�Ƙ�:�h��%>��ƥ|�h�&��c�Yi���3�Kt����6��^���e@T��y/����$��'��_�hQ�:�72B�}�-�pS���aݩ���5ڭ���lxl��h*�.�w��A~���\m ��"*��38�дY؆.+Z^ү�L?����T�9ɉO�%�5��>Rh�K�٠
��-Ap�-o~YQ}1�n?ۘ��͛"8O�/�9V�4��9,^&I�~N�I>p�:�5n����.�c3�W	���Țg���[�pQ6j�����> <��R5����F ��-�!z���-ݾ�g�Pp炯�s[���z�b�0���+��ˑ�a!�:>���LmV4~k��^�2���|$������܁�r";�D�e����֘�#`�S�sR5�W��M�ãmH�+2���[q,}{ج,2D��2"o~�!F����;n�n�<p�E�1��m�A�l�K��/d�1��$*����M^���C�r���+��b�>V�g�u�ՁW�U'�4�q�|x�V�3�Up����<�`$'�,�R�ܯ�jn��/�`Ψ>��|b�ɾ��I��Q�s��s���R�M0����5��Yk��G�4�����+.m��GG��0�J��-�y��x���/=;��yyܸ�66W��/������?�7>��ḿ�Q��M�rE,��@�N�s�'߁K���8rݛ��<�D�yC�y��jE���6�^�l�
N�8R�KK`I�;?�a��4��
�G)��IcV]��x������G�\DB�D6��j�����V*6�
�OT�5�=�S�!}��u-���j�G���	����q��%��-;�㒜,����u-VG'kg�y&�DO���D=�=��Ȩy���o�2�=Z'T��};�9#�K�,ڒ{�e�3��7|qLy�H�&zo��3�J�@������.�G?*_��ֵ)h�}�<k���M�$��`YFo���[���I��
�wѲ�R���1b�<��.՜�|@G��F�t����­!1���Z�k�
+ڔ�(�}�쉞l�8�'.{<�x,/�]�xQ����ih�~�����em9+u>s;����4z��^H�/��2B����?g������j�z�1:e��b,�&�B��-�fht�����l}3O�H0�·�ʷs�8��#��=r %4ݖ��JW��ȼ���w�5��ʢSyxA'��I��8�������~����k3��۶�	�bƒ���jX��m6���K���[��_Dt��%��]��:��.�)F�i 5�f,Jv�!��=���z̩����`����<�c"�A��=���e��DB�gB�V�L��}mjx�_�lZ��L��3�>,��z"���m��b\�3�/�7r�':}i|ޠPVcO=|2n�,�	���ho�} ���9�[{d�*o����<�6=q�v���hɛJ6���=�v�-���v�_��v_TB�q�o�d\y]��˽��U�8�-sR�q�D�ވ�=��4ߤ�����N{,��T��7B�3W�ދ�g�Kp.�=O����1~��//kܴN�zD�-������"��(S���X�m;q��C0�vΥ�*�VNk�t��PD/\���k����q2�-���ïB�%����z:rl�E���'� �z�M2�:Yfy�_�H̉w:�ȑ �ÿړ���h���%؋��J��̯��xe^Ԝ�~�S�>��!�ܐ��=��=~�:8�)�/J>s:����=4�d��Dh�y�5>�]�����O�1��[JȨ��/�+R��z�;�����ɘf>J>J9�<с8���7��Q���|�A�[�|�bNֺ`.m���W��ͫ��K�����؀仟}xzo�`�{x0����=���q0.�156�C9-�Z��;@X�1���#P�t��a�N��)�p�'��erB�3������$U�h>E������h&(g���i��{�$V61M��i�>��r�W��a/J�gO���(�eC;E���r�<T֯T%�#}<�#�	,9d�Daul�+l�~\�{�c��zFh�93�(������M�<Μݬ�h�.x�a<0���(g�x w�Y�k�2��hY(�1F ���1���1����O�[B�1���Sqc�1��Go�C��?&�#�o�ɥ}��M}�y�d��R2t�����q ���3/�G��=ϕn/z��u��;c��I/�'�d����J�NV�ܑ/Y)89���,�Ȉ�|<���d"��-S����W4,����_��#�w��7�>b#�f��|��[<���"{�'|����*��`,2Ф��+x�Y:�>�|!��m����x���2��%OZ��/�����~���]��\ߚday E��i���ѯu>	ֻ��������&�2<�7��t�I wd >�b,��D����!W
�p��E���k�M��с>�~��:�m�f0F�������f��xG��U^x ���%:�.t7��?ƂE���9f�� �ś݈�0�#�Q��mgl,}C2����9C�^5���ec}�gc�pk���%.��?t����'��[�43_�l(�&�tK�<���E��Ilz���m�h{��'dLh��޷��X@÷�-RƆ6�c���/dxĖ�V�7���	p�)�fV8���7S�!��n^Ӧȫ�@�r;�|�_��3��;r�k��'����c���1�h�l��6���o�k!N���_���6��/N�`g���|C
G|��3�'�{+�*G_������6�|��N��`yhM<<GX��9�V	��Q8,��?l#��Oe���t�l�_S���Sƃ����2.Y��"��UPt�)�x����e�o\Yct���?x�sU��#����D��Ӳ�`���� �xaM����2λN�#c����.`�$�10����h}4rS?-Ҷ�*��Gx�e�mmm���u���p�|[��\y�f�׼�b�}'L�aۆ�M�_��'}���n����~�]�l��B�s"/�2{��ƈ]���<�o2��?�g=�ßS�	��G�&;����Oe�xp_듈\UL�G�M$2����5q p7�z${�^�9>�9N֪�p��r��Ƴ�����,ۙ��>?=R��&x(�s|"ú�����",f�YXt��8bR��XJr� DAGK
�((�Ĥ �IfC���T6��'bXr�R��"(Z�X�y3O���*�R4@{ԽY� ,6Kve,��k����Rf���^���8� � n/�2�8Ub�ƾi�P ;��`�B��bSJ�C�D��_%Z=��<d��l9+��/��d�C�3�����������#�}�E�V>�K���&)Hy�I�9년6����d�/�i��:(Rs�t�Xx�$!��3m��x3�%*Oh���jh�@;'��2�al����+}��?��h!W�|��m�i(�g��Ȋ͆���]�d��W���\�f�� �!anyc'��1�h�:l#C�_����K�f:���仯�\���hxs��"?�@�n��1�N1b�ਟ_< ��_/oҒ��^���x����6��Y���7��@6H譮e�8�8���#޼8����~U�:����$O�����+N�O�2^w�h�	�����G7�#6]��C�l&cK�|A&ՖH@��d0�S2�E�|���D>��f�1��|�#㢟��/�t��g��f��S�\e��$|�r�ƃ��Ц7�Z�LD��l��DJ[6<�F�o�p볯@�~á3Ȏy��h,�3��]��������6�骊tS�c�/l^l^Z@�?o��g����Ϟ�$Q��Fg�ɤ��`��m�� u���U�ԛ�I�Ad�8/6U����g-��?r�զ��U<�2�L_���#o���l����,t� mZ#�x�I~�A?��y��c�z5r�ʱ��A��tr�uF{�5�)yd
�5;C�$" t��H:L{������,2᭚G�8���獃}+�y�56���-���P�[�'��6`v�v}�����~��H�5��� �,i��/6�I[h���_��-鎃:O̕i-+�|Z�+[G%_e�gFQ�RҺI?�'��N��g�f=S�]�ߞ{�>Zч.o��:
owG��=O�u�l�p[�Dt�X�>: l�@�r��|�;���{�^/��#A��3<�qꜼV{ᇿ�����k���z��u��J�E�Ӯ�ĮfMk���p���iú���i�s�H���ʩ�1�>���h�]�v�ት`a/���^�g�&���.v�k(z >x>"G��V��I�D��>S�L�]���������S���܉�˻��࡞�1P�8��3mlHҟ5pwoS?��_�ck��؀��Gw�[r��d�p5gC~���6�i{>��heP�p�D0�Y0�%H�&�Z�,���|�:-0pt�1�|��������g(<�8+�����Z���$^%<O�V�Pƀ���!CĈd���tg��`a������қ��M��&(^�;&X���˞�aR6��ń<}�B3��ո:G�2���svWN�6�0�� x�
Oh��q�H";��X+���7<�9�/�q�L�qoX�EM�,�(���H��n��/��u%��>+/���<�	���j9����T9�����������_4(�`�#��2 �M�?]�(ﾐ"��7O�?��IAo�o�K����hdQ�dU򥝆�|^muh^�WE��*�cK
������.�������6(v6��w�$Ѓ�y�`�v���"|�+�*zary�[���q(���s��o2��od�F�i)�e�O_����� �:/X .��n�#2���G��5�lBX`ៀ�����G[���Sc�g=��1�C�����V���	2~�"�h9�/���R1��ȀL��$�Tx�z�I[p���"����3���Ûa��H[���c�`�	�3�L+AN&1�ឹ{b;kܢ����'r�
��;��aiC{����sA��/����3����考�Φz��1�Ǒ�[vD �6���4ԩ����~��dS;��g��	x�чvn-���l � �6�hF���^w%#�����ӫغ���X��y�]N��?�t;t_�w�+�X�Wu�Z��e�y�(�	�1%E'|r�lx���y꓍�	���o�Ѽ)B�qaް��ae��|<9�dj�e���J?�Wx5[�gA�'|�Y��ʨ��*v���__���ʖ��F�#��C=�'|���ᾭh̵3�n�#�K-�G����^x.��h�)����"��~c�ʢ��Q��?��Y�u�e~�Ŷz��q���ؾCJQ�_Y��S�iz�Euk�]�I����q�q3H"�bzя�k�[7���m_l��[4���{8���ڻ��S|���'o��=�~1cI9|g>A����ʨkg�ˉ��o3���1ԽG���̏�"R����h''z�o����>�$�Z�8GE+VU�2G����d?���K����>Pc�.L'(�?��¥1��xE�<��@O��x|�_���?��z�5�aEy@��+h�.�2{5�r�͂o^h'Y��p��)�v�^il���X�X���$��B�F=g$�7��Xi�1�劏䜘����xMe�X��4A#&��`&t+o�y�yy�V��c�oew��D�i��(��`������:��gA"t����u�n@��DGȽD�PS;E��wN���q�R���L>W+��x������>0��yk���9���>�C�gC�������;�.qF��2��1Ƙ���@�����ч��G�o�Df�B���]�O�aA��}���6���1"х�,��	,]�l��i��j�e�_@&=A��Lq%��7>��O�U�š�3MN��?��1o�8��.��=��	��c�a
��VDuo�k�M������-���xY桎m�X�述��[�	L9Y��U㧎�����
��O����z�uMd��#/�I��<�O����`��/�*��k�p��^��?	R�7"V"��:����zAt����9�l�zB9a�W./-�0V`��q66:�s���:���r! 繆K��	��w6��B��f�ZR��Xpk~���а���`K�Lڵ��ג�e�|ϸLSsv�d#� k���ቡ=s҅r�C�Н�.������ +'��G Ȥm���Y�M���O�Jz�E�H"|��~�Z�y�B��#g~5���F���F��׭y=|3G�!�~ۜ�HĲ��2d���o@9Y�s�� ��y#��8>�x�cR�-d��."3_W�7g"�lZ����	�W�	v�xF�.��0��c�e��)�6�Q����DU]Im1.���<��tF����iJ�^���=�:�(]�O٘FN8!�EPi^X�%��M�dg�P�X[3�oP�9yz���-��1��͜b�!�^�?�f�t���[�C�Y�4��c�d~�>p'WX6��nH.~����x���n�'���P�ŋx�!�c����P2�=!֔e;W�ŕ-�&6�u��wd��S�e�5r�p(���M)��l`�;+z�zB�����_�{$�W�w�.y�:d'|��K=�k�n�u���#�H�9/h k�������f��C�[6D�CY�Il�i�.]���R�X�]��v�ē ��W�cYrq�<��6�f�:���j&�����c����n�4}˜�����}��c�۟��qa�H�2��zV<�-���"~�re�h�����5P0�I�}ʽ�=�;i@�K�eٙ����=��q|�A����G~f0&MJ���󆎜R�M)�R��	��Aah"k2�d�+>��Q��Z@��=a袨fL����BǄC��ݦ2�eR-Bpo��"���B�].�,��4�F�����u	�C� D�bؘ��Qt"Jτ̙�����}�ǹ| ��E;a&i�T�/Y&/�(�ό')9t�K�>�����D�Y�F$L8�G���LƌQx�.�Xɡ��~�c�D����{��d�.�̆e�,�#gj�-df���2a,s��t,������
�3�����X�:U��<!MJ�W)r/|�l��]�;+~a-4~����[b��*�ت����F ��}6T���F���Ü�r��yQ����\�g����/"��S��Ǥ�iƔ��U;�Sδ�_�$X�@���[���/�����4�p��z����+����4���}��]G>|Eg����n�g�lg1��������Kd�}�6K��4���r!�&8��ӷ,�#��:��^���%׾z���/��E\�g��`!���hz#Y8�A�����w��y��}�U��z2A?3��G�YF	�w�1�*�:���kF����~Ϻ�J6)�Ml,<Z�>�>�ZM���|Qr��&K������qd���p��D{���}�^�|�ʃR�p`��́�MY.z��!��64{�P��+�m}�6póu��g���P{���mb���k{�d��rx�J6�cPz
m�^^4LG�e�Q�9��w黢�V���"�M3�@���żP�^2���ʟ��1�Zȱ#�U:�&�q����M����GK�������1�x�_s��%=cC$<�����i^`SԿ�m�г!M�����.2ˍ3=Q�`���Ⱦ��v[�Oi ~�q�67�^6�`p[�96-����Ehp���5O��`�-���}%�W�X�V��
�'>���͵R���2�?k�u_��y�X��qA3�F�Di��ل}"x�=�ڢˌ�u�h>Яs����rX��m�ײҙ�(�XOgv��hV����C?�/Nʱ�s�a�'��e�x"�bH�e�ɑu;������_�r�ǌ/�l���
`��K�
���P���R��Ƞu�z��?d���ۛ��1��B�% �N�Gp��:�車J���}����m��1�k�V�,|D���8�Δ~��xְ�
Dȝ	�a�s��{,���@���7��?8�BEG�<3p`�L�c�C�B�SQy/K;W��5,&\��,�,0ìrf�Ǜ����P�/�Ջ ���|UX[���M$����Ai%���`�r�t,�s�����I
�����K��z=��^/b( �8�q�Ͱ�[
`Y���~({�<�zQ���^;�3gR>��$)y�ՆA<�Hl�� �ᣃ����&:�����3\����4�c):=x��#�'�M�V��b�4p��A˭ld{C�$�����`���@��J��2!��	�mZ���z;�d�����?�<_j������T��)4<��p���Һ�E�3rDn�#bX�;�2�3�韣��,^6x�d!���<����6�2�4���[���d���I_"�INȡƋ[B�ǖq!*���Op�����mz1 �cxQ�q?䗫�-����Y��LQ
N��Qn��L��"�����*bl3�fX����J�}��>�'^����f�k�c�x��gy�\D�K5�q��u?���E&/�,��//�]���K��MX�*6�4������qm'�cpz�;�@��ü]/�����c;Y���%�:��ʌC��/�r||�s��E`�T"��n�[�v�85������C;�-�fZ��/�y_���8Pf=����ӗ9?�D�<t�������:p�ò�� 3�ןC�E.��͸��t���cH�eAJdnK��;����n}?��ž�C(��q�WxFo��85�7N�1�^�Kv�#�f�辥��'+W�Q��9�`9ÏR�0M`�O�<d��7B܊n���Z�6��6�)��6��:�G��>9ya�m����d	?�D@il'��8Y�6V���O�&c�]��2�Q��q�S�j��C��ɷ�����H�3����NlYO���t�l鱟}}Ʉ��8�~)���P�����"�*���L�#���zƦl�ʭ�e��n<��S�U`���.{����k����ں?�?��86�x]�u��,�5��	�tQ�Vd�]��~ ��6W��[�	8�Ƽ "W��=�v�j�ã�������y��u��L�CtT�:~;Y�	���uxs�ڪ���B�ս�,S�'m�)��x��3'�Iଯ��0�W[��'B�,�
���*�b�Y덎�����bl�j^@�2a�(���ef}G��+��.�>2nk���^d'Z�q�V�H�h�����άM�\�U����^h�2�O�]�w�s�7����T1FX� �O0ņ�20����-�Zp*sG�P�D��~���D*\O*t6��g�<�_�FV�ތZ�)���D�"���"Y	2&�.�3����>�i0p�Fv�~��eW8&$)�en�Fa߼&��E}�1ƅ &��������y�z�YD͟S��?��_���8�Z�\���,ڤ��/��O�Ӯ�h��n�Z^�piC�Vds`<5���?1rF�\ue�	g�5u���	�&�=ᠥ<���#9۹��F��n^��_�GEdV�u�w��?���hb�S43�16ԓxr:2N�
8�{�(=dl=�l(��\�C��@h����@Gx&+�Sp}`"-xW�'l·e�s@��������z.�>������C�Ey��l|��i�N��{/��π�7�O��Ǡc�R_8D�:gy������S��)�z�Ү�|⇇ѱ�C��[���#�d��%9Y����:�����^��1����l�1���'`T�~����/���y�Y��V�k���\�k]�?�cSo���U<���d��':�cp�?��sܲV�w�=l4�ɡۺ��S��u$dӅn�L0='�G>\�eN�Ɋ��1m�ˆ~7_t�Ǆ�
�҆�;ˉ�5/��6,é-p�����qS�폾y�Q�ˏ~�SeYN���z����/���9��4�f��r��A�+Ս�r������"���Z�6��w�
>�2�*5M�o���Ɵ��v��{�����v^���t��t�e�U�;h`3h����J��<���v��	*� �>��� �R�='�p�9�o��9�K��X���͠��<�:L�o+e��x.�#�/|���ǝ��Lֶ�:����_�����E���#��^���JoJr�E��w�[������c�5[�&d��D?W���\E�J�2���3~��X��_l�ꡩ@�x�"�Gh�;���D��0��� �`SP>���=&��[<ڑ��F�@!�D�����o��X�,|�]3EN�S����qWq V#ɢ�K����"#�tG9 coBg���C[r��
����z䱠�l��2���`��U!:�9��f����_Nj��+F��yބ7p�V��8�ZeS=Ǫ��������)q8]V�uK*��q_�`�3��LΌ4{6�#*">������0��w�    IEND�B`�PK   �m�XK숤u  �x  /   images/598b2a10-ddcb-45db-aacd-6c87816d7084.jpg��eP@%:8,0������:�n��[p� ����;�-�m����j�ի��n��u�G�����Tu�-�m��HHK ��� ��m�� ���/�u$T$$DD�w((Ȩ�00�ߡ�cb�����BGO��>>>6!.>¿�HhHHhx��x����	�A�#�3F�����!������ pHp�5 �W����2
*�;�� x8xD����_��_������M��7C*<v��Tj��.|��#� �w�D�$�hh?��sprq��򉊉KHJI˨���k|��26153���rrvqu��{�
	�O����������_PXT\RZS[�ohlj����������_X\Z������?�sxtyu�������� �����?>����(�����$"�G6d\�o(����Q�D�r��Ш�(_�9N�# ql}�������P����F��y[` ��[0��E%7�3���p<����%�B���[a.����@:�)��t4y�\u��r�ƅ�i��<�f������\�����C����	��������/6v|��i�����%gΪ�<����]彩Ց���������Nr�P(�~O��1I~vs��jԵ �8J�_�B�y!س��_���[u��#F6$4�!���e0�� �4iN�6�\�ۢ��fTT@���T�L�fw��C�,;'�����S?������wd���;d�b�l�klI��*O�
�d���7 X��
���|�A��CM�}���G�H�k�|�&��^�N�~�}e��[�_��t�K��"�	��0N���Ss�x1>�#f6�}jd 0����r�𔏼�p�c(5�k��NJ �rh�Q���8����,�x���J������O(�����F���C�Z��Oc�s��em����R'��p�C.`��i}�ZG�����'�L�e��� �{��M�bmb���nU�����B>$������Xc|w'�W�)�:�2��[z)�D��|�ZS����Q-���o���U�������:��zri�iٟڍL�Prex�y�c�t*�Ҝ�Y��	{���6>��������͋m�2c��ja(���7q�yJl�m��� ����?�F�d-�������Vʹ)��qjqGq�|��Kr\Q!���T~:����ˤG<���{�%���/�^[�$P*lQ�p�炘c6��"\�C�Q� �m�P�	L1�cp�i�>>0�\�˿��0�K	�2�1A�~���ܞ�\=sVI��!w!�슬����-Ȩ72��@��j]�m�&�x!gu�|��cb�kJ�|��0B\��fZs��K��	�IB�o\�J�5�*f�H�E�}�{�w7t�lS5		��R�����޴����d�/����A� Dv�D?��A,�����U�ٚ���ś%E��`����N�åŔ~��AD�+�V��˼i��G(u͒�f�ӡ�f0�UCts�6��h:_K�y�\�^�+q�E��/x����#c���)ψ��������]l#�q�ʡ�����~C�u������W����Z���j�8B�/�MR��q����V�
]���!���%+�����)m��¨��j3|ʽUx3�X8��C}l ��R$��6�����{%6�Nb�Aa}A���Os�C���`B-V ϫ T;�p�w�s?`��=ݙ�Y��>ю�w�x���\l�Q��-�h2d��m�[�2^A��y�G�6�qz�I[>(`��d���e���� �Q�PFTɠ�p�Y��28�19Ӭ�F�a�(�}wR'�iv�@(�P?<���.����B��a�d��4E��/2�:@rP-��h�:�G��#2M�L�r[�[�ٮa0[�-�8ҹ*��g����]�����s��|8 Qb�L/��<pH�;j��j�-�4��/�YlyY ۴FZˁK����H���J^$;#:�k�m��%`�z�N�B��_�?v��c
A8.����T'��;`��T@O�zL
՟���J1-�k��·U�Qw��i������Pe�3B)�J�����d�;!H�3�"7�7DVIi�K�-�j
�� �8j)��5���^*�)v���s�=��x܊OɴB�
<�w~��6�ڴi�(��� u�b�7q ���E5�*���_���D�F>v��.Gݴ��
��N��tG^�R#�)�K��¿8?E{Q���l�-7#m�D��T4g ��̎��c�fۇ���3w�[��į�N=E�Lp[]In6��3Aێ�0R_g�T;r��a�{��<i�_�lBŖJ��	����s�G���&���C�2bZl�a�4�ԃr�E��%�n��oj��ncj�� ��/o������3�5A��1��}Ɗ���D�E��j�zE��� 
h����c���� �+���i�@�U��a�=�Gc�I���Da��;��Sހq�fW���	����m����({28����:D����Y(�ʢ�����l��K����o���T2��]�F@��=���9%P����,��G��8?bQV�>Ʌޱ*M�q�W��}����Zd�����p������\mj��&c_Zc�!-�p=o���]q\sSk����df<7sA��f����ŧ�e�氳e�<.ܭǬi�l��	Ŷ��(�i�EB~ȡ<��չ�A�:�ӫ�2mm��/�۽��H�h�fL�+��7�E>����  ��+��
S.�L���d�dF�q���O�l�Y��C䛿6�q���nϱ����+�g9�q�n�	Sm(A�޿�G���y��Zis 5�c[L��8/r>�u�Fv�8������q�����,�Bu� ءd�|��f�7v^���\镭����W&��~��(J3	k����Q��~�O .��e|)+�X�8��
y���S������@=����,{4+�i�X��ɤͶ`�S������*�&�f-/ŗ]t�6��\��O9k�I�6�(P�����{֩���
+�%��X�L�̜�֘����A�J����(�L�Gi��S�>�S��Bf�/+l9�ڻ��;���� �t�-Y&�*�Ǌ�����Ȉ�5�a���1�8��n	�ȚнL �6�7/U2Si�D��gL�S�����4�a��S�z��n�Ӷ�"��M����r��kJ����7��uf޼�oW8$/ߌeLo��o�|6^L����.���� ���M�Cr%Fo_Z�Ej�UT}��5�R;�^wX�]��ne��O3��@-�|��ޚ�h��9�8B�-����(�b�k��㘑�����M�I:C��Wj��9�^���ޝI)�u�ݯFƕ��:�ͦ��ҽ���#f�Y���f��O�b�͉B�L��v���,�{w[F�[K͖V�M�"Wt�ӕ�R���m�!['sk�7dl.�|&lږ���e�j�I"�g<K����C�|y�`OUŒ{��#�b�F�tawk����q�;�]0F-�A�c�ZtG�\v�~��/��m�-�3���5�g�d;ʗM~'�sƠfE�v���ߦ��|[v!���u��S#U�����Ȼ�v�Oٶ}C�;9l_�c�����~d��#K�Vb���^S�ć?$o	�Vm��,�ǳ�KVq휾�U�rHy�E�����˂#�E��%%T�)

̋Q�D�!���m��]zf���ͺ��sL3~�Jr'���ʟ^����ZYBBg�ʣ�PB�2~����Hxx%�ܿrN�8?C�1��rv�W�g��6J>�x��ߡ;��Kc�цԉ=$�g��2{���z��S{�57M�Y\ʗ�v�e��+��ԏ���g�J�ER&�T�_$	"\o�3ْ\���hz��\!s�c�)�0��@P����9󭴕c� �м��Ǩf�T*Q�/�ev������-��I����4���r	rR$ȟ\�`��eq������_{�Qh/�����WTb��FĊk���LM��mw�Eg$��SE�{в�t�]�P��H-Fs&[�i����͌�]����z��,F��sk�,��ɷHW{�pj������	��dǲJ��P\�j��<\��(��v&W�v�ļEy�i�H�
{��l:>��z.�a&�b$�i���س��RG֫:j^�м�:��׊4��5���oj`#{�ճ�ה��oG|�æ�������-�p=�
s#b�k�P���_�v.�?�g�o�%�H��/��|FW�H�� �;J[+�+������V��p��K���䣣��e*~��2���R��M��'�#����ȋC%PO���'l�}ٯ[
�o �������'.�_�\��g�Q`����gyR��>�K6 r��G�J�W  �	9,_�D�*y���9��� |�����
3�g` }���k�pw�����HS|w|9v��t~*A�Z����wh�xM�?�R�%ט�|��>|��$�f^�B�c��B�^b��%�r9�뢠Oיr	U����ͯ�T�(����+6�A%e���C��a����	ko�v��{�RX�&[�G��J�QG��񋼐�N꨺�h�_�;�b(8�V���4~��z���zC��j���O�]~U����Uz:�m+��H�X���S=�뉰qc����uU��/6�E*� �Y9�t�r�D`�/R���=��5k��v��;���$H��}E=��Ys�X+c�v��+��^[PM���J��%�vD�!��Չb(�Z�}/B,���[po�����9�
"��i.�Ӈ>B\_�%��1f����\�݌���H�O�s���"\'$9��I�:Ps5>�?.qΙFR�_���ى��,11cz 1_L��d�e;�$�-���9�1dDu��5.6���7�h��ȶ��"{���c��OG�F�>1��� ��4j!�h�dMj�ɨ:ϰ}ʆ*��u��?Rz5�!�������u4�/~�1s;�Z���=Q���޳A�N�Ā�+6�~w}_A�{�o5�|?��q��B�6|�|�?�/klƤ*�f��g��R��m��yA,�*&w��-����s��u��L��-�����:0�9�����\�꒗��ќ,8�:���y��!��p�d.����Qpu~c�9)���<%`���#�e��?wN��,��xTq���b_��RD�G���]�i�9yG�E!=���Zp#�fM�{����g�C�C[vhӉ.�v�n�F��<��k:�-쁍^�Ȋ^Fy���܌V䔳��@l�Cs�$��#�
��N\�n�G�N�Wb�dX3q+Ks!��D��/m� �eMfz_��5�(UG]���1���[to��`��'	�3�6w<~ c ]ldUlά92��3�6��a�@Om�������m��/Ⱦ�׊���jI�݋o�lye�p����`��$]�5��>�t�:D����N46�s�{c��W.�tҥ����5��������\��(m����O2�o�<�V G��K�=�l���'�%��"�����xyAS�H�� wn��_
^%l�p� �\f��/=�OSfSiIǴ�+y�������URJw����������;�D�q�iS�S�^K��m��x����8;ZU��v�zo���t���0��a�G��D�[��.d!��y޳<��,�n��$�Ք�j� 7�ڐ}{��
�Ⱦ�����ڴ�Z��F�g�t��	w��Q�Hx�ſ�k@�#��`@o�iu�&B�n�L� 5J�0JNy�͔<f�M�߻Ϲ��x��"WM����H�\����%�x��R@���~o����/��g\,���hf6����R|Đ�f8�.���E��b#���sμ�=ƶC�ԑ�c����8E��Գ�5/c�\EU�p��tCò�΀��׮%lc��}E����fV�=�9�(�{KX�{��0H�m7I?�-�8��L�s��j�j���{ �sX�S�8�e�k(��˞-��+q>����d�� 7�֯SW��qPsC�؜�>���.^��1��Ep��3)+���!A�u��gn2�BG@��}��g��������߭��g�D�߲
m�V��3�X}���ѻ�Y��=�����$�5@�����(E2�E{%��m	�.�u�D���_iC��� �g�ޜ��:�H�n};ǴyS������D�k6[���'Ix뤓���e�<K+�٢Yj��RI�F�J����O�\�}��#,����y0oъ%�Y6�MHl��@�ן�$�@E7k�X�kŨI�k<���ZR�����E]��ӿ+M���8wdޯ��V?+��bQ�p�ٽ0�0��Y��j,��� 
��~�5��p�Z� ,1�q����L��N�zm��c_3�Ě��a����y�*vz�K�X�	�;�Y�_i�Mq�%l#�+�q�x�?�g���6Qv��� �$�֗�O�hi��M��djCdFVӶ(�4v����枆!ޒR�"6��_$Rx_f"����jl�,UsdR�)k�����C����������JjIaڟ_c7�a!��MU���z�\�}��'�_A!�r)�RD1�����/n�ZC���0o��k�������/��(�8,�H6��A�!a�!����,��
%�g7�0��y�y��7�?7�2IZd/mk��kz�[&�4���g�ߝL ��"[X�8����������M��5��Ҁ�h� `'���Y��0IL���aܨ�ӓ����Q����'�L�&�L��g��m��ì�6���h�C@���F!_�<RCy:�]�Ȧ�J5���_S����4to��f���k��{�C�4��O�?W���"�P�p���Id35mab�����;��UE����ݭ �^�^y��Mb����>F�3�ïJ���9���-��5+�P~ %?�
����۫h����]}����̹W�a�ozP�9H[�7�9{ر�s�h~�=���yE�'e!.�C\��$��J������zXh<�Q�}I�Cj�:�݇�^���ޭ��y�@�w~���U�Kr�5AP��ܪ��2�x1����Q�쎮<(d$��k�St��I�����W!��!GR�_Dj �U��5L����/�w�lг��fĸ?���S�8�:�<��DV"L���U�@,,N;e%i�#Zr��`��������y�T�Lߥ�Bd� ا�ԭ����5�_|� �>�^!�\R��CK���:�����Xw����͓��;��Q��+~�1���]�+���U�2�2�[1X9G�q�J�%��%��!�l����³���ˋ�i3�ӈS�h>n���OW��l��rld��*J�E���f����n�9VJ���/ty�4�_A������1���U.�8�_ʧ�;4�@!F�H�VS�����Bc���J�&���F�0��y��QW��<S�	tg�_캫G�-�"I*��,ǒh��)��?��K�1�m+Zz����Z9�w��&A���v���}$��v���u�u��jI�����������tm)�;�Yu�˘��&�
#d�gCo�>�r�#�O�mb��\5i����Z'�����L*��W����;w�N�whCG-�r���$],T��^��ʇ\<}�����TW�m�7B�H?�WO&,+��B=�.�p۟����dg�L�>g�h�nq"� 4�ӳN��2V}1��;0�M�j��B��6����oL��lXiŷ|�'��t��lr=I [��1$%����q�W�KR�u�R1׫��iwҀ�v���TG�ǵf���%�Xz���ͪ·�":kZ�p֋�VK����JɻJG>dJ�J��K��3&�f%���;�$��?�"�.27�zB�R�.Mm7c�i*����>����M�� �U?X#q4�4�+��>:pه�u�9;�ƂQ�\����L����:5��VrV��(�����'�^E����q���i+Dz�Z{y5�ƩU�� �N[c�u6RD����}�H	tIAD���kkn �#$������7��{�7 \C��)b���$���e�Y�3Z������l'
a�CƊ�¦d�70�΄6��F����Շ6Ar�|sʲ������$�K�Cҡ�`�黜�uᚃ���1sn�`}���x�3�h�B<��r��)��ظPkA�b���|�3~���Oz@�T��8!�Y5�
푹������ ��M�R>1�D��Q9h���s[�>�P�]���YAx��m,+��G�7�^L��M���4�"�_�x2��Z��O鞤%������&}�^����?�k���.�
��_�_B�:��uT��V��[
�g�j-=t�k� �cO|�)�y(��b@�H��a���W�bh��}b90J���NE�QO����HYK#�i�x	-�^xF��":҄tfhY�rE~Q$�T�f?Y��7����\�����%Y�T-�Ū��՗���	�P�%������������J.��A[�è�}�t�qWq3z���Wأ�
̈��vH"��-��:�a7#��0;���2�`l���hZ8��z��T��ќK-�k��$Ϙ�)1�Q{�*��t���'����(U�!r�vW�=�#	3�IéE�j�ϲ�u�d$��fa���)/�Bi�[nU�m;Oܘ-�T��]��b����d�_���س��҆!�4Sr����g��GW��9L2��V����C��4���_�.�� ��k�+�ﻄ�+�*���j��য]@(��4XL��V���s{@�yi�G6�А��t�ԭ@��- ��}$� uRm��JV��	��)�*�`",��N���ˎY��Ҫ�����N�U!|F��� /�3"ME�^˃y�~M�j֩�Yf�Ɋ�f�-�2[WM����t�����;�8B��/ʃ�Ӛ,?��� =K�������aB`�o��A+�נ]��@�3v�y�\Z��@�o"غb����c
��+�F���h:�,��y��,W���J��=�6��R�vEe(8��@Sb�sӧgS��OĖoܯ*̾@�-�$��f��E]g�j�]�Բ�t՞-��q��ĉ;���p��E[�r{��M���oU �|���I����7@E�!�(<��۬��s����T�Y�Ʒz��W��%ĝ0ܯ����.�=�rY8��̅W�Z�W.�?Kփ)��\�b<�]3�ad�o=t�g�s �ga[c�߸^�G�������wê�ZDK:���VC`��{��縠���}����ؔ������4��pid���
Ia��Y����+�5a��2q��L��pN]��Leu���A�"lY�D$'	�I�����!�+��D\[�x��=���즂C�jY���~�Ǐumqj1�37���H^6?^��Y�g�������$�x��JԷT���������� ��,�t�,|��g��޻��j[�h���:~�R: '�����}@Ŀ�,�f���n�R��b�m�%���" �	�6��L�I.�j	�����a�
pD���%��|�#�N*�/E��C�hu�Q\W=ݏ6�L�2����1
���Z�'�rW�dk�]&�G;�8�������S��l����9�j1;4���(�{Wo�]���U̖��F�Y��q>d�~J HDD�[Kg̛�`���u]���ȏ�L�ۄֆ#r\�����a���Qb7S��g�h������`�&�VS�t�A�e/'D��z���
g���8t�.O�,9�t �XFA�c���*�˖��x���|jo*J����6�'��u�e/aFފ�����L?m�x��6�.~XYT[�[K�&�Hqs����9�6�ģ���WX�ȟp	p����%NC�U,]љ��e�T� ����,#cd�{���x��������ڲ�[���=�˫y��2l̂�h�q��z�>���z1��R�2W|+�m�Ȑ�j����B4RB%8�}��ԥY8e]9"'kd�W��kZE�뿬�s�}OY�:��m<����2r�ƞ�b%̒���B�.�f�Ȍ'�j��t�&��:<��_Ż�p�}z���N��ɵ�9����@`�'IJ��l��x��B�w'6�G�V���#��%���`p?#\��<����K�`�t��z���Q�ӱʆ�����}z`�e`��]��d� y�9hL]��w�<���d�E��$���Mۏ��suc�W߽���	����-�UG�h�'������Uw/
�����xpz�^�+��b֜?��H�ۺg�UP� ��"[`6�0�sƴ���]�V�8���㮼�̊kj��Ԓ(x��՚õlƪ�ta���W�����%��j�Xy��C�$_����p'��*^j-��ɑn~�|�x.��i�'z�%��uU����1���b(���O�1�C�V���B� Y��,�NGIͳ�d�=_�z��3;��q]�#m��[���]���ͫ�o6�'�8�H��q��ծv��e{�d�����}���n2�j#�����d�>KjpR�"B�A��q��b@^�^Hu�\�,Ѓ��^�G٩ނ��^Ҳ�[�&A�Å]O��P�WD��)Lq��GR�1Z}Қ�3=!� ?u��6,_�C\]DS�{����E%��#��]8�?@�ڙ,�).^�=�TS��՗7�>��:���ţ	��Nfkl%�ו��7��~��5�NU���A�$u�b��pA�~9�� C�蘫�W����(ؿz��1vw��JW�����8� &Kn��Kv��dW䓶��k[x��$�.^*��6[�B^	�*�=����N#��d!��Q�?�?�_��_�qZjp�y��wn�U�ah�5���[he�y���Ƽv��^���I�/B�XEc�q+e� ���v�-H0+&3�jj�ƽ�QN2قy�V2N�Z���εP(VQo�[%Mj�y��EQ9���%����*�|q�l�<���i�\*Ih�8D��chk�{�� �=f�Qd�~a�䮛K�.�uJ\�;�Au&�	���p����(r+� rj�������������B�v(��x6�K�1wh3��7Ib�%�i�cgu0�~����]��RK2�I_2�#1�ODY�V����d�Ð}�����.�0!�xYm��)d{��t�E���OU����t���i�b���c�m,=FT��<�p2�]��؈���JiSe%sL9ڜz��5��W=
��q�����L��c��84��إL�2R7�����e,AU+V�+{��{�!<`#�q��}��J/�K�_����nM��F�JV$&^@���nA��%�>�r�"ӑ�B�a�3

�TW
���ߙd��,���Cd-��K�����s'�s����?B�S+
TR���B�F�Ǘ'Bz��Z�~��I�Ŝ�I���2�ɱ{�����S0�� �)�η�����1/�D�|�V���m(m�$�Je���*��v!��� �C
�S���E�L��uH�Wh#^	 B�6��7@l�t/�ֶNݣ[�Ia�Q�r��r�����^2��u8�Qq�<���Q,��gvE�w�4(����7��(K�ىە�8.ҵj�q!H��$?ze���9��]c�ctb��\�1����*��!��S(��R -)�R֫D�ω��8��A��v*)@-�g�XbG�EN����t~��^ܤ�A�Vp�8]�Քy{R���3�2,��o��^㛤�~UP%�-�:]�@v�*��~w��v��J2�8	����3^����E��=]Y��Y�_H��ࢤU�d��ԺL�n���;{9E�'�FX���`���b�W�8JF��,����Ґ��b�����*n�7
"//*�}7~z�E*��Y�2.O��v�c��	u�э��ڐYh�j�ke���ݱRX�B=b�Q9��K��ȿ��0X#+R�Vɡ]9ǘW����߄~�׬���k`ڒW�P#��ݪ`�������Y��U�m�gvo�����..��tC�=�Vy6:X������-6��d��D��.Kqٷv�$���I(�n/�sɨ������9�,ձ���ך�����gX��򷍡OP0��"-�H���.�DjK �HfīJ_p��ڀ���8��>c_t���&��%δ�Űi� ��!e3��50���5�����5u�Ne��n��	��C��#z��V����u������W��ϔ�)�����8�B[?��tC=��կ��%��?)+�c��G�f�;��Z�}\ĭ�6�.^�/�j�#��m��7�ޚ�M��`qU��(]�E�����R�5�瑋��k�؞��ɋ��_g��d�Ar�s��,b�=,�Mk���Pv�%��v1�Ĥ�%�a�AU/�f�V�8S�z�O���s��Y����8x�缭����DsqV81��_c�����M)AD��"m>���y�t��9�K/3�R4_�L+�܃k-�D����vY���I5�t)O������ڲ��R���i
 ��E�F�������i��Jf���bܭ�I������e
���q�݄W}o��-|I�Z7R0üH���I���ϟ SuD��Di`�4��l[�%�$��n��zg��.$�J ����p3n#0S�sv}\��\]��4��\��A�'m_�X%�.����@��,�cs��@m�vg��aQC�r�4\���+1t�Jm��D5̃\<�S&ﳧҷ���ƀ�$�nG���/�9��^������I[u*i��EaMR)Aҁ�y�jx������^�����~��a�����k�-�?G�Æ9��n�q��)�>��/P8���zI��.].��W�Z0ݠ����ֱ�a�Frs`U�9B��ȫA��I*�p_K��c6��{�(����c������&8�}��T�������M��Mⲩ��f��7*�\V�V�bYZ��~C�r�۳�9\�D�럅O_�㄁=� ��ga��#�b�(Z���Y`c��[�1D��Gu���i�@�ƎiJ���1Ϙ���{[��E�wo�8T�Z�<�����.�B�J�5c�Կo�H�eR����|9��.��h<D�_���6Z����궬�:�fG��B��D�aܭ��0�sk=�i}���&�1��aJ��+vc˥I���K��Wg��!'��� #,��p%!�g��\/�����(�Y&�E�L?���途�W�Ɗ��<�H���6��Хm���a L)��*�0;�%䯞��ﹷ�H���?H����MP�%��$��� Q:Pԙ���hQ_*W�O���ۮ�6�U��3�r��ݏ]�l������ܷI���D��E��+p�'.|����MU���7��ھ���Xy;V�h�s��}`����հ�^a8�N�d��l�G���A���y�" �q ��I#-�w���p�p2������T�jG��%粙t~�Y�j̡S�K�W��7@M�Ɂ�f�F��\���&e��@b��e4֗:_l���"��F��CYq����u�<%F�O\���e�ۈ�����:`P�~���+Bm ��E�x�	wt����Xf^�%�"9�ֵ�>�6�t�7̳x����"$lj�#�b���=�f=Lg�zo�����%=��,�?r����@vz��$�T(ђ9��HZ���l�$r�O�ItǶ�XWO��i>յ/Y�5»�C�_�A�a��s�G��xF��S� ��㕮��\4l�M�[b�ׂ#�`����76�'�@�v�]�+V�u���s������U�PZ{&��z�2��W��3b#٦!�Ez�7��v�$�g&�z�+^�y�)�ңn�ʼ�>J�8]�B��:�ҳ˜�~��$1��hͲD�!�����UK��`��(9������T����rk��d{<"��#�࢏�p%�p�ԧ�5 ���x�xeB��	=�_~2�R���`����X4;id��Q�#��H�
y�6��|1i��_#��/
���\qt�ֽ�����#�U���Z�(�
]9����"5��פ�K|��!"�[�w�ըx�{�ɫ��hM�%ǎQ�n�-�T��V?s����"��'*|p@���8�AP���֋�&�	���G���I߼Q�fz��`z⻨��׈��k�dl�K��s|I�sǏ�������é��e���Z��鍭ŃG!2�{f�N�$�y����h o�
��\�Y�����٫9R	D����0�#9�
�aH��@�n֥��,NʹQaS�Ej�D�×GZ�p����H�w:��z���k�M�et5��}�!����F�ݜ�].dU'N�U�W��[tt3����`����SF�秪e����^�,�����M����$�O�*���+��6��S�T�����LK���9�{���+��2�z�[!4u�+��)ޑ¸�����&(�	��u�a<4>�e�Ϡm�ɔ�-=K�fu҃�Վ|�&���`�T/���O�W�:\q>{jZ�؉�nL�[�"���
�_�����µ�ړ/Ǔ|=����ڧ��L��W�	7��P�N9�DE�l�z�J��!���Gʠ�=h������)ةQZ��MUS�jv]�֕��}t�t��!1��71!f!ó�d%�n�4��I+�>DDDb���F� ���7���Y�º7B�}b{�k�l7e��\�%��x�}��o������K��%A�w���4�uR�ŷ�}4�H�:I�J����"���0��U�i[��B�Ȳ�
�~m�jn�M�1����̊�!G}���ˡv�{)�|	�K��%Q<�*���Bu�o
s����D7O�=�E_v�[�`��O�^z�j7~�_�h�x�J9�ѭ���Y��`WC��Z�lwպ��0����㐰��$jM�R��|��`:��{D&��@�w��A�,B@E����Օ�xM�3ƃ��k��5�p�(���?�v�9�нUěC9�ؙ��tb��M����>`�@v1�d��7=d���k-Te�������@�$ftZ��Ի$ǈ�$�{�q�p�6���>ס'�5̶���}�4$(��h���M�ݣຏ�Fo]#���"� �Z ʚ�w4!eC�n�Ny`m B���U ��p�9P^ƒ�g�M�tE��ٳ�9϶k�X��n�T��9��@��ܶ�����^�0�P��Q�M���|F>�Z���� %.Z��9��qa��{���;ٶ�7�DSll�v:��t4�N���k�j&�=#��½J��6��P��є�lIvb���:M���KE�K��/�(�؊҄y~������O=��G�����V?��<�7�� 3M�N���^�+ٮy�ݵ�� �Fq��nmL�Y�輽�p-1�+��<��WѶ�P�F�o�T��9���o�Ҕ��B؛ӰR�7�a98f=6�q{?-�����\�V�ZeLN���Id.gF�1*WJ��x%���3�^|�~���-�f��W!<�3��x�8i���h��>j������*��=��Ea�f�ι
�R�w�����/
������vJ�t:�Y�v����ۚ���4�F�|h��ģ���FJ!$�L��˾�Q�6i���F��j��S��Y��rvA��S2�G���όܥɔ�v��]z������o�tb 3+
��ǡ��;$�z�U���.�V��K]�$Jӻ�>�Z	���IQ�@��v��Y�+�X�{5j�t�S:�Y�ںQ,ٕ_���B4VA/)m"&�i[�rJa����d���� ����]���h����b�l1�ny?fq�J��޴_�]䴻/i���"�-�t ԖC�A$���{ErB�*.l�3/��d�sv�����B����z)=7��+�]�<�Ґӿ�^D�h�L���҆��p<�Y���o���O*����77B���8V�XGBY���X� ^�ퟟUk�E�Rl�� 4�R������OTH7��Zv�I-��/�֫�G�����?�$�A^ʞ��wJ�A�B؄Ba^���F#^�I��MB-����U�.;I*�*�"S7��Y�v����31c�&#�yB�����[h;��
��N�����\�h�F�����g��j���ȘsR�H�'�O�B�ޚ`�J���n.��Ϡ���,�~�*���N),-1��c��9��������~B�;?ӹiŗ������4q)���[�o#^r+|��C�pV��.]��jg�Sm(��?A�'?�B���e�������q�m^�xu��:e���k�C} 4��aMGO�b�]��Cƃq�CF-�믽��y��(s�F����;i�#̀hY�2�?���_�A��^�;����j����l	.B�
w)<��]www�[�����

�@�P�s���}q��t_̟����b�%�Q�eӞ;�'q��+�_B�Ē�Q�\>�0��o3��{����|���|�.`x�N^������S�V]����<��R��������	
�`dqe��<O�i �dOSVV���!v�
@A���)HZ�8��B?�T�zY
�$P%�m�)k
���ӂ��lx�	eT�M(r�g�n�5ﾯ��|���'��%C��y�Σ�`����ے�ړ����OB�j�]6^*+��d�a9�VU]h�`��-Nv-�e���C%��Z1�2 T���sQ�ٱ�z��k[� ��`��6x.r�V���<����3��.G��S��(�)	>O�.�������s���Wן�o��;��>}!)�I����F�r��A�HC|����&��G����`�|����w�J�̱�V����Ĺ3�X��&�x=�e�igÛ��#a<(�Y�����������H��=�C�\���8�����3KoC��N����(m��	��&_Ȳ�V6u^E=ۄH�dj�T�}��Q��1�+���,6�d�'�1�e����]����0����LiX�> i	Qv�Z	��%sbq�¾ɮW{Z��>qo$8ْ��f{)dA"'���ϽD}�3���7t��߯4����Qӯ�/�^�겋��D;��pf��2���SE�a�����bV�\��(DV߸\O���B'6Z)���-����u�P��_U�yeL�d���5I�q�#r<DQ�'��^�`�=���������@GB���:�$FC�T7���b�1W.�4F�)'Z�	����沧N�*T��Ó��7��py�L�ԭ(�����8��-8N�N��.�GU�瞿���M���>j�]6�������*��y�����Y={�˸S��_"T=֛��i�K����/@6&�>�v�!}��L/|퐬���Y�qq�H�4 �f=
�9.S�� �q�nH�ޔn�ԟn���=Ŏ�������-J[+_�v�A�����}�R~�'����|��gUnhn~H���i��MgF5S��vVK-HT��m�<i�ހ��۬�,e}.�:7��OM�H��MF��h󉨓����яٻG��/)���P�=�z8�%�V��*��MCFU��ed?-�5�k9��.e\��E��#ΰ��(߹N@(���E���o��[.�ڽ>̍��ց���Z{Y��:��s���5��r�EK���R�|9����}�A� ���BXe�m&Ξ�?N�б�U�ܸ�4�/�N�h���d���b1�xQ�c7*�6.6�̽�q�e� �^�z�PX��*a5�|�J@�:����W�g�h���R!ƻ�X�>>�U?��G?�K����[-�n'�J��1�`�m.���w�;�H����g0�֡��5��M]hsMZ �֔��ju���ah���������k�<+b�=�jq�� �X �k���<4�M�����-�pa�/+4�u)O����K��X�)9a�6� `�$+���~On��RI��N[Ɉ��"���+�gq3y��r%�S`+�����zD�E�a�y�Y�t���C�S� ̽}i�q���֤�Y��ϫU�3���fD-�*�Ga��Ɏ�����ڔ���Mm���y�
BZs�ȣiu:S������^X�E @Gh(S MUȏb���6��'��8B���3������O�Z�';%e�z�������.�V�)�o��>>��4����D����s�҂��b֞�}9�>�u#���ե\�������|�'_1U(���D�t1�n�]� ^�s�d)�����p'�L9�Ad�r��L�q���P���9�O���~y�P�c���b��?���M�j�.������i�m��D���[\o�2- �$�[��L����|�Z)�ӥ�r�qTh�f$d<s''�{�Pj�IqvwR�A�Ƞ��7v����2�@�ջB������c~��Ui&�j��6�͝�h��P�@*�U����E���T"�V�4�y���z�vư~��==�(����i���a$-��G{�on�Y������)�n��G<�0�6
` ��Q�۔տÿ�$��U.%/��e��e��fv�7.d�'����"W)3?=-%���A����Մ�<�Y�#4��,�ZlZ=�	��Ϡm]�z�]A�B������}�1�<Yg͜��"A�!�SE��2�����m�(��'.��G�Lމ��?�͍��KC^ɠ�'��07��%�]�G�F��<��|�{�L��TSu'�������`#�������1˾ZY�&8In0�r�V������^�O�+�`�!���|� c���岄b���撃2&\�6��xe�S�?)y.5�$ZS�-�E&�ǅ,"��#�0�}��X�v<	���뎰To��7Ga��j��[EX���"�2��'�[�S��A�����X�as#煮,f���v
x��Y��>�Y���\i]��J(�i���.<�,���M�śd����!/N�G�	&�F�D�]y����.�n=Y��� �����.n'��;�k�	6��]&#h���8���X^���/����i����g�>\;�v���,�����_��U�Ř��XpN}bHV������Cvq���m��YIra��9��.'*����[���Ӕٻ;�\�D�(�uޒ�N��?!���P6^{��ynOOc*���6��.�H�uPT�I�d�e	w�m��Br>�X4���ə��k:���b�!v�w8I��$�z�4���.3���j|-Y�2˞�l�_���T����Ae�a��y�/%�~�r��u�v��
�f+`Py�.$�B��a��8i6��<ZLf��hƋ�,[�oe�<����:��//���&`��ڿ�e�+���"�Gɇ�1?�����C�=�K�j"k�,vg'�.k	���q8sWN������I��1V��� ��W�	��W����Ws:��m�{Җ}�9[4�\��y����_[x��C�������ǳ��F^�b�JF�|��3%0^��	 >�j�gB��I�X����dr�^8ka�īxr��E��Z`�y��(�L�ٔUq��Z���Nf�LN���[��#wݐޢ��%�r� ��'����N��.�9�ݩP\��[߈i�q���5p�������%=6�G��W�P�Y��L������勇����:�ߘ���&ˤ�^3�H/��������~�@i�v�y���$n��_�����6ǎ��Nb&Q��m;r8:�5�<�����>"v�\���_t�tT]q/��E[匀��q��5-K�c�Y�c�ㅙnRi�4�y����Y�s�;	>N��}�"��j�Lk�紴�QRm�3�}�ݳ�@��D��{z�G�V���Z׺x]Yv#���3�?&�n�*�\y'������vn����l����D�Q�9͊O������4�2���q��\�٩�j�+Q��F@�Y��������iL��C�}��
�f}�*�5�'��?�=đ�F���������jW��������f����~�t�2��K�������4)�gE����r]��k.��BAwS$�nr�S��s �e�o����u�/��pq?�+G;�&wv�����d�֨F>l���P�VV�S�6�؞��Gx�>��Hxּ�^err�'���lq/�����Y������I�X���he�e|��	�o�|}Z���� %j�����G`����ix���;�J\;��x�+�x�t��-���-����51V�j=�/���g���xo�G��<�%���9�C%��z��do�<w���0��']	�&M=�g��I��3�T_��X�Mww�*�Q�4�x�/�)ֺ?i�?U�P�_#�=�~Jo��sH�ypM��?�7 ���TMd9�?�2�� ��T=YJ�Bg�5z\���3c�v��=�y��t@�.�ގ�q�K�#��-WP颃���lT���� L�*EQ]x_�}�X04>`׺tEVGWڂ���c�ze�ۤ`IߵM,�8����'���@H�����t*m�^��mɖ�1�t�X� B�n�8���i�j�U�O�����m�Aq����ISH6�H��R߶�����#��OA�9Z��Fl1���b�(�ek3䛂)�c~5U&Ѕ�����~�ȓ�Q����2>��
���EZ䲺;~�����LE��ا�[�Q�̕�@��m-���0^	sH���󢹀+Оyns�Xh21p�B��p��Q�l��h�k��Y���;l���9_��|<x�Z�0t��%3�����|���)4x���q���+#хCzS4���b0D�%��B)?q�ϊ8I.!k��3�����a�WRo_DD�44�J���~E��.^�_�a��c�.l�jT�r֪�F��go�}Xlq$��g-j�-?��l�L g� ��&�Q�>8�|d�*159�y�c*��`��5V�T�ޣp�џ
��]�QB��o���4K���P�J!���q���d��qu�E�wU��N�rw�gI6ޖ�j}U��vvl�~�'��}�J9�����s��C&{�K�H����C��;�١�!�������y}iL�\��6�ī��E�`�1	T��p�h��,g�K�5p�0(����f�њ�M�wh;������+a�
�f��-ĿN�'zr�Q��*X�ˬ�J"1�3r@���ސl���޾��r<�֋:͛�>*��z��@b��v����z"Hom�qW�?$�UGԺ$q�ȱO` B���IY�B��_g�̩��L�1�R��8B �Q�U<�	گXt��8��.�3�<��N���҂�9���IFg\�4�W$Ò���<�����������T�5M�_ʎ�e1Vi�<���o/��y�H��.G�b������]�{`0��k/>�KYM�g��n}�xЪ����"E�{����E'��i�g=��I_���cs�p� u��q�	���%�2?���#� ����ĳ�'.�� 7�b`ǳ������6C��H	�;#���1,��C�(�=(`�w����-�++e1i���%��o�Y?��}���}?_�6�WS�fO��s��#2=^A��J��Ј� e����V�{rI�7�<~���
�����5����]Sm ;�^E=9���;J�5�M�|J�� ��cY`�Ie�C������(0�[Q�wnU����i2r0�	����G"��"�d_���gx�\k˒�*�#c�n�/s�D��#�H���Й>�j��&0'40�����L�aq��=�ץ[�3����[�䅶�q�+j���M��}Np)B�2��c-c�\,�b�F�i.�����-��WH
 >�.,�gQƭ-�	��Qs�Q�GךA�u�f6��$��e��Bm��wC�_~M�\��&��&�Hr�֠>�6�=��޿�:x��N]�mS�z/ҡz&}�i�?�7옷-���4Ys֮m�.�em�1�ś�L$�(Q2>����'�l�00W���\���4�>��,�p�X�\WK�<��w��0����&�z�b0F;;Ӊ�;���(������<�dv���U0&XR��6��;vF	��.��#<[d>&�֕��
.�8���"���̣�︴�u#�>Jr�^NYq�ۆ�"�k�h�v��N����r����~I�h@{��l/���u�򈽁�R
��p��mD}1�+M
K���HRJ���T�H���ڱ�)0�u�݁N�y$t��c��q� 99<1�Mb��3�k�N��NA�Mg���=���G�����G�4%�í�e0K��p�dS��K�5�L����qm�>r�����<��N޲�]`;L'Yq��{���\x@^�vy������pټ�D.U� ��0FM��Q�� },-�˷H_N5#4�}e�I
��]��kKY��k�v�a��|2гD[�/�⧮f?.��F�+�6mت�l�q��G`��F������z4Z��ʊS�Ĉ^n�6�y�uY��Jo�|6A�]��N�����%/e�&�6�R�4�ֈS�8i[���?&$!�Cp�"�${%?#�5Z��?�� ʠ�U�=��&��[���ȇf1#�c��x�M�	��*8��|[ົd���1�<e����#��1��r� Nq��fLH"�ݞK�W?�m��q��bX'�DG��K���}q�J)�e�]�B���oӸu�`�0���Òiӓ`����gHc=�N:��D҈�Q���Uה��Ʉ������x�}�R�-YָU���Aj�C�����rd&$��2�G�o�s�t�;�|�D�a�kG�r���7��,���)��-4nku��<���4n��� K�`R�&�?��䱢���\���U�3�doLB������P��8B��u��$Dl�OS�j�QK�b�[��^��=a��.�]/,$c�!�?���q%�������b�U3���"�=s�
�ԛ�Č������Ѵ�ኸN����iNo��~A.�s�6�C�l�Q���}����\�^g�b�6�=��D�4��U�j�j�vi���\��>��N�����O �+�</�F�?�Dz�}R`7�(.U���R�[���7�����us�eY�9�>��U0A�ϡXP�6�CW=/�8%��@��oqS��_\�|F�k��o��:~{��_0�Z��{����J� ��� �&��'Li/�������F�D�٪�U�,:w���Đ��B��X+�t�lE�=Z�\�=Ь����r�#`B�N7Ӷ����`m�3|�F�V�KB��k°|�� 1�>l�sTl��ڜNm�Ǵ`σ��A�[A����ƙ��Y.���7�����ܰg�l�"�V10×��T��^��+vϷ�o�3'�A�=��I�k�����ք3v�U
n����C�;1QX�0�.����\�H�?�W��$�n�U0�4�˸�:_S��1�5�f���%M��5ճ�x�$�z0��^�H^�7\T�uq�ӻG�5WX{��Nb���6�F�pʗ����A\1\8weO�k ߗDp�%�|`����S.���]݊��:�5�;����X�(����|u#�;�'�%�����G7�$
_2��,�2���l� �R��N���+�c�b���D��sj�5JI5P��k�$�n}�SJ�~��> ~�	
	R��K)Y�^�'wFьN��=�x��O�DD}�����Ig�v'F���q'��W���W�2E9j��-�>h��b�˩�;�葵����1��,�q��}#�.��A.G��.�"�1���^5t�G�a�r.�LE䫨�c��ecz_1� �òe:��}��a������C����$Q��N�b-ϑA��©�q���X�WN�;�cJ���!<:j�°�SNl�t�/�d�p#���;Ș��:"�~w�}��_������AG7��E#^j��82��e��`�h����I���t�*�"��`���P$������߬��a��W�{K?���"�QN3ul �?,3�s�Z�e0�'�������~+1�; �`3�H �n ������мU+����v�V�/��fX����EQ�^4�
��ƅ����T��K�^al}ϛv`:��5�yL�I(v�їt,v������l��8����/�Y^q������j�,�9��vڍÆ����C#'l��gk���/߮�� \�(P<�鋕V�A���~�7�<C��ʛ/rV�`i�ﻠF�c�j���xy|>m�J����e�g����ve�&��G<h�:f�}
�(����y�ׯ����'��4����:\C.6]˨T-Hw��y��-��K��	8�/��g�F�i�q=���.���+B1vn?�w�B�8&I^4�͔�S�c!s^*�`ӓ�5����tSx[Dm}B{uc�춾�P�P�^�Dy������wŮ���%�ӣ'A��φ�:}ϡ�1w�C���*�v�6��9�<#!e*�V*q�7>&r���6�
���qks#֒w�K�
ķC�`�g�O��|_7��Ļ[=��e��y7b�?�=��q�"$L�ߵ��`-0v��q�yARH+�*���ծ4Kső�;䕎1j;��p��7<LQ����(�5FW��*�޹.eb��RXk
@uXp8;�9�7%A^�����1|�;��E����3�s䢄�AЏ�>B��Vq�����]��q^��{���`C�y�\(?��k��j�аz4�(Ҥd� Ƶ��l%C�k�GY��]��H��&"J.��p{�pot^�@{�<�r=�n�a������jV����Ɋt�v�����!�[7�
�iH�;fc ����YV��Q�)����J�������?�iG��6cD�����7�����I:��㋸��X<��w��.P���+/[�Dz�qn=�j�X@�y�	u�LR�r���\��ڮbƯ�K�	�q�Xhw �IV@n�^�I�P��>]�nAi��I���a�t8Q"���SR�1 ��R�̤kaf��~�G.������IFhΰ�K���{��V&EW�%'�&ۼ�K�E(��[��!����G��N�M^<���.�⦵����.��+�7��&�kA�?���4�*�!�v/���i�$���K��v ��Z~|Z���荕�u�e�WU5�B��Qux�5?��+���%��@�VY�VP߱�-�e�ʆ�xR�ȗY�F����+�u$��N!�g�Ⴆj}�����}��5a���<rDyx�����~�k�l> ߴp����\(��Q1��� 0?����}�h���Ω���I6X3Eu_����#Q%�M+�<����\HED�Z?�`r��Y�eJ�2��?�3�Y}hp�߅��D��*X���>>���-XY
�CF�q�X�&l8�|�+i��Q��D��'�/Ŝ+ n��<��C�-��M� u����K�59�2�#��맦����)SF��	�g&�Wt}�I9sj�uV>�Q%[�9�V�3���$T�J��s�^�CXD���%�ڜ_�X7�q�<�N�Ѩ�	�q�]���z�btD]�YJ�zƟ��lna%Uف�� l��)���i]�'�}O�D������`M�lҶ'Q��:A:9���(A��A-�#���!�s{��7�e�����=F��Tؕ#T��u$�6�A�4^�,�=���n89F7�J�N�W�lے����wM���!*��>}����d�&I%z<_��e	N����	..� i���άuG�:!� ���M�tkQ�UjwdK�}��짦��P��F8������~bD"V��\	y����ݳe�Y> R~��A}6�Kr��7�㦗�Wr�s��~:��z�k9���g�;L'���=����a �x)��F$^-��.^�M�p�AP��r Н.����|�=ֳ��e�g-ym�
�ݼ�nK�jO!;��W����?:���ܶO��d��Om7zn�+G3�*k=C��n���y�o��h���{1��v�O�9#���Ô{������-�,hl�ڤ̉��t������M^��ֲrW�Vb�� ��~C*�䤤�qڶ�b|�]��_��%�Vh�Q����5��He,�}"ͤ�v���p%a{����ǣ���-�)J�jSb�*��f���I�z'�	�~w�n�h���b���n���H8���IH�{��R�E�t�ϾJ2U�f1���P��^��i��8� �dR�c�ɇ��z;o����-ǃZU�Cĩ#Dvy��X	��5I�,�/YL������ ˤQ	b\����e���n�%��f~}�\���=΁�S�4�$+�$����Nwz�����#4��o�����!q*�w�Q�B՞܍�1cN�u��־>;F�� p1�[��Ɗ�㳨�Ԅ�K�>�,�@����Z�yEu�~ڥ#� ,��5#���g�;�d�]�Z��"kn�]��`�M�W���SL��������&�)*/683��AG��q�����2�����4uXP����dM��a�O�1�d�4䡕��`���A�`�c����<���w�u��@��W&����/�(
�?��1���'�dQ�,���Y7e�܂ٸ����B�6W�*��6p��L�)v�y�ң�|����2"���g�\춽y��ܛ�N)�7�{):��i�nϣ*���h�K+T�,����~E��B�qA@L�:_Z�Tޛ8NbJj�}���>j�/�P��`m�i�&}q�(3�mc�<p��!s�F�s�+3�m�����\]f=9:�"��$�Ml�;�]�b��>��o4e���J����tZ�i6P�"�`���H��Zʹ��5�a/�U���W���3�bL�@��4�d}oJɋ��?&��M�õ�C����t��'x~��, ��r'v�Ab�'������1��^!m�ow�4e����Oa�JK,���I��-��	��1�>�ں΅�J��%&#�Y�}�0V1`����(��DV�Р����� 	;��!�FO~���S���~��֍y�X,��&�+#Dt�I_����g����s�Iĝ��(*�"��B��ٲ��|ù�}�2̟ ۠�sKX1t@�����џR�az(�8
�O���sS�`��ߜ�{0k�6D��5�ev�i��[6̎��RX�tڍI�pmͪ�C�Kbb�Ə@gv9�IA��m�����"F�~mw���֏�=mW'���>Z
L|���I� ���o��b�
^r�6}m��3����C!�ӡ�<�Դ���>H9G$/T��JDJ-�뚣�a�_�0�d� ����7 �u޻�����u��"c|��R�R�~���S��دh��_׃4�
�l���l>&@�;���H}�<�R _��-r�2M��3����8-�@���F����܋�la�u
���y��7��j�t����*5���*�����?_��է'���;�bW�a�2^�^�i��C뙢�"�n'�έPOq4.�c|��<AB8A�K`�; *��ty�s[����ٹ����\ ��3�ܨ`��Q��3t�C��F�I{�.�������Nh4��������g�W���F���]r�Ps�����]�EPl������d?t����yv����[~�J���s�Y�Y�����ʱ�D� �X�-/j�|���I�T��{�v����<~\r�s b;K�N� ���a#�)re�>��Dlghx��i�V�`\����m�<*��x5��$;��)���7Kx����h�]	��ᑥ��l,i�Ȕ�@��e��gӎ�d�<�0Z���iM
�TP�Eg���Fa q��:�62�4��v	��RA<��4��.N&ަ�����|��-1�P��Ix��>��V��K�Pƛn����}�H�/N�'{���鍭&#Xݡ��F���7�u8��vC��8�mWW��I[�P�ݩ|�0(���`ӭ�sjD��E�����X�������]-��=}o ��H�ݻ]Î1��a�����{�=����yȎ���n��{q5 2�ep!���"�f�Ч/�ҙDR3C��=�E����W�.Ŷ����䘒�ˣ�e�j�Ͽd�G���tc}�G$��5�����_�L_���,(A##�����	�a�:W�GC��}�^�;���pi�d���>��hLp�*�&�1�2���{��g��f{���,ݔ��K*�:5��V�"&���	���{�����+<=q����t�R����r��";ͺ����A}���Є�3g�|��X_6�arQ�|%��-Ϥ?��L^H�ȐcA��=l��9����sCF���R N��,�WՉ)Cy�A%��=��}��(��#��&�]{���y� W��o�(
��	�=�ޚ��h�?���xƾR�캏����� n��^X��i��T�����G�g�I	��O�9I���~�AU1����� ���qo���P.�s�X����A�M�� "�Г�����@��Ղ��=�f�5���c�+<I��� Pz���G��&t���&�]�����kaw�m�:/w�̀M 9HM�^[K$��;'�5Յ�o&|�k�Y���=M��P��O�#��;�mըl�b�
c�6ȟ�3e'�eSfo�X���}�p{��-c�%%����'������$�!�<{�Cۏ�ٔSv��mIx� � �g�u�KN�4�r���-�Y{#��Z�ᑨ�+C�F^��u�!s8�Q����q< E.H�cK��n#��uY�#�߹�G���"���O��
I�MV�����X�a��x�1��|�kC��6�w�͚��+	e��P�D���]}(4��3��o���k�'��n{��N5ÃK�$'-�ݗ�a���D�Y�ԑ������y�jH4XWm*X�����=��@��s�M�C��`�Ue�`�i�mI�Tu]��CDAk�KA���1�,�K���ސ���RQO3�臎aңg6��zڛJ�r�cF�ş�5q	y`�?ߐ!�:�4#�鱝������P��q�G�z��Ɨ9!	?(3����Q����sH9a��9��y����)yEs^�%+T�\��*�9ѯj�n���)��:�̯��v7��!	��[0	X�;p����FK�m���Me��֕y�
n�c#��]�r` 1�W�+�|�R�,2���G_���ƫ6���N��jJ��F ��W���`�q���%�V��pɓ*4&��n���'$�Wb>hi�=Pm�P1�T6��;��g��G�8L���{�w��..&�PvV��_�Z���ކ�Sp��Y�>d�0�o� ����,�P���A7o��H��u��~	 8��o���T����gA��/�Z��?���҃�8�%����� �~{0�_%�|�Ƚ#�\��<�Oo5w�C~��(d6���G�� ,P�߳71ŴI���7����7u��� v��YNߥDс����QXB��Y���z�H���I [��m[>u +UL�e�]��c>��i��X!S7�Ym�T�uo�<��~
�Ђ�aJ��<�s3�t��Բ,Z�{��iF��j��Ěi�y9蚻x=,��Eu��W{Z�$�G�F�g�����aNB�����`Ѷ��=N2���%�( �U��Fj���>|��<���F�'��|��@=�O�*�b��N�=PD�~���}��%o�vK� ��-~ĩ�S���qR�Y�m���l�-���:�Z-�����%���N��.'��n�?��4%��Q���7��'��Z[������+��T!�8�!�DN��{g�[�or�\S��5Ikk|q[�Ƚp�&U�ޯB�wz%(��cUྭ�?PK   Jm�Xl� t� /   images/700d3a7f-db95-4bf3-ad80-33d56978804d.png�cs%��=�vvv̉�db�N&�mL��Ɏm۶mO4����?�K</ΪZ�ww����^��+JI�'2·oߐ���U�}���/�� �[�����o������.����9����˷o(���#�f߾}}I���yf�w���8Q�%nl�Xx,3/�}���-�
���\̒R�w��z���|?)�?!�=)\�����a'�� �m�����f3r�u!�V3Yyy��IXe��n ���������;r4Rj�?(�Q�N�H��I!��
��'������!���EP��a���+�̘	O�c�T�G~@�
���.,��폾͍3��?��{L�,M���tq�3}� YC�y��*�t�zm�%��W|�￘�����]R�pA��^p��9�V��i��\;TQ)��߹����{�U��jr�D(����{�I���$*�ײ��p����_kA���ƀC���ܠ�(��%�p���[}�s��H��a@����8�k����KÛd�x;���^"eg���4��"����S�h�H��p�Հ�B��^׺�������� �_��������k	�o�I�D���t�r�;�\�xm�Q�fiz�Q`�:i��_�4E#�A��Atݓ6I�3`�:$�C�����WZ���FV_��s��?p~�	�g�L0�>��ucVVV4ir<��u����)����v#"&x��`x.�gC�H	���U�<��C�I�<�ֳꎂ9��2&�h@E�uC��UT����ZiIyƖ�϶V��B`�(;"�Q �3l#LH��3f�bF��~��M[Y�`��U7�a�����m�8��(����m..?7�F�3��q���DO�8*C��B �k���N*0Wޙ?���Y4p�N7d2G�u�C[�n&#������\����)}�������;titm������6�0�TG�|��ڄ`��|��V�p��KZ�w~������X���o9�h��_S��I-տ k��fA~J��M���l��y>�R2��=4X���~�D&`��<G��a�`'.	p��|�+�((^�7��A��gW��r�˰�	����c�M{�e��v�0D�������֙�8�1�b�_v�1�-`��������D@w�6z;(3��S��\�c%C������	��g����p{��T�y���`3�ģX�ƎŕM;g���`v�ޭ��;�&����#t�zJ{���f�� �os���Щ�Y!��(��6�k͋��I��rm��F���,Ґ������8���slDV��7��(kð��.���A4n�cֶ�¡�$ݯ��.�3]:h0"����_JN�;��I���jC$0��l`���^����mm���c���[Y&�WQ��@L����N�qT0���*t���@�4�<^��Q��e ����[P�Oy�p���5pSm��D^�tc�Af,MƐ�Q~�������$��G�]} ��P����3@a�g�g ��KԴ�>m�Z�C���yH�?t`G�)�u���fj���<��WL��{L�K���ݢ�X��LpqR�ہ	[Y8ӫ�R�@���7d$殛1�I�b>J^���r�U�"�����(��F�l�(��:��fQE��Ѱ	��m� ̝��-N3	{=�o�\;<޷�4�9� شe��;�`�
�[A��3f�r���� �G��$2�oh��57�� �a��5`i�ɺ2���\f��v�$���O���YA�Je�r����#�d�R-m�w?	4a��t��ϒB�>![�E{�!}s���xC{��L!��%;�q+~iI3�1���b�=\J��y�z�m'r3�f�ukO��R���Ѳ�7�ueeZf\�td����}a�&|g��zz���E���:������,�^c��<AkrC�g�،�m����q�<�Ĝ�"]�F-,�0�E���r��QWϦɮ���Пq9�PT�A%<u�cf�;��Wba������05㓾�y�)y�s+��Z�pMF�j�T��ȃ�s�F�Ws6єܓek�:U0=X1C����*��=����F7qR�?#R$Ђ�l+�']�7���3>�8�]"�E/��l�����S�f�(ǛG�����9Hi�����˘�qf��*`��/>��xh>���i�i�Z�wT'�}�c�5b.���Jl�gkb�����\�D~S���2���*�[����-�p�Y��8x�G7v�Ik���V�o�qv����L�`�Jx���˿��)�!�����^^K*�bD��/N�o��A�"��p���g��ׯ�8�����A��N�e�����,Q)��V؊����a�����RLxGq� ��ҏr��AR0N�N���p�ѝB�7ivB�k��z�H�wRf���`S�ׯ�]�ݥ�C[W�J�on�aSyR]8�d,èc�ʅEf��Y=����l5u�^�FA�?SP�Q}t"�T�HC���G%�n5��Mz��-0�ݜ�eج�u�.	ԃ�VK��ً�rn��u��B������.��Ah���c;qUd�����p1�
�*���d��0�tO>P��|�w%Q��c���]5!�M�JW��}�%�횱�n�Ø�6Z�9jBI�\:�0e� �x���L2��YG�Z��/�����A�9�i>��eO����Npy�)k�f̓ah5���`�ߪV).
v��5
N�8��w/{���nҘ��>#�e3y��$5Qq���%ݲ?����Ǣ8�QV��k�f�4g��s��aIp{C��+�f��>���2���;�:ѹ�����1��� ��Zg0Wm\J�u�r���+Yѻ�r9�����R|oP"!�R���i���7+k���9�\	�j�a!�)����[�F��#����U=��:��H�d,?N�jĨN�����	�����]gkv*�H,':Ř���	�Oµ#P���0�*�����d�UE:`��{�k1�6WwZ��>�ܑrԈY��	��k��D�ȕ��6L��<�M��a5���������C�ٓov�%C��l8&UI~JM-x����hqn���g��sͳ�EA9:ɔ^��d;�	 >�	��LI�]e��,�/��RZz����K�0s��K���t#�~D-���HVs3q}ލ �n<�� A�K���c�T(Q�� ����iB�@Y��(�NíT�^_S.�?������Y�,W��|٘��n]�s���o�&CC
�NO}��;��(v:��Z>>�HQ��F%����m7]�>�p~����?�z<E��L=�k�^���p8�8è2J�<fu-�*�q��t�H��P��/`c�Ű%�U�����`���+��ǚ)��j�4O�xzĬ�+z���T�����S{����i�\1>�=vi �Bw���І�+ �b�1���Bc��{�*
�+a�C�Ns%A�#U�
�)Yi��o�+�tm�ЬǮ�u4��e�K� ���o��m�$Lq�lB�C�k�������t�<�1��9��Θ��O�E�悌�~3KLR�`�5 �l�{8��w�ޞ�lkm>�"�i�Y�}�Tî��	��8��<q�!/R/|���d\Z��,)���1O��},�����f�����B�.�4�*�F��2��!��`Uv���Q�\BK��y�c�I$�0�@#B���V��7L-�n�fy���I�?b��1m3�o��w|ȗ�Hע�9���V�%7=3s��n��c?�à�ט�1���r��ͣs�X"X��a%���*�i�,���F�)Y�2�F�:��`�Y��tr��&N�޹W���J�d�meܬ���p�ٕ��('�C�=[H�2>a�u�ڬ�"��\���G��\ȕ4P��ҜI��N �VSqg~2΄tȂ�&Gm�Ĩ��v�[�t�����`��h����J�ڔ{��fz�BH�ou���x%�<ǯatt�|5ve���l������B�����Tr�b��O�� �{Ģ�_��%�zi��-R�����Æ(��,à�NōB�����\J����xnҎ#r�z�e����)�V��o'\�#�S[YʰN!]�f0�ԗ���?��ǤC9yۢ� �9I2BQ��R�6���c��.a�r5q��I�m�p�h�=�����d$^s�>QW/��2�5l?���
�,�<w`�����ӺP)��7������s�C�&]�����c�#+]"� _��`$[D�է�`#�6����_tT\�W�!a����k�~���g��]}�e����/��I���RP~�o*�����D���<�Դz���^�YE
��;V{�ZGx	7��KBN� 0��5&�Js�f�6o�8�}�f��N ne5!��N9�2�/]?�:���O�9���V)�'Up�M�|LD4�����l}�Uj��Ǖ�~A�����|j���<�Q��/1�Z��!���Y�B�y�E䡞�݄sw�˚����<�wa�ؿ����e�q�;�/BtD<[�l)/��z�mY�D3�����a�0��T��@l��,3��}��}JQ;vXkC�-E��W���:�j�g����E?, )����ͫ0���_�q>���7Yh�yM�����ONY����@ǌ5�ELW�L��S�Ыo4���%���sBd4��UjTl4�e��[ɎL��i�p@%���ԫV�c�6��CM���N2i�ta���L�tǲ�:���F�&�'�=)9I�_NfŀH����7��y�>#a����H$�}�Y��;��ǘd����dȐ�?.>�����-�,�d�&*�?ʜ�-m�m0ؒ-���t��!/􉹇ڄv�C���ELvk�$�vM��Q"�2a e��2W�n2i̠"_l6�"B3Żz��L��-k��q�iҩ�@�Nb7P#qc��]{+��2#�P�%w|v�܋���'l�8ԩ�A�/�
>�Up�t�%M��MP�m8�y�X���0&�8���!Х�Ƒ{��\���V�I.�������GJA]����=���x��Hv��v���m������2,�^���Z�ǈ�����xYP�M�t��J�_���I�٫7gc]��������.dh>H�U��F�wϴ�C���A��C���-�?f�u���H�<c�x��}����E�#z�ȱ���Y�i|۰�)���9��ApMYE��f���N*��_r�a
e&<_��#|>;��n��x�9~����2����WMI=��v\�<H?>��=��u)�H�UW꺙����L�*��R6Q�!�w�N���k�rU0���ip�X�JJ��.7!�s'^�m}ޖ�[���h�>_t�pN*Ć��cԡ�F�mr#]��ʨ�1XL�@�;*���[�G�s W��s#��Fѿ��gh���0|���I�ta��K�]��6׃ej*.zJΔ��
Y�����Ke�U�y.G��%��^�a�5(:m�	��q�<���X�D&��ђ��)/c0c�q�<�Xc�X���,�,�'9Ԣ��*�; �� ��	#uuo��_�Y����`b��?�_!��0�OM ��ﵷ)��\� 3D<�ІB��Q�`�3Wə@E���C}X@G��f�FG�1$<����`A%Jǜ�U3�K @e'' ��n����xtAO&R����F-vR�b$N�eۛ~vS��[O/����ލv �P�)(��e<�ŶZ��
#
q�����T����$T>?Z4���P�pc�YF�Տ�1-@�������b���|p�B`���B㥅��B�81��زCaa�[[[���S��o���l0�ir��rA�8�-��7k�)=p��_�����G�OC;��O���/� UQ��a7����$̌�E7BN}�A7��1L�q��Z��J��߱~Q�����y���,�����-]o׻�ll_�i3�ݞ���;_}lA���������U��:^���Zt2l�,�۰�L��(�y]��p���5~|�,\T+~+���X�?*j��VQ�y��~aY+��Bh��G&YE�yv�Å�`
�V;�X3�<����/��-M�Z���È��LTaw�:�>�����l��V������C`ve	'��N� ]lk�|����L��a�Ko���ݶxu	�I��͗e�|=w]��� ��J�s���w����]���T�6�
 ��PC��>Y�H�����#k���	���T^���H�F���p,���l�� j��Z�v���)�?a�#01�������/�q��K�\]'�s�W��J�����󉃡��E�s���,�_e�=2��0�i���҅C�����3���
<���ک��/�}QQVa��#h����k:p$��ػc5��#6��]�y�خ��u�_��J�hn'�$eڽr�_�$�����&�x�N(:�M��;��D����ˢ� (�;6�C��ËW�Q+1��:��|�o�.zߑ�noP!����i��i��I΁��e�Js�ODD3RV��W�V5��*E]�q��s�!Y����JaR#^g{0$/��ݚ�`J	��Kjq�(�a�zCMW���U�?���ΟM�I�����/�`s��h-�|���f����w�����şBO�O�x�Y��8[Cl������iP�B�U9~�k��hI��AA�Q�t�M�MD������8J��EQ�\�'p�O��N�f�:��$b�N��������M��3 m�ũ"{��N���1�X�����4q?R��H���}��(+�A5��)�6�&�;%�?�B�S}}]])Lz``��O1�/���w`F̊kT�8�x���)�L�~����at�	��e��dÜ8��}�,_Ǻ�}������Xu�����Rw�V9R|\�w��G�������V����O��)�Q�-3)D���d�����Okx�t�x��,�*��0z䦉3��W�b�e/�qc��]�#g��g&N��.���ċ!����y�Ahyc�u�&\6�Ow�GՉg��͋e����������߰����UpW˽���v�"���-.{�1Us|x:�=	q�_b	�X�X�!��!�te���хR=���r'�N��P��?�nj��~=���V��S���!�XU����%ZW� E ��}���zqh:m���t�U����e��|j v�tJ
���Л��d~�;�	�h~�������\!�ӓ���E�"Q���25]A6Nohm���w%��!f?�tϿ�A:K��?���~����	�f��a���:ԩd�̀��L5[���Tx��#�`�����&<�iAD֪��j���'�����Y��P�Jk�}5K�Ŏ�/ޜ��-.f�w䗢�Y�������������o�-*Z���Xh1�J?O��Riq-�l�ϖҋ��k�k��L���YɷA�Рg���r�
��:���N���'�f�3��c".@��M���ch�f@�K�O.�-�!���2V����� �:e}��J�"�]O^[?	��@���nx�{���Mբ>;��+�8���aU���m~�B���*H�$F�C>+���'^��y��{�"��]�`q4�{1u	��y]��@��ьaf���S�S�?���r{�ɣl��]�a�����#^�i%����fŋ�@�5�jM����!!!vףݍ��m���DӶF����p��EC���+��
������:)~�~4�@�F�#���^>��M�>���v����p��Z��Wd#�����Ur^{s�YLEANV�[��F�2�ǭu��Wp�V���j���̖�}�X���\�af^`\�4��f����8v��k[@HO�G��SB�of2�^�M�q1{�a�I�=P�����n�lC���*��O�6
k�]�E'ѷ�*�(�^�>��@��:�d�f�\J�dl/�YE�bHD� �fZq?�]K�l�K��+FHM�M����t:�F�����\t{�BrrvF����p�� ��Y��~3��{{3��X����h��L8�#�G�W���T/z�{ِ�G���qծ���$XR���(���K�ix�g,;��:c�*BK���P$��l�\��%`K�]���3WZ[sm�A��<;̟`un��̲}�������S҄�XdڈT8X�mr}�Ԥ�"��l��ŷ��M2�W�0SA���_���G3�
5�jej�k�K[���6�l�N~)G�$�������Dv�����kz�z<\��>!0��z���Rn���k�GB�wW�n+����'�"�k�L��,Z��2�Fު���e�h+��;�z�{�kʶ�sL5�%L(h�7�ݘ���>��v/U����#!T�6>�'��n[�� 3��;F�2����Í}�6m$Ca$S�Oi��S�<�Q�鎟����'�Fg�,-i�]�Ӗ;,ѽ�zk�G���#���c�cs�[�Vӛ���$ħ�aP5�<kN�Xw?)����ğ;���jO6��.�����NY�&�?���ߔ��Y�m���w��V�hU�Ғ}�?�.W�Śt�C�|��F�In�v�V�v�K�Vi��ݧ�ZH>/=H�A&S��>��R�	����]~�`�V����\/���2%�g�g5!oz���GJ�A��WP#ܾk٫Y\��l��K~P��$�yE.c�}��k���+]�ǹk��9�R�,kT�}��F�fc���3�)	{�1�Vrl�8\��8�gh[Z�zu���8��ң�)tG�f�����5���M<t �%��hM�]�����oJL�2�ɻb���`9L�.%�籍�Vd���/�o2l����~�\z)=�<9y�f+���wP;�)��g�T��C��`��V6���#�P-�-��7��K�g(.�@!`�J���ͪI�Dp�����3��w�*@��@)D�3�UE�.b����s,�����Zx�~ڎ��ӨT�Xi\��Ғ�J�\4o���[Q�Un�S(h�b��.6�	5 �X爻	��5[��Ò����kF�J�Ş-�nLJ�����^�06ds,��&b=Z`�ߛy�I-��$�+��ײ8���m�gE~^�J�77����&�����g�n��+�E�TV�^�w�'tXe�W�^
1�;X�=!$���M#Eoj�`���i����!�s,���KI��F�L�D��7R��M�����z��0V�'���X8�kl)V6�@K�$)�P�'Fi�ke�����y�#���}��=(qf��,f��Ĝ��a"�R]���X�;����� �؏�i��MD���jh�����Ѥ�bF�9�X:����գϓ;íƇp�w���ى�'ȿ����,��s��
��,�Y�%�x��/�|�n����J�u$Q�kQͮ�,7C1)��Z$b�<\\#��K�X����THYz�^I�O��$^'R�)�|����6{Ce����Qܞ��*���?j�?>�����x�X�h�k�$�h� �)��w��b���aہޜ�F��b�%��.��Y��<M{"��2��0lA4=�sy	P�^��;M�'f�T��§;���/��Lٜ/=���!�2a
Su���_3���e��i�Y,�Q��$�Ҍ�	�AIе��r)F��`�Y g��[����u��$,s�����%���LN��쁻��j6&r)�����n��܈�����o�7X*�`�X���)a�����M� 55����j۷h��K�Uj�V����ɵ&On��V=\�062���]b$�y��(2��4���E�%ब��һ�p'rp�\����t��]��h�y���Ύ����t��A����9]6��U8_�X8��ӽg� �*�"^2�G��u�}4��5oaNM*�
���M��r�.�]�~�s\���a�Q�����%FT��gp�To���Y�����c�+�m�~^rfA&\�<_q;�D���D���o��xyO��z��+7	��ʁ���>E�O�^��K�O��Dx�������b&}|<<��ړV\����_���+��>��Y�T!�B<��ҽ)�F����Djc���vP�~��\=}i�g:���Lx ��iQCB�]�"��J�3�93���T��2���ҮK�>�Z���=?��^aa��۩�hTE\�hE��fa��	�,t7�W��<�N�����#��K��h�V��Q��,"~��Mӻ�pÅi�[i��g �
�K�U�<� ��8�Y�z9),;!���T�v��T(34���R��4&.~���mhN@[�8&͛�e���~�������q�u���<��t�D��|[]}��\d��{r��`Z�H�^8[X�%�������5?O�Y"�0 f�V'$�O����vs�����gT+�q�*��F^���/���uϋ_/9B�v6.Ur��of ������k��@z{�S���( Ib� � ���yGwH:�rTܐ�EI1��"ykgˀs�}���أ;KJs� ��at����K@��H��PEO_�˝ˡ��d��5����։�(�ppC�6��m3a�bh��P��c�m���GJ��$�S�=��_؍d���6d�:���4T���E{Ļ�n�Z�;���z�:�_�ڢjҷ��cX�Y��V��72��h�d0.���u�ۻ
��uu4�g�t\�b8��::�=W��h
��J�fO0��	}�y��qi!n��RsRoA���mR�bФϥ	���<�3����@���ܻ���\�������=A�`h��bĹe��bn�P�?�_n+������@����l;�iqϧ�u�u����M�]t��x�z�f 3h�3�)o�219���eF%�| �:@��\_���e���pȞ�ĸX1���
��o�e�;J�0��'5��ڣ�)����3��0�j����An�'5]C�&	����N���f��h4q���c���E��I��D	_��L��v����-"���j����4�5HXC
za"���dU�]��ek�kTHh�������$�\8�3���1�\E�*)�>���W.����T�nϥH���m�J1����6QC�oK����b��c��~FDD�`����[VneI�3K�j��W޿�	{Y�s%L���ɶ����~���,���)W%hE�~p�2`�-I1����������ͺ��3�@�9��O7�V��a�����ŹQ�%�b�%V�}|�ck�����ė�5�>r��{��>��S#W�ys>����ao�
�Q׍v#'_�j�z[��;r�v�����<�zI��f��S�H���7v�7.,a"��J���՟�I�	K�lL���Nc�<�k�K�J՚C&�D�˓,��F2E���?�%���������ڮ�+$���&O��|�;�2��qz�ez��T�����!���hQ!����x��H3~Ҹ��C�����d��b�'}O!�~��;�X�4k�Bn�Ǵ}�.��'��o�ʧ�����c�Yg�f�j�����V{�Km��4E&�����L���$3|���T���w��q��	uW�,��ې�@��8S��xc$���y����Ӡk����«������ˮ�����Ѷ>?�f��ُSD�'��J�=R���Oع�í:Eu���Ncg��Օz��QOM�5�밉�v��<���u
��#��R�����&d��iY��F0�����K���	˯ݲ�GG`�ٯ��،���X�No>���-�(���OL��8��{wK�hȳeqS����CLf��qę��ր�얞�m%��
z�*����b���Ni���w�����GU�l:0�p^�� -��ji��߅�a������V��>�*�\�,R\*c�qyzI�<"[J��-_An�l4U�M�Վ��G�U�I2�fR]S���2V0th~�i���dŏ�K�F�Y����a���tE�f��WH6����l��,��zQ�)@Ed�t7�u���s�P�,Pc��?��� 'D�Q�[P=�@iYS�ZR�m��U�ozP���|��@�=91�PK[\��������ʲ1��z"i��ҍ�<Ne���gAh���g������ǡ�:�����4�,�>�,}^�c�Z6�M4[�p��d&�w�:�
�a���+Ub�(Y�HR&jl�_�pG�GL�?��̛x	�oN�&W�#��OϙR&��I��]���B��XR������%
���XZ �p2���γ�wWOu��>��	k�;�*�
G���)61�<�J�'ާ	+5�ʦu7X�d���>���'?$���ǉ�����,'�`�˕D��U���]����A��_���V Z���r�%����R��xQL�6���U$�\��j2��c�C`�3�v9��+F����:8��kՇ�����k��M�q��#����W���/&�9+ba9v��_� 0:���a�W��f�Ϫ�)���`���\Fz1S�9���쐎D���rK�"=n�+��<+.�)%%�L$�RZb;��!N��:=�I3��A���+�K��uz�P5Վ�Bo�=�{e���;�b �Ƀ��]�zj>(z^�vcR���7����=��j	���1�S3�p[�lG�2�t��]\d�x �#q���>�w�zV��Ân ǀw+�m�@V��Ac��)�o�O���
/ދ��>4��+K_�e��=�=Z� >	T��T������ �m{��H���Y��w�b�aSPV(���o�k�ʔ��<�5���J�:$��XX�v���mH._���Z���/����H�z�qv��X���.:���)O:g�מ�TР9Le��,]�D��O[�T��U��|/����L� ��(r[�y�of�КP1�ֲ�l���l�{�Um�w�����^�y9��鑂�2ǉ��;v�G�I�V,�GW,F7�	(�T��yx�Ғ��L���G�i��]�f�9���t�h>Ԙy���i�F-J��́�����r�+��ӷ��:�V��S�m�LR����A2]�{]��)�Oi�W�ϰ%�L�~�G�DI&�2<9=�M��Fo��� �?*�(y+�d�,g�U4�mddOa�h�V�.߷x��+("H�kR|�̍�YO�kʩ�|�dj������$I�S�a��/�ڵ�c^�T�4#�+:�n�~3�U���c�M��z~U�!��ާ��������&5������/��&�sjo6���wV��M)?�Ω�|��f"����x�הl�tk%�dw^��"P��7B˩ba\�L(�$X�bL��E̸���9�e2NM�79t~�==�Wd��E��<-�a�Ki&�Nkݥby�&�q�f��3���|&6.oA��{�ɻ}1��]����̂,<`q�����%hQ#�=	��蒍�Ֆ�����.;���.{4������V&���=�l���Ant�k�v��)�%��Cm/kY-����'��7.]~[g+��m��o��o(�`��!�i����Y���\���9M���7얕#��������4�O.ۘ����֞]��]���KۜK1��V����e�C������B����S�v�\��Р����$�C*A��	4��K�U�RzX�?�3f��?�����k~�d�t�D�c%��A�c�#�Q���7|ZH]sp;�)&�̦�}f<����Q�������i0�u_|K�s��z�|q9 [�wyt=��th[�"�����(-�����gͱ���~W�J�-��&,��RB�%����Ș��P�ԑ���6�ff緣�����GM6+��B��uP�R���r���	�A��`:�\QM,1D��t������E=������x�%��Q!r�8�v�D�^��-4���e��v���l�p��!�3�qb�������,���k�C���4rwϒ��-�͓�ѣ��	��S�U��E��+>?��WrSf��OJ���#�%%%�G,-���>��?Zv>G��,�MK6��H��Bc%�%�1fbf�}ty�~7�6|��Ha @�����&k���q���6��I��v�o�����t]O�~���.�#�Ņ�%������ګV�����p��p�_���C+9�x�c�muʉ����*�*�h�2[u�L���
�=Uu��⠩�}Kd�!y�d���c��gYC���Hu�Z������m�m�3ycy������-��H�MU�/���h���% Q����RwZF[����=�B���h<�7�H=8o��1��0p�a��N�c���e�7�Mc�<�����Sy��Z9�7&㚑vE:�¶݅C������!�MV>q�4�4iH4O�n��+�Z�nM�[��,j�=+����gqe��j��2��kv������
6����b��q�� X�i�U`�xASf��(QXU;�S_�7B���Ma�q�0d=l'��������{��
6%�ǖ��#Ԋ��#'ɸm�����6<����q�p,uI� �I9R��P����M�v?��*lv��qУ'����*"HH<X{�Wc�[�"������7�a�����Q�5�5"?��B�6���sAo�aG�8���ϣ��n\�R	�{����*�]:�.���Y�b!�a��G�Vh�<�$Z������(���L��Ȓ��C�S]��巖�cآ3V�w
ei&0f�80l0s���oi22�;b[��	Ad�͙�"$71G;�!�u�u���J
����#��W<�O�>�	K�CH�	�,�Ue�#���6���V_U&�w�?�
&�BО!�'������^��:ʚ,3V?l��������#6�nu˫$�4�
/�,?�$0�k�<�OX�;���w&[�)��.��z���䜁��n�����gwE�]���N����5Ӵ{F���<�V��nU�h�|�*�5���13�2�p}ۖ�D�f��×�Ǹ��.m�v����w�-�+�����ы�̇��Iu�������K���5*'�����U2U�c�yy�y��lm����5�{ő�5�ob����z��uУ�Y�}I�/mƌ����<ӎczCZ; *I{S,�d[v��~���v�/��\���t?� �s��)��&r���m�õn}��{e��y�뵠�Fo�z��0&$���R�'O�����˃۔���<g6��d�p�,Vi���b�����R�Hӈ�֗� �����	\�>y"ٸ�N��CUN�1���ޝ�YZ�KK�	�I��(N��r�s�<�DǠ�n���i��e+I�x&�we����~��]x�"NR4�k^�(��W��X��~5�G���ٞF�a_ĝBX'�C�P�(�X��M�c��tft�=A#Y�[�>JAޙ�n�լ��ܵ�,y�ƫ~A��A"�kp�}�p-��}�'� ���J�ty��D9 �Դ8v�y�x�I��y@o���h�#
S�n�k<��8��Iw&������s�KZ�w�)��	���=��Uh�k��nDH���O9�ʴ�!!�z B�`Lm'Ak�����U�� ��i�ڃJ�mѬ0Ge�q[U���\�촗���e" �}��\8{r�>��=��Φgf�>��O��b��dџ}���
���\u��c[�����J���&̘���7AD/:00L.$�т"��ݬ��Qҷ�����٥�e"�`ngUZ�����AnQ((�6m=��@�~>� !�n����	�?�������{X"D# h�Ğ~�� h�&k#��ʿ�Z!f��U�����Ɇ�<�io��ry�S�o+n��[[����6_��W���캝l����ͽ�A�~���#y�;#|q�0𴆩�	V]@��5�We�`o��[�Q�T���q7&t�#>|$��F}H��l���/A��ۅ�������1z��y��z�u��;:�z��Bf��?���0H/WU= UAT�CJ4��rH�7�>�C5`�#i#�����[���@T�X�6�l�1�S��[��u^Y�2��i�ȷ�`F8}ɾ@vfz�6@ׄ^l2���y���Yd���a.�zJ=�Y�W`��J��`Z `��]�o~C���������JJ�|�h^i�7H�,���ߐ��4�F�24��I>2/��/D,��XW�l4�Z�_PI���i�����:"l����
�Л�Yeke۟$2�L��Gj�M��|ZU0�Xk�"�z[1xA��c�?J���$"��NY�T�¨���ˢ��٩SW�v�v�`�r���<\��������__;�� "��g�u{���l�Uu��1څ�=`��Z��Ғ����a&`,��!@޿��%��o[6�~'�%I�툵��R�UE�e�S��Ls4�eW�)d�9�m���� ���;]m�P$5�g��Hhϩg`�Y�
�o��~�P�׶��7�Lρm�ԩSp�P0�X.#"�J��ٰѐd�\*C1��8�Y(�ٌA���=y�ضm�������q�H(��e\H������A>�����ik,�:��3�>s�܅��}va���7���,�M���s�l(H7Bv��;E=T�\% e�ɶ���4����eρ^b[���I�@HL�\��)rd�:61}X�YA�.^��;����{����^��	}+y�M�~%BR"�$��b�4- �G�豰��l(�A�R���eo���Hv�tI9�Ţ/4�����ip$0��=}��mٌ�h��$�eLr��8��,Ot�lY�乘�LKڑ�����!�R*�8y�)���*+`�í��]�ɾT�e)����G�T�m&�f�_^{E�g	�_����l�Rͪ��ܴu{c(ÇU�d1	����%�~�/=n�����~I�nֈEH�g[3)C��|{�,$4km+�K�Hب�\Y&��@n�b�"'1�a�-�@�W�~��`W��	�B�C��K�j:����\�M&�Qd�!�V����ɻ��P#��מf۶U��ki�e$W�r��������EI1���-��hZ+8UK�p�02���Goر'�=wj�\Z0�Z ��fit��o��鷺��7�7����#5#���u��RG"�m�ũT�RQ~ڮ���]O��h<Y�H;�-Lj�U�^l�Sٱk���gF�ED�܂��sY���q�Çn�V+`ߘ��&�RX,*rQ��%D��,�F�e��Tww������` e�s ���kV4z��6�C!#L
d�D%J��g4<,±�1�A�4�l2����J���18�0��4�IE2V�@F���t�/V-������{����v��m�������?���Ӄ��k�m�Z[^��7n9��ŴiX٥]&O�kY�"���i����+���I�JWG;�jӓ�gO�I޴w~.�Z.�ի33�x<���;x`av����G���a��C��A=�cU��)_d�`0��U�3+�D ����Խ{n���̂��Fc��#PÆR@�$uoX�.��$�r.b=$)��Dv>��+��4x��͛6�����!�T�RZA��w��i-#�ԙ kr�fe�g#��ҝɖ4Y��-�gf��	T6�M:ͯ��F	��ZH�����Y���u���'�(�+u��l�"������*ժUs���b��}�r�d����y頣cV~��1M���ĳ�њ�"s��h�FU&�AH�I��E����˧O)���̈N�'�]�=i=��J�b�s#�L�Qqe�4F�����L~F�Hz�H7���ŗNu'�	��4!ȬO`Ct3�L�ö��J� ��҅+@�o}��6`�P�D��8�8�3d�''��`�p�����م�@�H��3�R<j��!���ɳ�%�l&SX����
��㑎� L��Ѷ��cZ��Ŏ��{n:���O^��pkpG��*.H���,�F��áh h�����=q�����`0���E"oHqQ0�bS�ӦC�SaDB�ڶm�k��I���eVI�K�g��s���GA\�,���1v����B�X6?H�v��ێ=�D~�#���N��0$W�u��V2p�@�3I֗�Ɔ�@�M�6�z���s�=��;:;I �����&V��r�UPО$��M�mm =���������e4ўq�x$�ۑJ���v���k�rg�}rt�ȹ�.��Rvj*~��H9:�����|F��@[��U�4cP����Ka\���*��f'_��˕��kєG�vݪYz���ݑL󅙹��م'�}����R��X�\���;���B���*bEv�*�}%�"PsYĊ�#?_P�t��\�p�s�7�a�0����Z�<,*��+*��
#Sm!��C:��-O
�N粅��6
�*�!����l���}��_F��d�^*W��<�������o�5�D0c������T�h�y��H�!0�k;���H�3{u�QV]Z�tdltnn�jVa���]O&��$ΎU�g���n�a��Z����Up���Y'�t$[�ee���G���L��hNho�iiUS5t��H�c#Z9Q�n*0�d����<|��F9����ħ��̹J�k�s�%�A�.g��sm�nu��Uq�=���L(�ҕ��Y��j�������vG/^i�}���� [�0���eǓ��e94}Y���ѓ',�}�/X��G/�T"�Dň�E��b�š�s�v��jO��ܱ6S��DYј!��cy���o��׿�v�z��#�^�j#\�4��A�P*G"�s�� |�]ӿ�b��d�:>2 فDS�̬�DR����֧��֯_ߞJ�&.�:uJ��(ЀQY@6�� ]����f3�xzT�}�X�"�$��d^:�i 	��`$*P�(�=55U(�!�����A�����ܫ�r^H��@�=XEe�z��k��b�2r.���bа\>C*i��$ّV"#c���LǛ�_�A)��`oO�l9B�>���M�Kse5پs��u���sc#;gf&�����Ba�5��7[�R<���~GZ+es�JA���HI-�B��z�e�t�L� �UWR���ۿ����	#޲m���t%�[�C@�F͎xh�4��9?3�{��D70�G�y^?��ly,7��w�b/�'�H����`,k��آ�j�"�V�g%H��$)�W%s��pw"u5.�
�����$a��	��������_�ɔ,/
D�� ����xn�]@���[O���"$
�g�pUi�)0�gKJ�z�@��R}�d��?}�������/<����E�V/jp"|�@�-�S�I?�%�2P�"A�	XE��v��"���J5]#���AOWh��D�J��Ԣ���م�:��Ĩ�U���ˊi�5�P�P$�r�b�kk�'xU�mj��`1l��""��z �Ne���Ҕ����c	�늭��4�B�`
e/S�U*e"N\��,jz��&�1䖊b��;�T�[v<�F��
Ma��m��U�ht`;5k0+�Yͻvf�$h��/�
�L0H�Av���#/=��cpSk��H�p(T���7G�qZcZ$+7�;T*���I�����^ߔ�
x:,I�i�+�DIՍ��+�j%_,�L1�%���@78�Db���`�C��P@�"b���l C�%���偮������}W�j(�1#�� �D(
M�m�P�Do�1��mUeYc�/��?������>0
�K��W�U_9��|fnn�$'�a$"Q�N�ܽyY0s�t2��(T��j5S����;���U*�Ct����皨弣��ѩDP�4	f!_	������.P�,��D���3�:�Kw��Ed�[������R�|��O�ģ`�0���
�uI�ʂS�E��x�%F���D*�Uʊ�]{n6����&�r�`�d�ir�čx�kx{���� ��V�bS�> �+ݠ�:��"��p8\��`�I�9@��
��?w����^�n���vv'H1{\��J�G�J_h����Nlݗ\��l�LHL�1A��U�Y�$���<�.���S�"!�L�&�L�C�������P��z�����B��A������"/Qa�WM����04e���Uv@`4�R�Ĵ"U*�Ј>L�(a|=i��ܡoh���BP�Q��o�(p����{��Q]�╻�:���I3iF9$$�@X r0�`�1�#�g�z�ڻ�a�6ۀ9GDHH	�89��tN������I�x�o������Ck��+�{���=��h>�,��!�B�x�T|�)�b���u��MD�^�p��EL�����&H�$RC%�hk�4���JC�+MG���X�PU.���h$���z*H�#�%;ogp��hx5U����L:����Vu����tmm���ռ��9��H��Y N�����|˭:CuΜY�(����㉄�t7��ʨ��\U���4���43�l������Q��q�B�D�bIBTT��fr�%��U���x�|Y0�f�VXx���g'�Tp_��.&��K�������:t�O$����Ν��.�-8X�QB����^�9j�Rxo��Ib9x���� �vww�?�=��d�ٴ�fG[К������6k����%�J�o��'�p^ziMu^�|������?��V�yV}���۳sG�����\��3�\q�屨+`
Y�������k���_~��S-joo#O��y�̜lMC�@V� Y��V�9-�L���Of�#�`�[!k���J�J���h���t���Kf7� ��#�hxg���r���>N�Tb 2�L�*�5�
�X�&�E�qaA(�(#Ͱ�C���dHf��@K�A�Z�Dx��p��G�sΡ����{�G���φ}x+�Z��v���@iX���{Y�p��3�!ie�{��e,�iɊr465x��8Ƃ_04#I���/�h��T�cy���8�?��*�����;��`�hu�B��-�����7���R�`��۱��N��)��===����6Y���37�Z;L�$�1i�	�,*J���'�Qu"hpWR�lcX��v`�%��H��+����uv���q
.7�y#����3�|R�0Eǐ�$*�w�nq
IR,����*�{ ����q1!K3,#��%�m(�T$�u<	�B��n�RY����/D(�bt�l�����8����c���nh�bXb��3_}�5p</ <zg�V�]hjk�.�K-˂݇y�'>����|s󛛷��#lD: �k��L�T$jpp�/}�k���$�_�h���UUE�Ne�6
g:�cnm�KDbMu�%)^�CUY���E�7�H:V�>}z]]]����m����a���kĹm۶��.]�m, <#�=I�4p+]�9��5nذ�b	7M��s�stlxhp����`�
��[��D]�4�&�+Z++�oON��A��&�JL F�p����{�}����/Z��e���W_yeU�+I��@w}ą�b
?��c���F&~��r�p-�'�􏣆GۧnY!M�m�d���g��E;�.x�N������.���JEi����ٝ�
�S���-J�1�*��4Dվ����@sR�d�X�}ˁ���1U8j-T� >ZM!���ӫ�|߫ol�-\���A}�h� _k)"�vvUm$����?�NI'�h����G�w��V�zmt6>E��x�+��@��i4�ɀ�����J���rx�	|�jJ�wT��V�V)���Z�� m]��������8���Q鱝L��r�Hv\�h�P���(���1��SIZ��l��Y� �JR���U�4;�+�0w�w���b(Ij ���Ț�RQ%��	�I�@'��1�_������B9m�*��(	���87�J��1p�#5Y������� #��]\�A��:n���c$�>�F���e�PU0�fE�w����&�B��6�z9��� �9P�1O�,Ws�ݻoxxxтEK.�hs���rV��S[w��?��:��$��.]
�`thx�޽�WfΞ���WdT��>�#��LV
k��v9]v�#�6<�A���ĕǕӣr$,�Np���1fss���o[�dq�iu-� �By"�
���2�|���y��_��|��Ua�7ۧ����9x�[o�Y[[=cF��hbd$��y��<�C����y������D����sv0��ظ�p�����C1����;z���?��c�+ᡸ"��/f�4NR���BTg��y�{��}����G�pۗ ��,�����mK|�BYH������pM=�bغ��9�I��Fp	%I���A�x$H��Z�;�j��8���?P�CU��w uo�M��Xd$��i�`yƊ
GE؈���!R�x��������ôo���u+p����'+]?��xhQ ��0���hM&ai����v���vu7��5ݪ`�q�짦n#���'-	J�|\(N:�9޷�~�/*M�hx}^�R	�,gC=f%��C�T��k$��FA�l���o�Rp%&w
͊�;6�
��i�Z15U_O�+��VM���-�?����̗r�ӛN_{FMm�O<F���.��l!�y����ϙC���ŝ�����/^������m,�	Wp�.��jh*���&UXѾN��*�#	;�Ќ��&�@�ιBi���I�T�)�
�tΎ��`S���t ����$���D*����d�w[۴����f���ڵ����a���i�QX������
�(�/j�n=A0��p�	��1������8MQ%I����K�6��Ɠ�XJ$�C%1� ��$h@��x#VQ�F�`?t��HJX�� a  ���������Y���|II*������+��ﾳ#�H�}�:��d2}���9sg��|����.�w�wÁ�G��Lk��w�)��Ne׬>�G?�qkk{W�хtuu��F"�_��㩊�=tr�MV�hu�����>x
���#��Ʀ&JG���n�M|�tQ���9���b4~���~h"���22�<�X�����E��IvV�Lpm�p�'4�Y߭�4ʒ�U�.B(XRȲƳ,ò�lR��7<G� ���Q��H�,�/Ê8�q�'!�ɱ�\��S�f�x_Ò�������eI�@/��#�ؒj(�z�*� ��A^&�!������Kٔu�Sp�/��������wQ�u��5부�H�,��}A���Nbi`�OR`�_��'�To��c�t���+�,'��pd3)o�xqW�q0[.���&�`h��A��<oe'�U[���a)}S�U5S�D�V�iLO��f�m��³��t���]�q��/mݱm�֭k�m�v��֜yV{c����1~���t��_�r]]�G?���S� 
*��4o4T�C���*��R׃s?x�Lǵ�<�Sbk��"��8ׯ��z�s��~$�F�67�3���X��J��/(ȪS��K��K,+��_�썟����Α�����~]�X�(�������%���餪�xĤ���8�E_� �-�؃w��nj��lY���D�{X��	 b�1i��SeI�_Q��)��}�Kjrcu��&���5�l�`�H�����5 J<c��c��G��K�r!WM����D��x�A���Q �����9�"��斖W_�D0N��Ga{Sc��hccq��e2�h$�'���!I�R�����Qͼ!k*-�M�u�ز�ўA��,��w���>qvM����̝w�9��cfK$�Y��/���O���d�p2���������8ɬJr��tM�^�	@����<oWu"U����ҙtM,�t�Y%�"�2L�B6W[W�dQ�e���Ŋ@Σ�
ǜ�	�jcD��v��Ȱ8�6��4\�>Iįi:D!�|�B��'j�L�4���x}�����jZ�ɔm���=<�b1/J<�s� �äm!�Q�EpIU�5��Is���W��%K�����������p�/E�3���$���5+j������t�rP���O��s��g�O}�SW_uL�W_�������g�)�"5E��3h�$�񑑚�z��� &u�Pȉ�Ұb5Y���9��)^���Ɩ�>�mQS�/�>/���9k�^6�c4A�Z�v���EU��3f���}���;���?	y�hu8���g�5~}�,Ow��Υ4Ccy��gslst�p�49�ì2�Q�Z0t$��o�f�f��h̾�Q�aF_ڴvU)����՝���x���F���i��D*SR`m#�l��zk�e��:D�:	����9�:�=��/�J�|���%�J������i��V$�9 X3�2#��H��`2��J%�^��-�3��J��o,ae9�I�]��Қ� ���#���&M��d��ɩ�$iN�?2@-�b�����
d�!���n��S��:8��u��X(i��s�ƺ�է�Uȕ39`���WOo|�Y�.��p��m�b����,��n����.��������o۶����}F�?:g��o��v$ٳ�Pum#�gE#lnw }g�{��k�V�`9_��6��c>���yξk��H�i������xTkO�`�4�2p���=�~����fTG�"���O�������]|�ڦ�EQ�2�u�܃e�-��A������������yN���w^غ�����'ō/>_Sv��H|�}��S�P(�@bL�0*��鍚tIF�v����$��Mf��s��C�q&����"k�es-�CLðN����m6��i^7y�9�;:�O�t�;甕M��F��8�!�9ƽpB0�`���G^}�U���_''b~7jVa)�-1u�UA �j�j!�D#�B?� El����biX$���qk�����=�#��n�U��J���v����dca%��Fc�t�b�捆(
.[]>�AHULi�磀��~��E� ���(�</��ȋ:8��vRv�P��rU��s��������S%CuG����=����j��鱪��g�ɦ*�@D��I�IE��u��{;n�X�`X�e$�������;{�~��{5�t{g��n�����}�t����������.8K��=G�=���_�k�=����vy<�U�V=��#�vǷ,�J+x%QI;�"0�I#��|�FH��)�_�v������[j뛧�^p�����-�Y�	����e��%0V��z��}P�Z$���
�܎ې|'�d�嶛�KJ-
r1 Ia���gL�^u���=`��˖G��$)�&��S� ���|Idm�D*�d"��l�RY����T���蘨��:�Ģ����B1�����.���ho�`$�= �"��A����i�n�jJ�-��@G<�D �<��S�۲���vI�g�=��:ƚD]��XS�)r>��W���O�������z�W�h���
�5����O���'�i��X�2��qe2�^T0�岥RyǮ���\�vqC�8Գ��'�yc����܌s7���{�pOס����B"d��̪��e�S˂�?<PA5#8�h4���
���mq
�> ���q��B�fw�	�A`Y�n�%)�D_��;���R�����ֲ�����㴊�Y�?,"�6����]�l�aRTK�|n"�#�l�8ۤ���p�����4U�@M�r8`���].Y)��B�R�$"<9��0�Ͽ`���k�DX	�l��{�\��-������!8���3Q@�'I��mFIQʈ
�a�b2�3cJ/���kS}F�Y!�����.2�B����򢦹팢�&��D����]��U�|��g_�2\N�%�����F���\�P[���QS�p����W��:�~¢��R+��F�w���3|k����sg�[����v\���E��SO<v�ӣ�����[oo.�g�夼k��sϿ���ۻ�����׫�<�^�����(MG)h$i�V�;i�b�w!zu<��"�ݹkw����}}U�5� '�`s�!paŢ�Ɉr����3l;�pq���DEb�O�̘��jh(5���..�;e��i��m�[��r�<�MPr��a�t�͡r&	P̓��G8}�T���m�d��P����
�jbs�w����G56L����q���`yE���/[��c�P(w�g�bռ��eU��k�P�(��v��f9p�.�!�����S�h��i���������g����0֕���W*�}>�����*,,�7��k/BUQe����"�T1�G����8�g��9%���ݱ�=�  ���-p��=�c#�ۚ�9��"�� 2i��vX�Oh�=���'3䆕Z0'W�?~X�����'�/4u�C��"�a���VhC�� D���)���Η�yo猎v�!x�X������zj^{����D%�7h5���a���L&�- ��4H��X��`s|>�\6	�������+�T-�Q��f�XH��9-��*���V����#�P���i�N�s8�����xWWW��I&'lZ���c����555Gz{�gMU8p��Ę|a�}&�A����W-N�c�8F>��봦��oxp)ǰ.b���{�. ^�\p��+�yǼκ�������.�k`"^%�����oo^�jumC��	�u+Y>���=��U�~I�U�gUC�&αP=�EG�zZL�BN)�"?�֖-���@(��g:]D�T*��;\�P(�N��l����b�puu��~�+����Q(��͇�/�H����a`��R�b�{~w�u�DY�皳�UWվ�uۿ���I�sކLF���t�Je��vxM�(1�"�q�lN7�tX�&n:C�!� P� >��q�)3�ˌ��d��U+V*�&������'&꼡�s�{�^Z�vly�eZ���s� ���\b,u��U��V�XG򜤈No W*��#Y�x|��*8[_0P.ʂM ��ϖy;ϻ��`���8}�pX
���w�h�2pD�j�	2Z�YR�M�Q�r�m�l,<����4��g�����	�vhI�����I2Q(� �Kz���z��t���Q^p�m���M�(��%��is��8:�'�y"�N��{n�W ��d�q���5�ؽ{w&�25%���D	�������LF����f(1�p8���qUU��wp��7\b�	�A�9uz���g�w�+�՟���U�5 ��8]V*G�4�����`�c?x�0�a��y=>x�:v~0=P|��7P�/�q�d�	� ���ڐ���ѩq�~��������h?�HW/�Uݲy�֭[PCE"VY�JC�4	k��/Sѣ�HI� ��H��W�4Ȥ��N .D�a&�5 ��93/�j��*�LV�D�*�X�0�Q�ʪU��q�w$�^�t�믿&��e������p�0�rS��ܻw���(�؞�{^yecGg����ۢ�ZU��X����Z�$Q�U���ԒLa8�J��e�.�Y]M�$��d��>(��Po���r:l��iXh���5�W-Y�d߁C���5>�<��=�]���$�k�V��12V�(�����?�sRÁ5/!�M�3�$|{|-�>x����w��w�'������B�n��}��>�-[��u�]�ӧ�t�Mp��L&���˗/gnt,9{΂��B�pg�~���#��iUQ��LKs��j����_���7�t���m#I|���[n����d*����W^�5%���s��+��?���k���l ��Z��g�!�<*���:]*�Nc�N8i��d2�:ԑ�1��3��p	��� TE���1��N�	�H���𑙉�G`cA๚hP`�xB�ݶ���ٗDaz8������|�5ii���@�iO�rA@2�O)����dQe!�d��E�5^.k��C�̌���X�Ɵ�^�y��D"�s`�y�y�-om^���h�������|���F�X��2�H�����S}�M���?ީ����\���z��k#���1��λ2�4�������=��68}p?�w�7j����,a�[퍤fP�Đ�%l��X�w2/<u?��eBS5pwo��vb,/ ��3CEº�Ex�p��K���$*�����LM�7���F}JzUU���%���?8�O���z%�]
�q�ORh�l$��	��fP���2�5�Q��hm#��4�Z捱�8ĉ�
��Y%3$~]��{�H�mvEt�I�����t},��u��9�R�]�XA%�%���V�˿��򦷞��X�������8Ϸ7�����-����������mjߵkg�'�PiY��#q?�o��%�%�flNC�"�
j�ŲG?�S�M2���Ӝ+U"�� F�"O���D�l�2I��mV�u�w~��W��|Z[ۿ~�?֟w~4���|��T y�E��ۿ��L&}�}��4{0��lV�>���lSS�D:�`��yN��@��4;Ǿ�֦�0�T[��u/�����X8R(��~��#G"��(IkW�^*�o߱���hUu]CCS�40j������M7~�_��ϱ��;��qZ6���9�s^u�Uv����/),��gppF����3$��X|�����k�9o<_*j %QTw<����q�{G��>�{����/���` ��o)���LGe#��`�CcuuL��=��cYS{��ZrlbZC���̧R�R���˛k{�^yᥡ��PMՊ5k:O����EqAG��ŋ�
�h��*$D:(o��b�MA��#"q�PH���$\81>�����>b�4��Gx�{��D?_|�܎Y�8r����z��m��\sG��@�T�.�D�i�F��Ñ��2�g���$w������۽����������}gGww�ٟ8{�[�[�M��6&U*�{����v̇����s����}̙��c�����_���* T��9�L�?.�(�����=\n��
^�-�L<���2J��la9�#0:�����n��|H��W��c�i���C��{jP�O�����aqW��#�s�R����ŀσ�qn��M���  j���;|E�����<���:��ӌ͡��(cwBK�Z���	.����N�,jCf�,Fr�%�$�_����&�e�]`D�t��_=�� �2���w\��h�9��U��*�B������/�B>J�̜TB�+�i����Y,��i��Ǟ����we'x�i�͂?����՝���/����1��l\t�y/���]��;����K8��G��כ�e��������1�������5������E���>�-~7d��� '���9{���/�{-Y2��<�&�6�PE��^�N�sI����g�������ys�c����s֟2>�7�Sjh�7o�Ï?�+������t�c/lܽx��ށ�#�F�����[�}쩢�In�ozjkI���*~�;�&x�(���*ߑ�nŤ�/[��ם*]Œ(_~���"y����{v����w��;|0�yˊSV�C#�R�["�dSV��bH��F��<�/	��~y�nc���τ;y�p��T<RW��������kN?��<�ܳG��H�?e��m��������Y���D߇�&�ꂵ��pu�f4��5L����1����w7�Į��r�
�Bumò.��	�uk�Yw����\�pf&U��� �3�RSR��J��o�����<����� �d��|����O����}Dp��y�pWs���H�X,�۷�P��vJ&n��eZ}��˯x晧�z�	Eע^�M�]7��-������ސ�P���r:b�����E����H�I2(�Ұ!�Z+gDR���Cd���P=	 q�����n�t�yLF���fS1�ڹ�^~
X��*�f(E*�eqdd��6,���A��S�I�<����ށ����C+���ΨTpQ0k��M��?��'����^���_yi|d���*5>|�����၇�7\S�ᒋ����˛�p9=vϪƊ������ϻ�����7�|�Ï>��娮%�nzP��;�H�(�`�6��#=�]��g�\����2}�=��GPL#)_0:��l�;[��@˾C]�7�T(��ј8�!	�ƭ��3�M��:-[*ٝ�dУ��|�Î@}�"��[U[V��ƶj�]!$��k�
�4iЍ���:��@fm|CS�3ׂ3�	�}{�����b��f=��3��ٻ{w|����~�i��<___����%R�`0(+D*�,��N0x��O^�/�
�;<ħ��x׻G7���w��4{�qٵ��,11!���Dκ�d	%���c��z�8!J�=�J>����xQ����F��"��8�ӭh�X���<�g:�,8c����M���\�<�Y*v�(� �MgHJcQ�1i�`��RaVC �T �s;�R)���������H�Q��WE���/��/�D#���=����=v���s��FV�i�;�~IL��q]����^��jT��"A�b)�sUG~ �u���u��*P%
�-�Tަ�2�$>�;x���*��~��������{}^���B���h}����Ύ�魝G�v�$����O?����1������֝u��D�k ~���%mb\����m�����^���	1������رx�&V
J5U�+?�6SQ���T5>6NQ(��A���QC4��2"@F}ZD�j�I�c� '�IG�!ǱբU$W�6HӦ
���>��O�G���4�n��r��c��G\� +���A��jRܛG���`dUdí�Q�v�a�T����K�}o����-[:���S���r��Ǝ��o~��^{m,{�'��dn��٧�~�"* UH�`�^��+i�x�Wym�wZ�ۇ��>}q_������pç���n���u��%�w������\4�s�����s7�����侑�''IJ.����J%1�t�l_2g�~��e�̳���4����/�p��f�-�4� �|,cVW�3:[EQSu�H����DVʤ�h���w8x0�v���f�d�ƚ	� [�i� ����oۺh�0�pO~�_ �\��s���;/��B�Db�.YV%E>��� `��靆���.\���o9���������坁w��>�o�ڕ��-�����f�
;����}��{�E(d^��f�U�_�AD�>Z�=���E2�-\u�'Y�V[���֮\.��T��	�Q(�zl�N�ݡ���06V�����v�ݹsgr��1$w����W��H'}����{��̞H�,�3sӫ�����=>��S��Hw�����X�1*��R����o?9c���V̕�*<&�dhW�ѓsK4�-aqT�\q�T�Y���2��r� Ɓx�P��M')t8DL�k��1H��M3�X��:�"���D��c�h(E�'y��������Rxq�r��Ep r�?��Ac��`l��i�,I�m���-�e��ۛ��f̘~�%��
EѠZmnm(0&i�2��� �$� -i�䘒(b�6�ۂ̋��'PAiH����a�US��0,���h�P�T�w�PY�{ܵ[�L�}w��׶l����+�PJ9]/�e~L��IG��Ge��E�QC*%k�qw��#���]�%IǀTm!�4��JUu��["׈���������ҝ@�	
1$��2b���8�t��kh2(v�ᣉD����- �YxʣO�x��S�-Y����ھ�m�gLk�|E��58����Rq���4C����+�,������\���oh��v;�X�fʂD�bv�|��ظ�������\ΰ�	���0�˪�3I�X�t�$ePy8��$�X�!�}���v�qz�,B8ė�t��O>w��Q�۝M�o���>��}�ʅD����֭4,��� '5�zJ2���c��6��q�$�l87R]s�Б��;w�:�{��Y����4�ںeˌ3�p��r���k���o��8ڎ9�_z�����'�\[sn����W֮�p�֭睽F̛-�̂�3���?y͋/����޳w�k��b����^��a*ů�|��]{e:g�:ʓ몯*�kn���6;�E�;��$������X�x�p|,q�W�Y_���w=���-� �R~"����a��l����^�l��ΎX�nL,9x���������|��L���_��������ž���������o��z�Y����KN]���#���,r0d���q^����L%ʐ$-If�L��v�!�,���+�V��-�"�㊟�;��ޏ{yH�8.sG3�]�>/H��	�[��j���?�s{$�lo��{�s!����s�\��� �����C�r�a��PS��@���iq�Z�R��}�SE$����[-��!j:�@���2�w",>��A�ܳo����=SV���$A~L=�IG���	m��D00�m6.�8t��ϛXU�f�ǃ��HTʨ�2��Fog��J0���A��'�d� 0@ϿQW��"s7��KX`��矋�sN��_�i��#����p"�H����ma����޽c���ˎ�l:�l/4��e҇�����eY�.��ض�F��wp׮u��q`�'�"��/h�ԕGRy,e�|��j¾����@�� �|q�¢+�&��N���5�2���E���˖�u��b���_v�&:|��676��y�����>u��A|��߾�����hrph��f4I�r��)�S���N���5iA(�Ļ�շ̨�60���6矞z�����;n���W_q%�Pv�����1jl�u�>��S>��Ɨ�z[�b��"�hN��^���y���5x�U;Z6\����{K	&A�6�TM �=���/�7�v�Db������Vp��)=SP8�^VقN��;�G�,=�����;Grɤ��D���hU���O!DHh%�x@�F;B�\��"����\3�4�����=W�IC5I�j�n�!�ȝs�E�nz�d(ZU�z�ڽ;��q��o��d���P�:T�����RrrN��)��f�NL&�?(�vL�MZ���d���5+�ҕ0�8Q���ybM{�"��=�?��ˊ�&����?���6X�=���ZPI����W�6���*6���ؤ�b6W�#ŻL�Q��֢x�w�Q��A�J�������T���yx|�+8���J%9��ə$w��yQ>�ݫ+E�?�q���w� >.~�#��ì(?�V�{.��\}�o}`��VuYv{���w�)�T��S����!NB�*��/i��3rZ:L�d95���8�)�hӸ��K<!�O~���;8������g�Y���,��=�}��V_w�3O�v�����.�v�]1�;�z�@����3v⋷~C-��u��3v��fn|lɬ���l�a?c�i>�s��'�������ˢKbј���ѩ�a���Bj���{{{Qr�C2�i�M�j�g�7j7�������! ����q)�I�ygkkx������o�c����Z�A�>�j�ij4c�;0�?1QbD���h;�ث�U?��Ӌ�, G��׻������"/*6�;/jz�ё�x2�Ȗ�-Y<<F�w�����B����4Mon�WJ����8v��%���D6vm����]���Hٳ=?[/���RU@�R����3�)ٶ������6n6d����\vd%b��;��"U�gN���U}z���588t���B>o�sр��S~�� ��HE�d0�~��4�Hg��H�(+:}tp�?����ty�v���_���x;kh�M���-^<o���5չb�/UE��z���E������X��*]~ߜ?�|��Q���4�H�B���a5T惗�1��+��H��"U�%�i�+K�0��x�����1k�GC6�Z�11�,�9�������<EB�H�4����������,ö��"N]��FI�KvYF�[.�HTNP)D7����)�SK�ą�H��e �&�bQzR���14��:�����Ғ\�9�p��T
+�a��@�����#�P�ȑIM�]���v�q���]��lя��n���;��:�k4֫#�8�,�y)��� B�e���3��U���ǣ0Q5&3ST�#LU2�b,� ic�����֟�&~��o�+�ի��j�Y?���Z[����??�۳��=�^�h�x�g��fM]��U����5O_>�O�X�|�+�sf����z�������x��_����q��룁�R��r9M���������f��Bb Kt��������y��d�Y�Ӊzqw$����n��b��R�a������u�����ǿwuuo���3�<��u�<.FR �VQ_%C�}�|6�zi\a�Q� %�(�ƖfX�&���^2���W�6��+W�����=�9;�pW�Plll���ih��d2� �zx�i��@CC�﹧k�l��u�=��K�.>瓗]�ԣ��Nd))�?���}�!����]?�CQ�����U"}g��4շTH熎�g?:л����޾�����T*[�6R��Q;���t��������\RQ"�#�b.[*�xd9(���B�(����r2�?�]�o}�_����'��(�S��L2���W������i����Q��͕U	Q��Q*�����n`I�L�C���5\�e���.�0�G{'6���?��Ofu�>{�yh�Q%~z��,^�ti��������Lj�?)��*��o��i{��K�i��o���p6���Á%i���K�"��eU��*���#*��;�������#x �C�!�]C��O�����?�a��wx��F?����C�ۿ�Ͽ�͝�]w�/��'��W)��$��-;�����ʖ���|,y��9U����/>M�o�"�����9�aU��j訅�hQ*I��pl0BtBw������Jь�c��~�{����>:���u;uB��G/H�t�yL.kѣ�o�s@���9{Nq�QHB8���8���p���}4V*@s)Z=[.�!*3���iI}�� 5��*,,����_���.�g����s�[��M�<�0UUU3��V/w�0̲��N[�1u~���\��e�`��|�i�羻cGȹ��6���7����^_y7*����NM;N �[Mm���&����c�����S@�p)� �΢yw����z��3>��o�9��pMJ��$��αMM�k>��aZ���|������o~3��B�l.�r?I*��zQ#`c�p����"J�XbU�U ��o/X�
��WW���b!���W����w|�k��v��|�gok�[�x񫯽��4y���XʷOk$�����U5t�@F*�z��?32Rlj
����1R����r�%�ht�_�ᚡ�!�ȬdD�L�h�TNǻ���he8�0�ZU��ҍ��H�"ٺڠ���r@3mȨ���N�"{���3jw�9���+�0piL��Цa��r@F��4^W]!4���&�(U)ds�G����-�����	�O��M���Ɨ6����֦��ֆ�8YM��:��-��f�����a����h�1�)����WTH�#Ӳ120���Iu��LFN%���d��+�,��lw��e����U�l�>]'������Ų�͜9s���޵MYZ�z���jLTb�Ȏ�S�ZFp����dl<E3�L:_�+���y�̙�櫊�Qt_�`�$!��-;�Dim��������ܩT����2�� ܖuB�(]���(��r��E(����j�L���ݼˠ8���
��2/� ?�F��X�'��1*D�'�m��a��E������LI�)��8V��p��F5o(q6��M �,f�AۄX��E$�m%��(�$�Ҍ��X�4�6�/Y ����8�R5E�ı�.����X+�����}N����IV*01��@>�'p�K�+�.� F�g����4I�!��z��ۦ)��<M)����\�g��t���j��N/8�����0�0U���.�1�	��^;�J9rp<��;555�����	̉ʂ]�x��b��kj�5�ѷ�~늫>�_��s�n���?���,�`_��N�́�!�]P� �dN��7_��U���g��V��UѰ�%(��V������S/���C�Ήt?u�K�rzh������]=��a�f���^O]���[6��߻�;:}����74��3J<��S���=1���E�6M��<�D�k��Wi�K�G�E��wgg���f�wм����<8Pz��g��	Ä���K�v=��+�l��s�Y��v��R��@z��s��KIMX:��(R"�w�*Sd�$Y��[L�s����'�@_�ܹ�����~_}�t�����曛�����wp�:E�0�5��R�W�ڤ�,����q��Ի���_2eC�_&!Q�LqEQ��D� w>��8A�i�i�|���>p�3��d��B!�K�)�x:1�ٲ}����U���>t�\�h��O>��9�{��X
 FJ�?{߉㽷���I�44A���h�L�o`�ey�[p9y�ݡ�fO__O_o0��d���$##��l����i$&�u��I_8՗�~V޿=�^8L������ݪ���\�K{ِ��]P�@�\�#ձ�6���ebw��kkt��8�}/�w�8���q�/D�$��z��h;����I��0!��&�r� Q&��(�|6�T�!'��*�U�Q)���	�Z	�`>�0�u��2Gj���
�V],M-
&���{]����mZs�Y4U�
�HB��Y��&��cý>��X.���t2�#�h�_̒φ��������+˲"�v��YVe�\ܹc�Y��N��_|>����@N�r���h�����B-]�̀起����F��t�{CF F����"�+VU9gMk�0b`pP��ŉe���_��*k�v����U*��,d�Q�>WUw��TW'���#cC��HXURWrq;��VN=u���6�&N7;�)���{���T@nU  K��W���h��b��$���\̛���ȡs���J�TM8���V<��kxS5���H�ӂU>�A�r:!N}c#m��vg#�b����F/�p����m;��y'L�����Mw����sn�9�q>fr�:�!vuc`�,��LJ3(�a nB��b�0�G=�@W]�H�:�E��}i��=c����ڝ�XF��dE� ���AVj�I,�I�S?�S�KH��S(N��j���j0eŤY�����vF!1!���#����@7|BS]�eIp�b)'�%M���d���Ej�拲J�Cc�|�r�i��F8��`��` 8��]C�E��=��ߝ���n�%2���Ɠ��z�\Q���%�)M����`����
�>�Ϛ5��?�>�q�im�� ��߉�3�T�+I��S@!�x2cؐxCc��͈s�A2t&�B�i��Pn���bI-�2��U��3��D�,�4��)OS4��؀�� >Niғ��C��L� `Z_��Q����Y��U�8-�=�?1�/d�+p�(l�8���2ĉ����X�`��Ȱ��FeYX���v.�ÿB��b�7MI�Y��4ڭ1\�+�\,A��ge��d
�a�}�
5��h9�r���nEX+�B��,���ǵ��BZx�m��j!�%p�����a�ϫIh�h���!�N���믾��e`A&�c�P.�J 9E�;�������sf;���X,K�'	�BA�G�O4o"���M�`��T�!���i�L�%Q��y�����K�g�N��17)q��+��O:3��MX�h���ӿ�7�v�٥R1=>�{x��N��v%߿k����E����!�dw�T���u�ؐ8��s9>��[�}vI�R![HN���y����,袨e��J�GC���xjd"U(��;9ٰ!E(��k�7��m���>,�/��5b݌�JRy�x���M���*��2��R�kL.8������"mv����X�G7l�bx|~@'����cq�!?�!)���55�6"��4i1�J������ ���њG��w�A�����/��N 1�d�(\,FYH���"t�b���(�U�2��Ձ�-ʈ}���K[߸�֫��M�y�`�(1��8 �]N�F1v)J���b>��(B���P8PS_#x�Gz�5�w����"89��[Sō��TW��l��w�|��w���|������Y_C$s$ŒkZ&�\{��`/�s��Y1��灨���'>2�pG�t/X�R���L�ӿ=�l���z
Ƿ�T�c�#8������Y�e�>�G/&�v� �m���%�K)E#�j��Z�y�M�/+��N1��O��Ϳ$F����������RI,�\���<�`�f���������#����>��x���c��]<=����/�6ށ�	�ć�+�̓D�Y�7H~*�g7K氃�D=_.��52XV��q�8��mU�&thKZ=�&n�FG��g���98Q]�)C��C�^���G�Q�0��
߭�S�16<�jj��+񂣱�ч�W/��3�ć� ���)�miU��T�_w�66W���Jd2��<8��+W��hz�bI�MwQ�`��8)�"Y�|r"�]~�0S������\N���Hp�,iV�T\:gֳc�ܵˤ�k���ZVzz��n����Xk�
|��5���G�m�v�W	<7�eS�]tq��u9�T>rh���\~Vskc�ּX��e9��vW�#�������F�bY26 �D�D���-7�������r>[�SFu,��Rzl����TaBl���rY��9�&�-1[��DFQM��py��Nt��|>�)�W.�sypn��1Y%jjjJ�B2a��O^Rćy��+֧S]����%�l`�=+qW� ��AN�r�`����,`>c�T.?:�=��>M��F�����]��(�Q�$�z�eϹk=.�eR��G<~7g�ű���`��e=�H�Xa��:���4�d�PT�'�mn�in��88���l'���?\+�$��$�"���l0�o���:�.��p�PPs:(����w�]Wu6|z��N�ӫ4��w�"c�b\����� 	�BH�^Bi/!	��c68��2޻4Ҍ4���~���[{�s��2N�?k{�ߔsO�g�U���D�򕫭ŊZ,����{%EV�"�^��Ѵ��ځ�K�ެ�]��=�!D�$P�x��I��i��}�hy�	&�i
�y��4�����ꚨGd+�ә��h$�)�m��F��۸<����qU^ј���;v���l��FE�4dXO1�C��'�E��8�~��1N=�O}�,�M��T�Z[�n#���;���e| �3{���At��;s�D����g����$!�G�[���7�� ����yGud�
1�߆��htM����B�B����zҲ$˲�!\E�VS[Ӿp��+#�2��gn�zi���ea^P��p�Oܰn�������H��_{ئ���8�'Mg��OP5�*��G5��tV!�����s/���#��6 �ñˠn��q�Μ=y���3]'O�
�k	�ڑBͥ8
I*5�E��N!Ch��8�����K���/�#��Iuw���!oȻ~uG��ED&����'wk�8�e�j�^_�0lU�w{���s�_w�uׯY�t��Ǟx�*JU����(xBeeeK[k+�����[��<<<������d��w��'����p�o�qK8Z��NMNN��+�i�4˃�n��@$*�/��������^[�t��z��������2,��\Y�1%��\��*BDoSpSW�kNuu�-��4"�Ԕ\r�G?�c�������4�.l�4�z���c�Ǐ�L�&.\��0�����<-������
P��X�_�x��������m��z��{6m\304���I����ٺ��:9ҭBm�Q � �� i��u9g[
���b)E�f9�s�cl��%DA0F]�8���vr+W�����]��"���?����#���9��]H3"XM� �wA���q�O�ي�oY[���U(�t;�����OW�π5�s���f������R6
�F� *d8�F��	�P���7�'�k�砜Z��z�_7���*f�d�(0��Q5����}���P*�6��E��7�q��]9S����0�����{�8-G-l*N'�-�ҫMOO�R�+W�۳[���r�b&nW���^LGB��L'�dU��2]7b9͛��A�r�iUD��h��Ă����EK�S��.�A��(<jQ�	�����5���ɩQ���(�����($EQ~_.D��M���3�Y���];������'�/�����|����ҥB.7p�bem%8�/n{�2���w<�hj�����민�P�4>6y���De"�/�ڵ�k��\.ua_*#�x��@0���w���lS�U�Mh6q���{v�݈�\�F�����ib�+σK�����P��s��k��w>Oj�kթS�E��t-�>����tIs�PRڹsw.WHTV��Dy�̄,\�pb||`x�|�酋:V._b�ڢE�R�\KKMA"���/vw��z�-$*]0��raH9�.�P��PJ9�K�mC�.�7��剱��Υ��u�����e�];w�\<��͊l�����DQ�<�H0̑v(�++���F���ږ�g8d?�R�XM����I넟���ڗe)���"�W
�:��Dg�׼,)"�Cp���K���u�m`�$���P���/HŮ�=#�R:}��$��"lA�xA���ҥ�28����BE�����?�+��͒Z�̧F���u˒��p<�����
����4_US��:r��JZ�����%�'v�ո��h��Hw�).��j	�'!j4�_��t*-�����b>�I�YL3VՌ\�PYQ��,a��*����ǣ>�7Bq��6�Ɲ�����K���s?4�Q"rH����0jQ�жx��n��)���>�PX��\='�h9Mt��j�naA��|k���I�P��o���᡾ʲ��r����Ј����Q����apd���5�Bm���}n�^n#>���4$2���	��w���)�
���*Q#�y2��0p��Ν]��T����vdd�����z��%'��#�,��֯7-�����Wwdr�.p32>��`V���<B�#N&#����utL����[���>�������{����ǎ˒&ѱ���>6q���$i����&`j�_�^�T�����r�RGǆյ�jy9�w��-l������e�-������6�i6iR�֭��.�0��`��5+lK3f_�?����ǝY��u��S�bi'�M�"&TX�>�\��� m�-K
���ַ.��;�$�	���([)���6t����\:�inmj*ߴraS� �С`8/�Xa��/PSM}l���u�mfsS�H��5UU�>t��#�C�<y�p(���{�<��u��<%`~�S[nK�k��T�{���6�*�PU�e\sY(�|�ۥA�4x*U�`��U��Q��C��9x4�km�<sa��<�C��֮]{tI2U���+��E�FM�a�r���q߉�>a��.�gC��k<A���}��ܫ)2����,Y�t�K����������U���3{���W~�o������`A+i��ul^�Ij\H�XD�����c���d�qU������T.�	����ka9rdي�Uu� |/\��� D@\�����Z�ܜ�XR�e��t��l'�K�>�Y<�Z �2r���a	ЂH"�`�
�cF���/c��u�B4&v����C�=�Y�[@�t��c��¡U�VgRI��/�30�H#KsyU��A��� ��Fᬄ#ql	 �T�-H�e)Dnn%	E��[����r��8FעP�e0����8kke|D'��X���!EYQ�ӓ��y<peI��̙7��G��jrd�PԊ��*_�T6���x�/if.��
�i���VWW#�O���:�
X���*[��ig����4e4�0F�3
�E�f��*�'��4�#Mҝ��xK��<CX~�X}ͲHH�@���ӧ�$�d��(�t5��8�!&w�xvn$w�B�I�_�>���.˝^��̼R�aS"E���(�����ŬD�O%*��b.[����ɦO^8#+ں���I>	[f��[�X{��|���ζ�R!�­4����F\��g�~o��UgO=�=06:޼t�DFRT$�@^ֺI[���D��hkP7J�v(tp=W�4�)�W����b�&��U���?9A�Mf2���3�u! �+�/^r�M���<����K�I��_�hӲ�|�]��<��g���P��|��Zʹ��٧����>��~�A:�����[_���=v���o������$��K�I~0�UE�>G����������l[M}H���Od��6<|D6�e�YSSw�ԩ��HÃC��2�ӧ����wם3:�i�F:�y�Y˔�f�w�c�}�(�r%7a;�H�!�_L�@���f,� �J
P$6C"� ��B?�x�(8!ڡ�J�"6�LNOMM�����Ѻ�����0�A��A����ԃ�����GG�'(Z��kH$�pD��R����B3�V���\��.
�:�Щ�D��8�I�~͘�1�jX��-����a����P�_�x��+�65�<2��<����e```r:�V��/�B���� ��bU�����i�P^�0h!���VD���C���@S�$WVV&��XyEYcG��+��"G���i�jI�$[�j�uC�!�D�c��MM��-�%YM�Y����L��
~��D`��͝�u`I���U�n�FDi�Ӳ�p����g
Qi���~���&��~�L`��h��E>S�{G�k�GO^�Lfj�rN=x��X��h]����4힋����TP��{tI3�j}$	c���b���N�]�>%��Q���3'y�����Rӓ����J���5v �����������!M�i�Q
�ݘ$�`<�4rj�p��9�>��R�s]1�#�=��%"R։����{/VUD5uzp4y�Glmn�	v���]'O&��> }Sm�?B�"��
����x���^��&g*.���䙮��L�0��=��W�(��u����������:���	��k�������s=�Օ,��p�Q(�g�ŧZ(��"�o��jL����dæko�������<�m��P�ʊ���PtA[;Ű�` l���ч�l�]�v>��S��V�(p4c!ɻn� �k��%���&A�h��6�1�q(�^S��57Gmc�*~MJ���`H���I����B�9c(�	^�Ν;�������&kjkSɉ\&e��
3�H�e��J�B;w�kEBA*�u�I:�8�'a�"b���c�XUN�6�s�:|g�
��m�
�+B� O
��ř��d,.�6l�P__kUF�bBS��������L4�����ә{�v����fz([QU雜.oY��mۨ�,��T"f*E��(���|7�|�@?�p���#Q�2���&4Cp^���ŋLL���Nʙ��������n�7K���U�R>�"LczJn����wG����JC9�&�2�y<�%�ܪ��8�!�T�R��X��3��v����U~�@�Hӈ}�O�����o}}����?y�OK��x'&�`~�~UUM�﫯��&�G)��uS���ǎ4��R6ux�n�3�aH�z	&�ر�,Mްy��;w�z뭲,y�^�Ǔ������;t��ɻ�ݰQ$�ƕ�$�XT=wo8�{1IaiS��<`V�ἃl�q� �f1��pյ�RL4.E�R9e0;4���A���|��i[YI*C=�`o��������"c~?�_�����u��#^ݾ���iS�_�y#��߸���/��t�2�m��̴T]�inl��:%��ρ̱z�K��>��"|��_m����8��eo��6X��Bdw�%ހ_1��^�k�ׂIK�<�0~0�G�KD;BS�I=E�<��v��g#��O�	�_���d�r�����Ǔ�E����容f���쐟�瞖��k�Ϟ,����� �+*�I�$���B��&!�,J9�.���)^�j�́;USU��S�㪜߽�Tr��Ţ�T�$��>���m��<Ϸ�-���*B�R�0�A��N'M��,�Ք�1>���N��J��8rk"��e M`�-��M�*e��T0fh��|�1j@2|$�x���c��M�b�C�i����d\U�fX�O%Sű]Y�-�REY8�%����*ʅP�W��2�Y����6���0UI<>����,�G�p��:���jӨK���xo�h�U�\y���"FFӊbR�,��ohY��DO��xeuye�aP,�T��f��P�z۰u�?���膬 ��h�y|��]�.#5�$渌s�,"�l�ޢ$ͼ㮻��~�G6G�������W.Y~Ͻ�ۊE.����?q�\�����%���{�ū����Z�[��\�l{{gyeŒ�K����?���򃹭mj�m^42��-�ˉ��M7��X�jZxVX9����Σ�4�l�GYf�g�ֵ�8���3�mOL��QP�`lT.�[�_�v,�f|t�'zG���BlKÒ���Ύ������ǎ�����aI���r�A���ڲh�E|SNJ���8���e�"s���8���\25=��4�47���g���d:k���ڵk��Gw��:x��,WF"�������͍-��2RU�A�r��H�)�"��4��������7��h ��$���>�L��hk_�lm[��W^y��Ұ���pL�������ER��Q3��N�&꜋���`��a\�@MLN��S/Դ��A:99�܋/��ֲ��çw_�����s��<r������ٱ�G>߂�F�����H��(��[P?��֦s�ݦ���������8�e�QI�t.[�������y�DH�q��h��#�q�y.��B�`o_�Þ>z(�k"aЗ��dP.��2P�\@�e���I��ő����PxY�L6���G�u�#n�b>K���ճ�� ~,tZ��B��n�f�HU��:eꨛ��$lS�lxQV5������"M��°�0��B*��J�R��N�:_�G����6�\�%ٜp+��qE�X�lnj��8�:JO�,�s�JP{P����"G�,��,��E��������ۼ�lq׌5�ˁD���ڂ� 54����=�U?��s+��:�����c��(��kgOu���)���՚��r�C���lkj�5Ue�op�k�^8�J*�*J�֖�ɉ�ӧO�ٱ�*xޚj��8K����A{(W�۳�K)���g�'��sͿKRf�K�֖N����?�ZDk[CMS��Ԃ�O8�u��V���?m�f}c����ps}�����\��I����m�f��{�j�	��#nX������ڀ׫x�ڪ�<KS�P�,�n����.�XLD��t�b�I����ǺΞڰv9Xp��(>��wn�	�| |Ag\U���1<�~�w�[�ݺ��?���;q��w���4EN���c�[j�x��R*ϊ~V���1�.0�}�|����U���,á�ۧ��,j�/$�_�Ӣ8j|2�o��5��o�mc]]hdL�����0�[���n�v��q�ׂ�u���p�o`d|2��6xE$V0�an��lUb&G��e� M��������z���-7Yu#��)�Av��H6OxB�e���X$�ʚ&�5bo����˜�<eS&�ٚ5:2�����"�qñ`4 z���"L��uU��� ��Nq)�s�̩'Ϟo]��o����e�PX��؅��=�]~�bm�E93�I�~࠮lD���)Sa��f��sQ�NQ
�N���Ӗ� -��r�EHЌAr
�[m��485R M75�إQ�8���@:��t���W���Y-�77�����\!b�ްamkC��㞠�,�&~�&-��LS�+��:����
��@�&����=�	��)y;ČRt��~��7�a����=�{��:�P�'j�״���?���3�n�F�i1@s����`��m���R�b��p>�O�����ɦ3�T�bw���ȹs��}�>91]T,0�N]|i�
�����EA��s$��@�!X,4�_9��\\���g�8�ϯ�Ý1g�ΘJ�`+pdgc���_ٽ퍗=���|����+���ʶ�0o���SU��,v�������L�}�RP��RpRT5�<Bt[�I�BU���rT �IJ��k+?�;N����;[ZZV,n?t𐗡�S�U��M�fҙ�@�^�v���s�P�k_�M��"���k\U��gX��t����{>��'�q8���cay4��s`IF��;n��/����1yDU�߿���mJ�̽w���hI�]E��&�c�F�ݚ9���?:9�g����AF+XR<��=t?˲ s��6������o��<T�'2yk��#�-m�t��pU]>wa����ہp�;� F��9���y}��w]�����)�ƌ�b�t��ȶ=���ʲ��"����)����	�W
�4L�d}�Ԟ�����u˖p�޶���d��TeʒT�0P�����Uh4L�F�*%$B<��M9�������k�oG�<OK��o߾�}:p���4�m�0 `���P����y&�5��"XuQ��A��4a �*�!|�a5��y��$<i���D$B��/Â"=U�GGG"��\\�`S0�ŀ��I�v����h�������k�p[(M�4!�T5Ux�BQ�*R���#��P�T��,x nY� h�n���݂w!I��X�7�>~��s_�2K���Ց��7���(�I+�U���fd3�������3�����ϝ<��Sc�����yz��l�����L��7���o��]ع����3�.bU@��9U��C-Z��Ia�5�Փ,Q� ���{Ks�ڈ����W_}��/<�?>��?�˯��S�i�yM%^��f�j\���'�����]0���֦뮟Ne�t�-V��"F�o����:��K=UܫϹC�х���X���ܵ�V����o��:�B�7_�]=Y=uw�V,J��|��T&`Uh�"��c�%f0�r�u|`�UExE�2�H� K��;���-�G�8}�t*�^��VUU��<�0g�V񆕋��ݨw(e~�����#F���U�^ҤH�4MT�M�6�������U���D�ۚ��ೊ�z|���ᰠhF.�[����w��7UUc��,�?��l��x��d2�����Z�A�e��6\�	G������3i�.*��dm^�jͺ�����0l�c��
4���T���2��nkoTUT$180��g�j�D�L&�����tz�uA�?H�Z*d	�`�Ue-'�6hs^�P�4������`4U�ձ@��.^��oh��P���Su���������L�E�(;%�����9FJG`I��Y�ќS8��D��Ȋ\��xD����T �� ;��Wlst �	�6�۱�먒�<#Kq5(|�E)7�v���� �m��`���Sp�<��e�|v��ȭ�q��]o��C*��ߒ��v�C6�ˢp�aIк�I�U�]��=Q/8�#�8Һ�����|�����0������H�P�"��N k�������% ���X�S���/`���+J˰(�]S���9ՠ����)���E�JV��"�$#(��	�	�)��+
 �	E1m�\F�T�[��^���V��6J��D�a"-P��u�2A"�����9�<�g�֖0I[�~��_�HT���/`��D�z�z46�����ۦ�I����L7]��f"�P���+�森�Ł��(��;��O�(t��]�ж�Jυ��R�x)��u���"ί:!˞�0�T`��"|cf��X8,S�H�Yjig[Q�M�h�%m� �8Ґ���C��1,�x�^L;K�(�@w�k�KW��o�G	kο�_c�(�Ե,V�_�Z�������yC���>����^�V������/�A�Pd����߶mttL�巽p`��6��	qJ�(u�
K6�c:c�mqbC��rg´X��������z���Iax�o���U�^ysٲe�
ߎ]'�|�-����m^�џ����\a�(f|,���Ls��"l��| I9��,�0=��Baz27=n�>]7h�c0�FZ�FC�O��<?����������,t1 B��\ !���ʁJ 	���V���	HLщ��lͤK|��q:��H��@hGEv1c���ıs��"��i�@�8���3����,ޟ�+7l�c˵kR����O�My��O�6]fZ��E�S&�d��)�²%�u���o~㛭5���9�tE75�����t�8��M�TY�.{�f�VKH�R�3���ǏGM� !P1�o�^�#�\*�-���rX�S�i!eޤĢAh 0@Ͽ�	/��hC�ek�W�2TNm*1�Lq��[����������x�3?z&Q���6-K$j~��y)�UTr�H��>�qU�u,��͛�c� 0�.�w�.��^�?�ĵ��b87��#1�ts}G�t�-�M���~���0��_�ԁ��/'�p �(���c11+f���r7�;��;y�?t\U�W4���\�A��/X��F�l��8�m1�]����YW�"G u���J�(�f(��3Oh�c�鐧����l��,�^��s���'/҉�%Q�����LT����.P0��:nͦ^�ŋ_�M�!�_Qq��@s:�[N���=��$9�$D~L���<$:�f(���ɩ���Îŝ}�#��/��rYM�K/�<:2TQ[/���_zc��Uͭ��=�ئ�Y7�8Zg"95f�Y.T��9��f�|�bE"ˡ���ue��\6��4��Y�?��`e��'ah���M���J`�C�,��o���6n�+���gK����}"��@�RBƔ��bc�:4I���S馃;�a*�68�S:h9�H��L[J��t�F�s�<:*����7:1�J=r��<q����<%�xu�(A�>H�"d��0,��w�j��r���9���#��RK��49:��f�Ç�X#ɉ�p�[�et���P3>>�LN_�880�nY����p�;�LK<��έd'z/�o�MZ �|p��ژG-f/t_$~��<�鮳:�ŀ�ㅍZ������������Y�)�3a�â�eb:|����eKM��58�ruj*�d)��XBV���t_�P�,�j͆���
�y��_�����^n�\X� ��E;:�(Ѻ���(]�C��
�PU)��u���j94��^tJcNu��NFv-�"��S�57�B�,uxU��c�'#K�b�N��7Q��u(rXⲬ�rgaдKى��E�qh��4��©r�3��V?;W���
�oa���144����r�����?��O�m'�
|w�}���M�����q���jYGۉ#�emZ��r>=
�޹zz8o9�(}����6xǖp�����!�>ec�Rd~�T*u�}1L�#zn�r{(����?���_ D���tz͆��N�:1����Lz<�ۙ�t.
rC����cj�K����U�ǉGC&���x�7؛��eYQ$՜����#���$�7�sP=
C�r�8�W�~$��`Q*�2D``�UP��r,�8�^/�H!�i�qP2�)n+97n�&���,�3�dI"�ւT�a�I������"����`"~v�w��U˗�[��ͷ��_��/}ipK�,�BamÆ�
�+
t���w��()G��?�S_$����
Y��o�a}.�8t��H$��������j`�S�}(ԡ�����q���ꊡL�0�fx��@�W�G_u�R��F	b|zph�P�~J��"�����X_�2��KlK�1׬K0aͯ���\Q.'�������=#S#L����]�D����򣧞in�?|� �3�co�rK4W��~ĺ��AG�"�4ʔI���KC�Aj� ��t.M�FSE��1�wf�.y7^$�O�Kj;���,Q�=�ϜmS�X$��)�Ylq^��:�9.st����{�}��h
-#Ul�~/�U8>��-P�$Â�D�}� cu�p��$f�߭���X������B#S�"���/VWľ��J��I��tuumS�����<|o�Q+����Tѐ���p0��c�O~�.8��P�/����$3J`�f��;=��΍��EI^�8j(��ųH�S�&*�A/�ԊO�ؓg�k�}�婈���Z,>��ݧ��/�&Q�"ׯ*fQ�X�KY�,�
z��h4�����d�)p�$E�I���uKS�B6óLvljb|´h_ �!��4�㡜�-��aF�w�ɤ���Λ�h��8qu� 7pc�'f�`0�qI	B:XNoS�
�E*��w��hg�X��	gQ�� ���34<~I�	�H��DԂ��1���׿�PC�g�u[����� �J���/���xŒ�5�N5==��]l�4�T�j���xn]��҅��i}��{���E�&�VlI���/��j�H0\��&'��x�G?���GLÀ�`h
��#�R%���$�ѳQWG�<�$���Ϋ&7�0S�I���ho}U��`,�P���t2ٸh���x��_}o˝]�t�V4hK�x+-��ҋ���z-�}�$
!�lGR�p�.a�Esu��������w�Ŀ=��W��ŰWt��mvvv�w������`�n�kkc}�i�L�x�����_�������'�$K����TU���S 
��O��'������ލK;�+�9[qPY�=������/X��}�Ƽ�:���.e0���S�D�.=C�l�_B!�����^U���p̲�2��pҁ��`e�O@;��f�8⁔���X��n�]j9��3Tj��*��\���꓄b�&M����$��C2�l����fP�LV��xye��Ng�L��zEgݛ����^!�i����5���c��bF�;�^X�R(I��,n_�wכwl������7�h�{�E�g�aɧ�x8|`��֖�"��B���?���7l�@�!
��c��>�r�l�[,���0~?�z8�^��2�ES�e}M���p(
���ݖ�֑.���,��ǘ���h0'����L0;<<gs��R�e[ �,Љ!*2P�!��q�9�3H��E�'��#gX1�~�����}��C�B�B'�u�NTV���c��{�Y;�g�\����)������]v��oּ�b��%Ek7μ�(�j���Hdȑ�b^&%����,e�EC�-�Do�(�4M_��军��bK�B�#�"�(<�PM[aHE(D�vL/'���X
j�b�R�}�JIj1����.*
�IMO�Ri�秧S�7����qA8H�	�XRJ1i���'`l����U�����}��@&B��Q��,�X�ڍ�B|�qϞ]��X�
�K�.NTT�&�\�3k1��i�XR�UUJ!WQ]G���n�O�����7����~��G�=ux�k��y�Vm�$Na�宙RA3A�L	Y
F�u�஝8��u!S�2AZ�e�!-�,Eҁ�����_>�*�+�����P�h�x�807c���S�Q3B
k�����{@m�E��;|��Ν;%U�Xl�����=��( k�n���e�e�5�SSSp-pI��fi�9�$���í��?}��c���vOgn©q©C�r��R.U�G��@��r%	)�^��}�/^����E����u�p����XYEe<H���;���sg���-7��:w�����z^���
�P�5VQ�O�	��&E�8��q,!)DF"
�)�fZ1����[/.[�9�ɖ�W!`�N��~_�o���D�d�cM�A8�!�I��pM���kY�aZ�d��\�V0@@GZ�5=��eQ8-�ς}A�m�9����u�,�'s!8C���������[�����J�Bc�\A+�w���H���������'O�\��҄�H<���
���%]H����]�U���rL���e�FF��O��j�]�qW��hP��Vx�:��؊x��Lv�5��Z�t�šq��T���b���\���G�2)�4`Zi��ߘ�/�d�J^7�d�h�A;�MN%UJ�	^�t���Db������B�b:I��2!T�V��-�����Y�.�
�%,�;K��Q�E$�R�B�C�⏞}����x,��xbqK݆U��Z��5����衽�\���]K�tvttlX�F�Y8��bQ�w�.Ɗ>6H��^bdTݺr�*��>r��?x���ܰf5M���|ɈA�H���K�PwN��a�h��	���=�p�z	� h��l� 
���4�*�_y��d~���!�R��ʇ�� �l�W��痪A�4ڢ�e����@ �����ۻ�/�=N�D,�v٢X,V[]+l�! q��Ⱥ�������'\��#��L?&�1[��L\.]���u2h�ɳ#�A���,nim�Y)d�LO�{��;o�	dk>����~=��Q�FM����E��i/퍚
+��G��MH$�������!hI�Gƒ��:� U���k�-_���́����E7���1m�B/�4�s8tI��(�E�
�xA�ex#�O�d��э�FQ*�U����T/HS(���LҌab�Xk��7�8|N{�YE�%�d8�?�  Qd4���������{?{a�h.�X����A��B���_ھ�U-ܺyݪk���o�0u���U�I2��� )1[c�4��7�}�SP�w���>�?�.��I�������<C"+��H��>�^��/\�m���â�0%
������ԼI��ڡ}UJ2����N(E�i��������e��`��\�G#I5ÒL�
L�޽�cզ���E�%�RT�2*��}ݺ|q�\(�Bu$�e9����.���ah]71y�[�hh�������X���+/���
^���~�s! �L.���H$6M�,͂��LR�(�e$��)�[vJUr������u��^�BNwܼeͲ���[ߺ�#װ�E��Ҹj˜	��mX�m�����������m�]B��~�M�U�t�Ws�W�;��n�#���u�.z�9Uj-q��t31�cV'�:�|�u���^t�m��B7H3�
5+Y?�����l�F覇"{�O}���>�����Em��u��X>�IYQ��D�\�B2�8�a�(���>�?HK��bg�3�c����Xt����&-CÔ_��G��)gRQ/�dr(�چ&�%uݵ��[�q�or�Ӝ���L���*C��O������+��ޔ>�����$�2�74:����[j�����Ny�:�L��=H.����.�#��zрmF<u0��ł$�a��� �V����t'����U)-���y�pB���	}��ԼN�H��6��:�����+�;fL����C��]88��Btn��v�E18X�:��κ��fx@Xr3����ٳ{�JN�]�v՚5 +
��������>~�̩�����K��|AQ��X�qR�w#f�r�'�bL���oZ��^�0]���ʅ��t�"�}������tɹ����W�������EoP��r������"ᾞs6,�麵o��b�T�,/ˤ�_zq۱��׷F*�X������;�l��w�u�_���}���Y�<7=ViK�%��-̭w��/t���M�;�dJ�d9G#*�ls4"o9�Z���j薝(��4���c�e�[��$���(MS�>����L�"J'_=�7U%�|�����^98�<�3��-������}��K�ZXD&�V�yIF~�,�X��<�#!o�F�L�i����Q��,g.ob.��E?��ɉI��)%����E�#�Gd�7 ��0� �E�����dt!�Y��+_7�s�=�z�������2ΖhKE�����bww�������?���K����X��}Aۢɡaa�ITN�`�K�v�����
�P3�9U�4b�,�w\�#�8ڂ�0p�B�"u@�H��4	� q #:�]B�.m�uM�N<�ů��w�3)�p��||����S�z@K�I4x���ٶtŲ�4j��<3Y�����s��e=4���$��@����S}��}6�pp戋'��,�l&�h��a�j��X�Pq%���E| {���qIb��˃����5cJ�9(O�*o(�MC���-�1Q�&���¬��Wk��.�X�ȟ$ +҂&����~���V�^�t��_��646o���'N,X�\��m��~�M�Ϟ8155����1e�1-'A�XS��f	JSz:�1,�(n�2�a��?4=GVcC��ӧ�\�a}X$�kk">O]mM���$X���i5��(/���������Wd�B��A�B�#z�<H���7�7$E6�5|��_y���5U� ���$� �.�;�3��W��qhS�?���xx�<�r�-�U�򼇪����OMɹ<,Z�/��Fǆ;;����3�N�P�dQ似��
����N����\���?v�Į �~�SwUƹO=p���<����d�D�HD�y� �Ȧ�x$�O&e���Q�(>� V�_`D0�t��*��L>�x>����X9�W__�������1�
_�&B�K(S�C��������l3�drN��Xt����XB�!�-�v���.�$��d�Q��Z�n�\6|���=���_6�,�U=�/��rS*�7��itYG���7s#�ى���E���%-hchٴE��LE.������
�t��)W�ɨR$9s��L�Ω�v(D�����mZ���NEey�Du}G[�C>� H[�R֢�X<�ϤA���yE����/@1f�����i��$E`KBD'-d9��{9/����ځۤ�㋄=��4����a�C�b�����
����Lۀ9^�,�Ɣ[. �z���[AU8��8�ct8�]��<p�� B�=��}1����GoK��CQUՋ).W2�V�}!���~������x!&N�!���Ց�cٿ?E������S��x<4x�$Ѽ��~�����蘥���}��7��-)8�������p8R,ʢ�W��$����k�5���PCSKe�g��7��*4-Z��P64m��o�v���?���nX���>!������s#7��i�f�'`'Z�ʕ�RE�}$�꨸�B�oR%i���*d3S�b6=5F����ۛLf�3��+�054���LTFEۓ�����������L��g&5ަ��\N.�w���mj��~�Ò$m}"��*�7w�����,M�t���o?z���*�"�|���������p�o��꾳o�9[U��rۭ{~��M7�X^y���A vǑ����cgN�I��񠯘�h����>%�*�Qt�b��\��N��UE�~�R��+2*�9�Ԉي�+9߲uI%P$st�!�����=�>PS� [������W�Y����gҹ��ZE�Q���E�B��mCwhՐ�1����%h^3L� �b,��1`cPp@t���J,ԉR��lH���&���|�;>1�+*a_�����XNs
pqհ���k�	�@`	7���P���r2W�,��GH�j�$�� r=�G������T��	n��]D���r�58"
���,K� ��1���9�f[aл4 �K6ӻ�CT��t�f��u�y��ճ�(!����>���qƩ�CǛV�V��Ha�I\�(�@8����,��j�E��؝�v���+6��>�RW��W}����K�"���ר��-;� �
V6�o_��X[c(���օ}��O��5n޼9�Ss�"�(k׭-++�d����W��Ł��xMsy���f�H�KT�� x���l����ekRi��O������c5E}��7��vsm��|������$/�q��ԗ^��k�n��;ߡX/�T�4T�ց�w�����ѪD�sQ���{w��,��{�&iŢ�(��m۶��Ə��Ǐ754���m�����/�J�Jc�ʤG7m����rZ�3�ni�����v�D�ww�)����H���ܰa]y��,�88tqp8�tA:/�>�s�'?�����4H�xw��M7\'ө>�ʪ�kz&���#o��N�蝖xoY��\����k[3C�?��߹����tab�Z������p̅>��{��E��;�#�!iT	���]���;�C�c�95��r����_���W�C ��kW.ax.��#g��������t�yyN�dp����04��m]�o&&&����ؘ��eX^1M���*��|������#������7�����*QQWU�����ːh��E{#�J��4��a�F�vp7v�t"��t��#+��2"O[��G��Y̯��$�.~� 9����@��ҰHM=L��Q�,�Z�A��嚲h��D{[���	��q�'y��-��&�yE��k(���fŰD;�;\���%g�J��'����L���f�S9C0�a#����Uj�A�:u�}��,��Ӳ��7��|&8��%+Z[�(Kh&�#��g�&0�ӹܠ�"����{�4��&�w�+���FϚS��ؘ����Ç��z��ob*�cED���,����?�g �9z�.9O��"mcJXL�E�	n��!f�<�"�\O������3�������������p<"�Hmm5ˋ��S�hMSEY��!
Y���)=t�'��TS��������?����{�G>w�?����6�^�P�Ry ^H4�܈�V�E�iv�AI�m9�h�eS�k�g?�0I�C�o���<
���=���a��x.v�f��W�{�o�_����/�[��t׹D,�h&�Z�֖��h��7@�E�Ou?�Їu�<R��,�l��T���zw�����sa����p��cA�ƣ�^]]�����c������5�Q��������&SHل���M�U��'�|�����s1���gsg��������?]�����M` +IΔc8���Gxu\:)`;�i����0��8}��!��[J�U/��a�����ISu-59X�멮�K͍��3���q Pg8��E~�gE�p9�I
4_eU5��_�	���AU7"��?&�(�_XŲc#������pí[n����^��[�V��ps{���v���Ƣ��iʭ(q��P���v�����N$��q�B�94͈6͓4���+��`,�5x��G
��.�CI�a;��0� c�H� ��0i��y�&�����p�g�1&a9ɻ�G�#D�B��pE�,�.d��8k�%K�v�55\�ONʲIO%��7�>�������teM���u����Sk�N58����CH���?�E0����o�f�%�s��G�G���Ő�v���ʎ~���R���Y��4��_�N����[1	/�ܡ_��%lݺ�������a���H�`ț�L�2���aD�`Ze�Dye�-j \.U(�#өL��t!��z�̇�ԣ)idj�+�Z1���]���J��������޽��a���G@MU%�L_���[n�����ܙc�dx�e�d>�*,lYض���뼁	>i��Y��x4�ge��RS�[�d؆�Ⱥ�3U23M�S�
\2Z�'��6h]�c##��ի;��Z�8t��G>{�/��ɛ;{dMo]����E��G8�}�
��-���[�.:u�0IV�(�gNͧ��k�{_Owar���_y��P4B��ٕy5Gxu�s�9��k�������|������,-�l��k�~z��Nt�f
��D���A�WW�i�����g��<v&z���9�ц��6�z�����<9����o��5+V~����M���𹱉������q<[/��y�e�tQ�u�"C�hmc�����Ӫ�Fnq�
�5��������������pq� :�t=��F`':�Yp��l앁.3t�0���fS���w��J*�aoT(��)���d]�٥;L-��
8�t7u�D��w��)�j��H��`!57qHb�p�)��B�R	��J���
��඗v���k�Ս����\v��k�z�{O�l3�hE�Ξ�O=Ա��F}YA���*1���4��qy�41819)r�Ƈ�._9�/��KWT��l����BUeV�*�D"�gƧX����8f����=�q�Y�R���� ��E��̱s�pEE���X�݃l>�����t.]t��W��i�`� �j��q�a٪�c�100���e�]����˲U�u]߻woGG��������S�%��w���~�o�:���D|�����Uܹ��&�ɢ�o��(d�JQ�0�|6}��������'b���s=��)]ӽ�Ԟ��Q?�e��M7��f�N����U:-s�J�U׊���|��N�2^'B&��d�}Z�ǫQ�����˯�S���nپ��5U[[�V�p��c����7-����ʨ�e��Ӈ��F�������U&jc����]���O�o������{��qUi÷rU�<9�fF�rp�-��1�{��,�w�%~KX�e�e��ƀ3�ؖm�m�rP�(k49O���\��{�{42����`]ĸg����s�{�{�\כ�S���#�u�5zr���0`ꬿ4FXM�Y�\�Tn��br�+\R"��n���[^����- :�g���_�B�KcccCC�MM�V�Z�j�����/���e+V��kj�0��L󢱢�՝�G�cu���ҫ���_K��]��t��Nf_߳?��d�����[V���ַ�z���T�`�L2U
��P���i:��j��u�60�嶞��$�[�4]�iʥРH:8]��� 	�	.��>I�G�,�5�}�T�$�;� H��JL�p���dH�)�`(k��e��hVE��#���.Ӓ��y+�)�����7	$�e���][w1Q5����C�5M�C��M��x��~� �^zq�^�gd�¶m���&::WwIr	�?|�Б# gL�
 �2ً;��n��S!֪o�+��q�X�������V�<��+�\��;GqYUӵ���W�<�\}mM{{{�&s(�<�*a�[Ć��h�v}��ZH^�r�\*�v�i�Rɴ���jsd	�ٵ����Y,�糍��".pL��ӻt9�|E���H���Ւ��[�{�Б��� ���ܳW�Z�H�\����	xK�o���{r�𶮔�:��]g�qʹ�lx�3S#���lza��%���i�����^�e��f���/��\S���jj^�`�\,������¯�ı��;o/�bA�ؚ]*iŜ"��Wg��D���70;�|��e�A�QJ��#����v��~���������,]�K��C$6I, ��-�|E$��ӗumٺ���55%���YW��-g��O�7\w��?�⫯n�x�j�TeS�ە�b��폓��-���Y62-̸��{B�\F���HUu���Q��c%���U45���{�ϯ����c�a����o�������Y��gnv.�ɀ`��ګ@bnn�୵o:��������{�[�;�uM7��ޒ�5�D��;���_���m۷O�%/��P���������6������cvZ��g?�cS�y\b�j}sK]c�nZYUpTPb��K2�H��§Ͻ��s6�Gq4��G�����<�w��d*���M��M--7��],��i��������YEUA���>���哯����[�&H����W�[�R���-[_�ӿ_�0�N#��>&P/�x�U�X�t����:��#8P䶉��dx=3;����Q\�a��2I� ��Tp���\�����,��X:ǡ�mϯ��5q��ɫp�`e�u�E0����k���j0 ��-���M��շ^8V�̕�Y�����֒ON�r�Pm�ei[s@2"399�������޹�u��K�~�.%'�颛'\!sw��#�?
P+�7�v��?����B���P�����r���4�;wSu\g�<#R�g�	��T꾶t}��}�?�2)Y.=�iS]���3΄�Ţ�tft|,	'5��UC<ޙ�C󦮂�Y���p����0�<�R�m��.km����F�X�f���bk���!��o¾���Lݜ���Y���9藎�P��T�Ucݲ�-�<z�J-��֘rf٢�\.�O�9؟��׮^����߿���	�ndd4�б������nش4�Y��պ����?6�ߦc�<���fSKC���+��h ��v�կy[�b��{���<���v%���G֭�e�\:5��hܠ��K/��h�2�`&� ü��/8m%�[���������{�b�k��7��9 �Mk��4�'Er����"��ǼDØ��#�
>�'w��X�U�jdt���}`8���I@:�I˹lzvfth���ى���4X�MM��絵����N&�E9��z �|���E�h�X*�i0�CR,�Ś�g����_s��u�O��mA��_ޫ�Q6_�M-�DD���������<�̋j��*/zD�����l I.�k[�@�⎵�T�r��)�G�M����^u����3[�]��@�\@{�����W�<44�e�����}�&�dQ�X��+���{��e���łJSH���vw�h����iED3N!��a�BU�{�k�y�	� ��(�'^iӽ�d�^�M�J7�yD8���ӫ�:���x�
�0$�-�pq�1y3��]�אGț���f�r)�����6�0, /S-�v˝7\{���&Gr��9��G�rH�V���8�d�B:7�U�S&�(�̱��Twʥ+��7O���Ё0z9e���d/ϼz�eh�H���麶��v������׷ttt���	�b(����.C���HjB1�pN_�l��׼긭d)H�V�>��M��Hg�j�'LA�Ē:!F��ښ�H<&R!�Y��;ogm��.:����O����H0�	��[������Fx�-P����w�9.��v�$�^�%���|"(3��"L�,Z����U+�e�z��7J��F�wpj(b[�[U]�L�x�֕a��ŀ��ljdT*d~�ӟ�J5���?���d��f����%3�#Kw�
}�I��*��M�)xL�$�e�=�O�7]q�O��{���+���wZ(�:;ښ� B���\R��X�,�醞�5�����p�����3==k J|4�uvfjbjr�+kןZ};��k.޳��}�]}�MsŲ�V[�ټ�w��>O{C�m�U����gAYj_�r���^�J�m�k�`ڴm���Ys.�/�/+�ڶˮ�������ܰa1��F4�G���	�AK��q�P[{xl��Ք��M&���gw���O]w��<S���>O�N�7o�6g���T�M@=�WR�B7�.4���y�G�j�l��ׯE�2xP5n���ٴ��|�ݼ�f����������Kv�ν^߾�w�*�G��X�&V4����Z��"��m �l#��׮Z�~Ͳ|rb�H$�!mLfF��r�bEc�6�����p{Q��/�p4Y�W�:6��"+��H�lJRX�w�4���
�L"���SOv���^�jbb"5;�R�gʲ��xn�e1ɺ�4ɓrc椰�k!v�S�$����vC�4Iªf� ����]n��Oʈ2ennv��j���Rt,���Dڎx�����Z*��TrrܴLUW0�!��u�Y�����xI�"�0h�6��d�R�+T8n=ͱ6ƨeY�ҋ*mۂf;�Æ�<n�Kq�U����������񥈾��6,�e&"���^X@�_�����	Uy0��i��#E��Ȉ"�`�W~UM{x;�FO*�?{P�)I��'�+o֭Yջ�Y����v��r�۶��1Lm<V�������d)�E�y��Ro{<����cc��5}����&��n4u����GP�V�>؟A��=��KV�\���&��h1�ˌ�>t���x��jPfN߾gg�V��D���ݭ�+�/�lkin_�F�����XO_o����Ԧ�΁��l|��IqȎ����&�D���z�i��,�<R:�w�sy�K[�����.��,�[��V�G�9j�9Ύ�<�ΖAZ��v:��,Eq��/9��|]��Lǚ�(ō%���$܍'�N�[�z���?��1-���U~t�f�6Y=aPT��������i�&�(t�y�����˖�{�r*���6XA\����߽릐 �S_W� �ar4á<�������xWG; DG�9V
�<��|�X���
D8�%�V���,+f���
Oӂ�Y�� �E	����kv�����xI��e��R.���������`2�X��e��F ,<��:��J����x�K�[�*ohCHA�[�H�fH��j)���؊nZD���Cל�`2ڶ155��z�w���MQ;Z�֮[�n�2%�I��=��7�lnlPg�|���nik��OO���׋����#�t�-[�>x���G��8�V�fx�w���5���0�ش���l�+������u�^ڮ�Kp*�I�%�[.d X�J��bBm��-����"�B�N�x�n����p�n2�[�jSo����IE���BA�:>�iaq��_�3��� "�\.��{���=��cK������/����9�q���A).��EÙ���((�R��	�5�#y��d������|d��Ç�;::u�H�' �'�۷���_O�L���jS}�Z,r���7939|t��w�V(il~��X��с{v�&0��T����{���J��cO=��[��	�,��9%�<4;�44�?�+� dL��w|��x׮�;kB�����}>�K/��a��#��o��Ɩ���:ôжmۯ����_:�O�^����lj��2s�_mf*7�F�����zIUk���� c�����7�n4g��4�]N����+<���$���K�ktP������S��X�Ϙ6��VK�S�Ө�QT�)���v���k\�;�P��r��%�����q�tCs3���!_&�	�Vf.����P>[p,��Aq��4�-R���C�`!�Ɨ�9?/�,�&��	���A�c�,ok)����c
�)4<8�kY�щ3���e'�+5�������;D3(�P(����mۚ��/_~x�p]]�B�$OLM����Y�\*'��P0��}g�J�"�ˬ��(�������	Z(<01M�	�"�����#0.����x�fJ ����~��9���l���u0(��,;|� r��S��С���,&W���IDT��1�2���]�i�a�cc#}�z=����~�ç>��ƖV�F�����,����B����(��gK��I|��wG��ƹ׸�
 eIKs�M��3臘\�ܘtE��Ȋ@ �K�	�ݖ�.'w��E��o�T��X���>��r��,���-[|��/g'&3�,˂h�-[SʥBq����{zz�:����������z=���jA��ˊ,��}��8�w��T*�83#������0::Z��$I��m t�f�6�H"�F� TZ�R�t[�0Nu���D=�𙴬P�e����Ӳ�����)V@
$!�L*��Z��"K�榦,�edY��G�>��a9���_,��P[KH��ގ�_�|��������Dލ]v�.�ˈ8��3J���[��&<�&�T�ÕM��؊c�-���G\��&~��y�A',�K���t�����~  ��IDAT_W��sp��CkWZ:�y��	N�
T!?��*��fA��8����h�>S��['"�]T��y���h���S�C�ˡAj�Kb(�;<���Ьh;8Dp,�6���7��r��I�@Y�av|�PMM�-xáp�T��:K�C����g Bخ`{�<?6:�r�Ͻ�2\t^cS���u���/����-�|��M�[�vQn-|�����7���l�� .�� @���Ԭ\Q�yV�z@�kX��0�(�q��/��6������l���,�������r4��Sg�A����x<
����H� �F_�f}.��Ʊ�?���)(��ˁ�	ԫ:���f��7&h�I�]ʍ�V2�]f�?XdBR�0�#ͻ��i�r/��$>� }�JV��=t<Q�=�IE���w�n�a��~���� =7�x�SO=u��C��r v����M���8�nin�����xpf  ��'��qM ���ř�9P����^�w�=^���o�֭�u�ҥ}+WML��̅��9O�b�mGw;�ă�j뚮���=�2��Z���v��*Z9�IS,��N�e�+dL$8(ֹrp.U�V�{����B�����-9�ݽm��%��Pc4(1H-�v�`8�r��zt`�&Q
ј8ˏn��������[G�pO�Bw���+۷C�t6�&�p)+Kc�:��s�i�p�ۖ�D��a��j�:U���mjA�-�j�R�B�*�ݪ���ޅ$�U`�/��tӰ���	��T@���[Y~\���P�A� 5@ʿE�-�G몚�g�Q*�J�$�/�Gd)�CO,����-�x�U���duZO��f�'iǞ�ƸK��7)J��x]�;]`8^��C{�����X,�(�����*uQ?���^�2���\��mё#GJ�,�}�S��S(fzw�����=��2�}����&��^����9���vU�|ҕbĀ��yU5)���4d�H`I$>
IV-S6���;�X��q����tLd�ͲM�+I�B����v\�����"�\�Dr��2J�b}A�с���I؊�tJ-+MMM�l�b���P-��4� ��%Һ����v�� C���-kQ8��aD+b+��qu�S��q��E���n�>�2A~�����&)%d\�A'�eN��.��[�����p2 �9zx�e۶o߼e�ZRHŕ05>�fժx4����=Q� ��F9�,o���搋�A�e8?�h��h��	Gq�n�,��`y�M7
��'y}�m�-����7���DMc���t)����l��f]�χ�� �
�a�%0�E����q/�XĄj�����|����㫯��`��Ç�{׏�-�	x�Z�*�A�a�z��E��111��T"l0cJ���Hb[*�����}hfj��%���/� P3=���Z5K&��r�s���J�V.�*�"[u9e0ϸ[�N�>�N�}ۂpo��@aQ�K�Iy;f��H�������2b��Kjs<��M��J�t��+�n�i<˙�*2���{�"��96=9���K�hL���P�Mq��pY$��	�"4i���7A�����|�-�8�<�G�~2Q���KW�ȗG��-��Ms��e�3�V��R����%�A�O����'�[-�{C��T��4L%��m�E�kO?�衣�W�94:���(�mP�*&t�-E$�s�'�4x��^�jR�����7�;W1�3�j㗞vc}m����{	b�m�~�����.�5��!L� ț�`#�����j�inn�D"�4�t��4�J�[�΢e9��J8+����e���ۘ��6�2)�@�Nq:�~�r�<������!�M���D<�-��9�"�0;0�2Q�� {�i�Du���v,�nR 25�N�!�-שN�m�ƛ��l��C0�������"|Kc���Ɣ]��w���0����_���kW�&;��S��W"�nl09�.Y��z��5㕭�m~�垞8~{���x�^�7�̀��#�Ȗ-��j��,��Ӑ����DqCss������z_z����¡���yl+����l��JQ)s)��8_���}K��2< ʬ.�}K�_q����{?b�u�ր^[��FK�&���Gzz���D���q��I�n8�=k��O�p.�+FQ���&�5�L=��'_۾=���ʫ��xCcs틛�=���_���m}�߉�;v���g>}�%�wףUKú�#B�	&�ŭ/��\K{д�S2����3����l:�mb�a�����a���ˁ$�y��j0�4G�}���!ɺ�𞻒������y7;��(�H���y��ñ���-]�{���-H���O�¸"�U�VF"A4�l�æ��>���N]G�d��*"�1mQ,ʰ¡���,�ڸ��ZA�/j�l�?��c��^���ڶ��&hS��<`���AW�.�6��ZU_:��q�F�F��LO|.W�m�|�A�gQrv*�V��̵}#+O3���ԙJ�'E*\�4��!����l� svfv*[8���Gg3�+Vvw.��ܶ��|�?���?����H*�r�zU�%^�di8j�
��8�aEq,���422;$�92<�I�ᵽ &
�`-�%����IS���H4>5=G)����1.����xB^/����N�z( ^w��'��>��e}Kҩ����o~�����Y�B4Ly}�7��=Y)13����7�����w_u�u������O�ybn6u�5W�3�ihh�him	�w|�T�����aEk��V�Xy�5W%"A�T�$��c�\U�g�]п��IE��� U����>�L��y�X���;т^8<344B��(a?�������j ��<����|.��'Ѕ�q�R��V.%	�sm��ʊ+�6���V���KQ{:Z[����T6YS�}?��7�j�ZΊ�?����]��`lCKkC���C�~�L,�8���:r�P�A�$0n>�	�q<j�J_z�������3<<���^ѵ�/�
�q��w�<-K%�*�R8�������������Ҭ�vQ�N�-q��'����6#�(����uc~W��e�m���gaIZYeW�;��?�:��XAA�Q�\��W�8\�����(]DUi�w��XO��N<:<�&���)&\d4���e�r�Yf)b�c���3����G,����ݳ/��f�gێ]���-@Q,�D�f�Y:����f*�3�BF6f��I�nG�s�,ǋ���G¾"��ꄠ?N�k�����3,j&/�[?��5e�*��'?�wCc�G~����U�]vGD����Ev�c��l�v�ǧ�p� �xl�7��!p���m[�t����֞�������Ri8�^�������h�&N��u��V�Y܀�&@t6�N�%�Ţi��n�tQs�jQ5L0��[����<�f�H�"r,8Y~�?����[�N;��� ���4��r�)�,���4����dt��%�7��K�,Z҇]�]!D���^x��<�^vYGO��#�����}��(�d�ܟB��2��C����.D�|׭�-qYF���7����Ͽ������Z��ͯ�|��G�c����6�|�qR����F�"]y������=`�/�8ސ���Q76���-��ó�����UQUP�n�t!�D��Ԡ����\r�q�pn�e�od���N{���L&}��vn������O����~�L>������&�:�&�&��j4-b;t6S~�7�|��﨏#Է����%��1VY��ż�ٙS�t>9u`:7SHɵ��K��p25Y{��rf6S,���|���)�G���=���<R^-���;�|��\)�ɤfs�W��276t�M7H�᥌��Prb���T@d�t��� 0� �	q^Y�(��$FHWa%ƃK�M��m�=�׮JM��%�S�
�b�Bւ�C<H�͉ߒ�?w�o��Z�D����ݳs�4� �6'�����[�O#�0��
<�\f��;���Z:-�:�����p�S�+�������t*
-�5%gF�>����+�}���54�ÑH,[�,�`����!@&��p̊��ݻ���ݰ&3,���)�36�
��?�O7%��^{��m��Tۼh��?����/�(�%'��1�RI��$��65��2I2��X7��[Q?�Jz�Ԉwp�V1�D�ssC��_޲���g�r��g8�*��� ���Rc�������(=xT��g��2���IOJ��cǎ��
�&��R�U}]����Ε�ÌT�9h����I�G�rW��~�y�}��f�P��;���)^��J|�(zZ[�jk�*Z���?��D�7<2�2_�=<����h�p�pt47:2�z:����˗���Q4�}��_,��	�cYAE�	'����6 �d�T���-Y��e�X,��q�c�{��_�j8�3��p� ?�㠂����s�(E.�<,ΣӋ��HX`��~�Ƣ�N1��l6[��`���}���߻����]�����\պ��Z/t4z�Փ۶<^�h|�m�O��՗o,f�s�G
��\�؁]J:�qMO"���F���7�8}TQ����l.ŗ���>c�/~�+1|m������е�eK8�óx<sٴ7���^x��+����u]�����?���9v��B�p�����U:�7d�<68����b0��aɆURU��U7��"�JUv �]D�6� e��%u�I�o9жy��C�ExA(+
�`Ƀ�D*h��$��w+0(���ߖn��:�r[s[�D�·|1I�(�d�O�A����E�ċ�ε��Q�A�4��-[���Wu��*�;�zaf:Ű8qj�XCy{���5gyAH~J�\���Ekjj`;-�h�9�<�;��(B�@'9ZX�@�w����o`x$F�,�J��|���I����}���'�G�o|�޽�-m-�n�BF �%u�t�R��H��P��DZՔH�D��?��o�4�~]w��p
�j7�>o������ۇ�?km��HO���G�|6�����2�7$f�w>D錅[n6�ł,�~��x�!���r�]W]��oz䩭��e�ͤ�#�C�uu�M��f>���ڵ�
�,e�V��4������*�*�t
��ͱ�|၇~�4=3���l��_�	ͨ�_<�ʖ�aM���O�^�������M�y��@w�T�oi��fW��1�����]��V�&��~B^�S�?sR#��`��<_,�E��g��p$hcIm��+j�T�Q�e v4Üy��tj��=p^�aiU-��?o{�5;w�*��ҥK�����4g����<�Rz.	·��4���Ԋ�+@Ԟr�)�\�X��ӈ�'�G������W�'gK~_p|4����Vf������K��Y9�������э1/��k��^y~�K�n:�����ҵ��/���3���;�A&�zi�ֳ6��-�����u_z�
�HPu�mٳsǶw\y��S/E�������-}��v��N�)�Ѿ��U�2�Cl�&|� [-H
&��<X��NC��X+X�"��9��,��٤\K1���-�:K-ܹ���(��Q)�@�Ò麊S��F����B��7�Qi�UɓA��T�;�����O�)y������s��X*��P}��tnێ{X�r�X$���|��+/����LnӦ'���%]�����o#��qn(8�zcR<�đBP��lY�R�I{��b��Wu$���;���EH�/��6�(r��5�x�%۶c��Φ������ם�r��{vw������snm%I�$5qO��w�7�byݰ'g�LD�"1�?\M���^w�˗-��=!?e��hUK���$:eŒ��Sr�T<,(x�ʔU�r�����l$�%M��� �])k*�1aYs�)taH��H8�L�M���P����)�d��&q�c�	����k��V�U�ۼ����uk_y�ũ���6n��⸄8�M���S���;g���<zڙ�76�]��3�������RIP�Q��?�>EC���7�/j[a[���K�6��}W�p������Tm��C`'���J_�.h�"����IE��;̡����y`�Rٵk���+_���B�<�79����������l63�u��\�ב(�6��!���>h�� 2�h��O��׿
��r�x��a���\�����T2�u���Dþ�\� �Z*��Z@���_�)�;��bY>�տ�4�6���t��s��+/g���ehko�hm_������ b�5�׮[��������.�bN[���^�����>��G��Ǧ���̍��f�tV�jRs�mk�,�[�y�՟n&��ǒ����-��qL��A�D	6E�^�v���[��e���e�.D�E��+mHt�],��:�Is
Y�����MS�4�P<�캖��+��U�_�����]w�?���w�|�S�?���WA)J^�����s6����MO�ﶿÜ2�`?/ς)�a�듰�IGdT	�D}�[�J��N�<V����"M֚È�:�p�����~��G�\[N'O[u���ݥ�%#QDQ��:T����<)��Q4�G��l��r*�}�n���X�����E��[��Y@a���ه� ;{��5K�����8Z���u�M^���|��!��#��	%�z}>�o��tc�1(B��S�[s7�D���!��t��˾g#�OU�n����?L�}v ���u7��;e����G��)�&O������u���W_�����/_�f{zv�6��r<��Xi���T��=`�j("�;n����z;[n}�;����7w����s��g�Ɯ�od��o���IE���£nS�?3?(�8:���1A y.�fYv.��ַ��~��b�qpp��t ��"tO0���D����ٵ{(�`���H���ƬU>��ްiY���������!��o(�߿������N��>�X[{[ߊ���W����f%��=�y}�S�Pp``�������%� ��q,�s���\&ekj ��H��U=c�x}}Ǣ�w�����撢z%��	k����G>��:;kKe�u��7�\[#x��s���Ce����[�=��&���̏�L�5t��5��(q"�Y� ������_�j����,1I�p��	jϡaE��;_DS�r>;�ET͐YX`!����,w��.��r�\�Q'��j�50�B1Uw��x��������_r�e���fҚp���zI��4�FLM��﯑x�"�j�9)�fi��!ڥqoCSЏ髋*�Oj!˨M�I#N�x�=F�dz�?�)�%Q����2�^y���/<�����o����q�� �2���A��[�v�����MT3�=������,��O����?���p�M4)LX1�LjZ s��T{{��\������])]y�%��d�hz%�}�jY�|abv�$�m�u���L�qb.Vo&��R�k�j4�a.��zvf���R�-(��`�O|�c�O_V֟qZ}mD/�mM�%=�H����,��t���a�575\w�5ǆ�}�5u�w�z�)睲��.&ZH�Մ�c��o��i�e�a��ݵoX_NOt���ĝ��ݻw���EB���[�C��4'r�$��t�{�vI
�>�3'�_�HC�#mñ��eK�J��Mg�[[w�������RX�!��tR4	�B�lc ��I�.�3L�e����9�m�g��= .hV8��󎎎�%}�_~9���b�D�SR����*M�[�Vr~�_����z���uu-�Hޟ/��6�,)]��/������{���y<�� �MZ���f�4�-�Yb����\I��x4�Y�~�A�cS�HDr0"��7� ���J�Pcooco��Ap&����(�"��iZ�	ZP��%)��hq}�M��0,�$�ɷ��+�U�\Uޑ�����T���RC�M0�#�c՛9Q���F�ĥ�8g�(ڠ��YSg��|�������#�#3��+MM��׃�&��{�D��٩T^*�mln��m��CN��w�c)#spƤU�mg��Z��������T�yz�*�uLjKL>��ar���[���L]��k��0����Ox�(��"�o���HT�p..7]�^Y���7T`\GK�'?�a\���������K[[Z������0��]����O}X�LA��:�"�OMMfYlʂ̘�3SCǎ�eXP�K�a��Ѹ�Z`�⇭��kA�S���9ۘ���Ae:Jv
YbL���F���GI�uE1t؎EY���+9X�t`l��}G����mϢ��%=m�-��������EcUo'g)H<:}u������Y�td���W_V(Ɍ��u5�^܂H�܇)+��)�����&��o�T����oS��]s����(9_��k���Z��99>� `��� 0q"hN8�������K��@����~�2l>_V���:�(R�;"������ᡡS�8����Y8��ȡ�s�;��w|�K =�pi���r���#>�<v�{o����L���BE��,����l7x���<R[_��a��:���B`�NLL��i�/��"1��ۚ=za��s�\�I��D�T*�]�@Ӡ�e�;�}G�����XS�ٶ���w��M�Eڤ���iV�@*un�K��Lҷ��� G��@�� ?q�ϓ�%�f����B;�2���~/�Q�Аbt]#���ވ�
B�e�"x���ߢiX4��5�u6�!ޯVY� ¼y�����N �� �K�;�����~�G�w��.u����GǦfu����{e��S�,������ 1f<��M�Y��������c�GF��fsy�;ap;�����Ϊ]������'���2޲��A���
��e��̀E�b��4q&�c"�m6���Ye��g�4ֲu���&lrO$�2����h@&���%Ckom�{�A`.�m�� p�F�_ټ�`�D��R�"+�g�3m-u�fs�:�d�9�B4�3[Ɍ�G���8���ƣ�Mm�e�u����\��:'�h0GS���6l5�y@Wr�7�J�ZA7d�t��ODa����ǎ`��.�O��^N����:3B≥�XF���΢`���
N�®w�oӨ�?��B�v|�T���eW�`VLUU&''��H�����P�h��f�,�&���Vֶ�gB���0�-es9� "c���0��M���&���(����~�D�O/P�M���˳�dY.����E�k���f�LE�}"K��h�R�~�X�P���l)�i�k��O���������L���$v-n����d"�Ы;��޽�������d��������X}[}�ށBA��,����������XZt%c��ܜ*�6z��9�`�tGm~Np�
��O���}�RD��j�b��9�7MYv�-̇:�&%e��9�-�0e�G���{��.L�"ߟ���r���u���K5�#csO?�ҁ��4�
ȁeDL�pF�����Y�l�g�y4w2�ljj*�J��mo�@��|$xb�Ӏ�k�	�R���nB�)�;,��/q��d3�v+��^�LZ.��C�%lRpFhM�`�`>�J��:N���`2S�Ú�r��-Ti�*���q�`��+�C���YV�Zq-/mUX[�/�+>��*�8{�Pr���Cy�����v���q��y:��z���|rnn.�͕��m���Fn����k�}����������|�y��p�k}6�lll��骫�EB����2�ޥ}�#�� ���ʺSՌ[
�E�r���К^�-�Բ�=���U�K떩`3�ry�bm`hjW��@.r�nm�h'[�mP�t�D�B�Pхo�qR��"�6�r��Y�~ࡇW�����b�R�����;x�6�E0�(:��	=�	�n�$S��cy�I��p�-�)����%7�ŋ���J��������E�kj�[6.�����RB�����`Z�!��@����w��EQe�!y�L��������W7mݴ6�{���{��u�!�>p�݈�"�Ⱦc����_���T�8R�LN��iy$]�0�b�����B�^�h�2�%�� �q�[*��&ޝRa��.I?{K!�X�",/�y)��GU{���)J��i�̻�H O񧱘4�&Ho����h�1���D�cU��%c�4(���љl^3QI������Rsi�PϹ����Ѝ�195��e�w��,ni���h��^�4o���ɑa�W^~I>��m�h�bX��EB������u��Զ�^[��#���._�ڦi�a�?�h�K��Tz��=�ML�&Щt�ou���q+�t�u*ݱH�Bn�=��#�A��&N�v��o�b�J�&*wP[�t�U3��W#�y7z�ݿ`�<l�F��8�lDO�%��,��G��W__�b���/�2>��3555`oVa;��*v�����e7���36l���~��>����.g���0Y$�iR���!xs�M #��"K\��qUO�;�%С+z����(B�$����TۣT�'4�X�Q�T���͈��k�D�'Ǜ��;���]�EHM�v�w�����������_�C��wu5��)ܖ��G9�'���$Ӭ0cы�Z��75vvt8|��r<>�R*M�͞u�9�(�ڻ���}�^}%���q�ᣜ�ā�}�/=�;=V,)!Ƭ�l[ҜȌ��|B�c��G�b�T,ȹ|�,�.��{s�7o�O�b��2L���&�t:���˿���t�|��|A~r˳��O�_$���+��ŃY97<>689VД�+;�u1�E"[�8��Q����6v)S\G]X�h��lS�uJ�xU7a�L'+�-W-�ҋ&�Ot�A��BUT����U�jU�Ͱ��C��W�G��x��Zհ�D��R.s��*γ(+ʼ>&���U�`�Ia,��E��s6���8O���(��L:�1��h1��on65A���
\����T.y8$xE�)a�r$��y��#KQ�G�㘂��,nhjQLV���_��-Z�n8Ζm;{׮��K����v%���Ln�G�
�e�t�d��'�\dF*��l���6BD�-H�A����TJΫ��U5lS�������L�J�G��LF6�BMM�����"�%^HtuI��X�������l �S̈́�8i	5�{�ŋ�������;�ZV�s�ݻ�����>_�nCG̉�9��M�nH_h�d�Ҍ���c�)���Ja�sT�p|�l�P�����]*��<KU��$X�kV�u��٠��]��T�oq,tP|��	r���AW��	�7������328���6<<<33C���`�s�NK��2�4�Yq�9Ғ�K�ar�TSS�� m�L��K%Ͷ˺QP��}�L�D���XWϊ���ʊ�A�KO�%w��߽�@MMm![ڳk��ޠ�WHg98��Y�d�,����ٰ{�n�7�ѽ��_����M��zq��M� ���~��%�}G�'':{UEG����iQ��x4	x���,/f~��%a������O}�v1T�ҡ��#�l��Rm<����k|V�.q�bke��!IB'��$Ƅ�].�S�����X���*����O$�t}�6��PU��
�F8Ut��.)���Q�����J�N>�%@�;�˩T�c��S��q܉8��J{Sc�����z��%/?>~��f 7H��Ge�^\�r,C�,�\+������[B���K�&\~�ځ��h<�,jp}M��4&��-�u51��umz��?���h;SR���p��H�G
��M�Jô�rAӕ��:�{���>�4�v`�Xr��01�)�f�k,É"�.�G�<���Ϲ�4I2uC��ŘU���� �J�>D��|����J�I�zc���4q�;n�C��u�2q1s������B%�80A�^��s>�||���g�,�<��U)��������n�l!ϋpH�����̳6�+p)L�縜<�a�D�m�qD�J}d9n�: �-��(t����H'
�'��������:E�į�W�;IY&	G;n�(�y���7'�_2��u\;���t���|��߾��{���A���e�ϋ{��`X��H766vvv>��oAP�y�� �DQ���+��?�����g_���pt���8���
�r����ό��Õkjs���k����@X�!Vo�N+�]���`0�'�T���pA�מ�{�AD������mH�F��-)͋M���B��N��>t$���X���e�V�Z�l8cn~�O}�R�?�������}�\�\(��~?��Zcms4�(;(Ҽ.�}��O�2*,�	�Z��
����mk���L���$Y�ZXÀ�����1�������8�[�jn�q?�޿�f�ܲq��M*`�p�M��$n�W���l˸�FQx�^�������Dat&q[�mM��� n9�����CUm��i��/��?}�szYغ�e�2��i�x��}_�ʗ���р����~���������/��#~�>��l*�ޛo�ynK�J���=�4�>�#Q�K�R��R"��pCc����կ{=�H(�
W�	28�)H�e�d���^|��=]]��hf&��q;!��b�ihBU������¸|lDa��L܊�qKi��"ؕz��4225-+I�$����v�֯�����m�/�����a��]��0�^*�[uh����E��iq"��1��@!�~ÄQ4/�7�a,QS�bJV��N�N�h+�\�9�Z�Ixw�p�%98���<����:�	�*Q���w?�m�IE�g�������ӡ�����#ñ�:77�v��C��\�j��səd2��h]afB/ ��]��v�_N��i,SlX����X]EU3G�h�&�!��>����[�p�_ӔQ�Ύ���HHt��r��$^ 	��/\t�-��MIY��#��`���X����λ������Cùb���T^�;w�Dʛ�Dm}ď�zNeyrtzl`���|Õ�e�7���526�5diTkc#��Y�J�B�}�e7��`�<�Z,E��Sm��~������	^�aXˮ�[��n�����D^T	MN,�����?����x�|Z���X���C;�>�"A5ڢ3�鑡��,h\yF�,z|�'���KU9A
��#�zKcL׌��ᶆ�ν�3#=���s澣CmS�<����+{����ڠdvF�>~�FRqo�ɣ�~�+���k�2�O��b���H�������S�=9�)��l.��ݽ~ݺR�;��=�U]��#�x.�?t���]����-��J{=s[8��8c-���ҕ�^e�**�v���j��,�+V1|�I#�
1�<a�Bu����|��*p����"l)@��4B S��DS��SǓ]�!y<�d2YUU_�؀��������9�����J���uF�b-G��cY��m�]�E�k���4�����.ɪY�I+B*�N��+W��4�c�з��<���A5+���7�{ðߒ���[�P���J�؄O�t����:U+�e�1�hx���A_�r9\>H�JUSi�z���s�̳ς���P׷|�f�6ֲBIN�74�J�G��oÆ �|>Om}�*�&�K����l߹� �$op�����fY<�X�#y�hil
����㑦هG�|��G�y�X��m0�4�8mY6�v�x�~��ώ͢@P:��s ��\���K����x"���Qb�����6���Q�@?����`8���t��-���6�?�����k1��X�`�y�OJ&�|A�ƹ2זUVJ��X[╝WQ��V�θ���gEY*�*q�1�..L�EB��Y��eq� d�g3��[H�p�1bRehPb�~�jD�Z���E�Ь��	���FD��D#n�U�S3��Q�ǂ���r.u�`)��yd�����i%�JrRMs��#�oi���b�T�m��;2;���;�F����_�c�e�o�r�_SW���ʎ�������g���/�hnn.�����'W�X���g�N9���	s����_0d�����q�W���3wz�43�]�lɖ.�����t��H%$�d7}��l�$�dC:!�$��7�m�E�wiz��έ��wF������y�g�E�gF3������y��!��3�x<ދ�j]tEH3��-.#��M��	��@�J�*��
`�oj���P0@��W�n7����{a� �C� fn����0�b�����Xl``��,"�A���ΐ}�Qn��R�L��3Q���ר��l��ajf���^]]C�55�4Ut��<K�ޓda�Et'�r�Ӯ�yE�ˈ�c���Q�TqN�KL�AA���3sg��Y���a��c����A3A�2��P��'Ϥ�v��!�Ʀ�l6&L�kuY�EEQ�F�����͆
���U��p����1�:���hr^[���B�rY�hV�)�A`�@/��`��ʆ`!�p�u��S�<�j���h�g^ ��+���z��W7��.�6Z��ZZ�I���\�c�������|">�H$288��� ��J3<�p!���,�^�=�3���k[B�^q��MƓD"���OXy�9��{��]w=x��`��!�8���r
��Yl�a����,W�Q��ƙ�>�	Q	u�L���%9@^�ٗU��Xb,O%_��� 
b�:Ѣ�rCs��<0�0��o=\���R�e��Ql�[�;���^E�P|��@Y��z�3�$� �����{]V�ko/W�rgS�,E���1f,�Dt��:��}���~;Ӿl��� ��+�CS�����W�����?~�Y^�����e^)$�T����x���FS�c��*�byx���O�uW[������?�䓓�ў����ɉ�D�$�<1ܱ������7����6R�x��M:���Z���%��3�!/��.�Tx�2�(���h�|]���=���6���#���c�GȊ7�xcum��n����FZl�\f� �"[,���oC��ʂ��U��]38�}|C	��P�1mva*����J�ÍWQ����� �eN�3����U�w?P3
]���H��6�f �ͦ�}_������w~�[�sj����Yٯ~�#���諯����-������zˇa�ȹ̃>��l9�e�d2i��0]&y-Nu��	/�����⏙�j�#��Z��{�� mE�W �g��2��p �!3s�â�S*�Kc�o���Q����4#w�k'���&bo��\T0�R����$��6�DM�Q��y(>�N$���Y�J}<V[�066	k�LeQ�gs�\N��~����ѱbeǪ�����q���Y]^Z_Y���fmG��_l�o�bX��v�������L�-[������l}����~����/�r��A8������5��8�^u� D9O�NP���+���Ԯ��	��+�o�����̕W_��$���'�%�����*e	�0O��2�c_ص;O�8� ��{}�\L%(��Ɍ���	��b��(���i�؈Ų·�/6�@�����O-]��64�j�tA���"�H!FP�
�t��D�������w޽�Ƞ��::�:���Ͻb�~�����������������;��b�T�,I٭yB+x����ٸ~p`����]N>�����P˲���k�������j�;X�٩m�����c7G��KK+Id'P]����,6���]���f������DxC���'��'���|'����8)�L�U)W$��J��n�4���U.4��XāI$I��.�e�GG�8 �(�:L 4
&s��#�P�-j&k��g�r�$°V+P�\�֏�[�+e���
�%�Q!��g��f��)����А�=�#�o9m&���l'��,Llx�b�Ck�H1��9�x�;cf�*���:�+��x��ͫ+x��K��}�ӗ\���0��K��L��"�Z��O�_{ݕ��R8��c��La]�.�]�dS�E�58��W�3����tz�X�-���F����l%p�/�Ӷ��nU J��fV7�o���ka�s��}�����_��s�"���L \�(��	�C�*j�?�f��ېh��`^B�UJ�`Mp�&E�%!�sY�wX8M9��s���<�u�V�P- 6:�����\k��ޡï�z���~�ŗ��w2^g㉡��[?���eG��}��K����_������}�k'F�|�Gn���>�}ljj*
���-nw-��������:d��H���{Z뫻��e�ψ��u:�/������%%����_���[�M�h�ۣ�L���S���T�%_�iH���"QX�,QTwD���,��Y���ú��+�b�Y�� N/7D�nX�M_�<aMfV5��͙�K�
ߌJ6����^|	��w~�Hr��G�U�N���P�NO57������O���O�c��b>�O44_iPJ-������y[��#���ё�'�/\�!%�O���u�5W�?a	FW,u���ڕU��ԗs��`8�%�6��,�⢄���\sU�}.A&����Cs/�~����b�%Ae��G�zr���6�/I�-��yUW%�#똭�+��*�:P)�C��+�?���誚�(S�E/����j���Y��vO��#G_���$JK���\���q�x��]��f`{j8na�R8,�'��� !b��� �	((�9�ݠ)�g,��3p.1�^�P5�S��%Ŏ(C��0x���X� D@���lR<:8=��r�d�̬l��[H���=���Kw\t��;.�򵽇V�j�xK�j��VXф.�~�@���6*@ ��Z������:�Q��=0� ��=
��� �[&z����e��WX�8
�b
O�8>P�^�u"85 '8u�{��g�'�z)����a��m��B��QYY%����3���ߔH&+**�'Ƨ�m�׮�����74�l;X)��0ٺu�o��L���+¡���R�G�䩱���x>��lס�,VcH6Zu8>7o�������}�HW���tY�$�ȵ�-�����ùm�y��?p�@E����	�])�KG0�HS�Lғ�>���li��WG���������?��SOHb��	VEJ�Ɔ�s��,qρݏ��N���ؕ}O�i�3�P�-!�����@a�wpruL��D�8.�ҮX�;X�b��-8f�<��B������$�	�O$���9��I��P�1��[_��T�7ܱ����C\��=\����g?vÿ}�ۺ W�<�=G~{7=62�m�"
�L*-E�7nZ�0�nGUMe_�����M믦m��px:��������7�-��+���=����ibߞ��6�GB�c�c�<��vv�Z�o߾���P��O��9��l�TZ+k�����%����_?����o�̧���##c�s	�����p"����b~L�-3�FQH+V�y]*�Ro�q��T*	5f�2�^-��ظ�n ���;�gߦs�����ycq��UW�̉���(��LSO<�p:��#'�<.��p��\�Xp;�"КչE*
��4
���GC��:N wFW
.N�-�Ҥ��:N�F*2�R��q����N��t�4�є�޼B�<n��{���m۸�,+O���~���m�Y?��_~��[^�s`�y�Be^I��,�/���_g��]��i��{<�����b�������u��$Qܽ7�8�1du��R�$��Ӕ��P�DVt*2�+xJ^���&''5%�NƳ� !R���p`s��vG*�j��<k��.IX��`i.'5�$I8q�,���Y��ff�ʎg�z5\R�?�w���<|`ks���ڿw��+v��s9��m���}���-)+���L��U�Z�A	�<�Ϫ���_���o�}���1���[�_׹�n��{�>�''�,c!��!`�Td��;.>����G��c-l��86�*�䦿�������Y�6����pM$<1p����#�O@u���|��Ҭ��C^��(ۥ���Ь��;dV��iw��M� e`��!�r�Bu#�H 3��7;5pa��E�p�3Q�:F��b��n���-+���n8�������`Y0K��x�wOͬll�'�>�颹���(u��fb�x�1�K)9RV���Ǐ��ƒ�e�ۂ%�ё�����GҢ��?����������S[]����~�����O��7����v����)�mmpO>��ζ.<ws��QVJ4�����]]y�v���T(��W^>�?4*�&G�J���0?��n���?���J��$�9$�QF�>yUy�G*++]n�(f30�)X1)�S�N��12<�r{ᘅ��X�$�j�������>$�Īu��<x�s?��ۿ�o_�HJ�K��h_I�䢈8�a>���J\ր�K� $P]����,V\�D����َn����"Dznn��٪�NU8<�A�H�F;٦�����2�4�CE�䉫wnn_U��2I���3�:6����Ȧ����-[�����$f�_�-�ձD�)M��V�d�]�ӓ��5�zx�@Da����U���)_�0� ��=3,�%Oӫ������F"�j����@��g&W|���`>�%#�q����W_|��^x�ί|�� �3S����D"(�T����fklhp{�O>�$@ �
H���q�X����	[��'p����b���Ӌc�������������?L�2�u�y��G]�����`��%�7����s5�4�8�"�a�%���x�ꫯX�Z;;2F�X�b���o׮^py�>�̤��8r�EF�
��r9쌅b4�X����s����K��dsY��l��^]N}�d��/8����G����w,
�[�j��e@p�fǢ��%��%�����V0:�[�Ø�6�p�w�����A������qlI���>��BQ�~+�w�B�9Jq���.�_w����Վ;N�M���+p���r���M�l���j+�**C�(Iwhv�f�҉�i���	�2�IfR2X[���ٴ�&��W�c@T_z������^ ����}骲��K����ګ7������ذ�i��&Mw�'JC������C��u�� ��j�8�5������J.�Ȃ$�%߹r��n�Ɠ���U�	��n:k�u���ǚ��f�@OLLx���T�bcj �����T
�1 T}�2���y��eNsk�E�z����.�'�0�^p(��K
�\���f�&g���y)�N�aY!a�рn�,���4��c�- �G����2�7�D��)6������C�f���%���\8����öD.�o���{aד�'K��鉖k��U���}|t��q����	��G��S�ݛ�J\�8��r,������^R)�W#�R����)��ڬxc	b�-��V�&K�A˨zZӳ<��+���J��19�)-/��ƛG��/_��.�{4M=~�8�.���UTED���_�=�X|�:ߊ�_ݳ��� ;�y���?����`�?7?���sV��vvv�'�[���
'����X�F2zN�*�lA����I�e�ֆ�r'�����hGG��-[���ۛ�KJ�2�$���m:RRv`��D<����3���Zm�K�z ��z<4oɋ��陏��$�NJ`"/ؾ}ٲ���dm�ǳy��es9,M��"�`6�)>��@O}UUMU��fs�+	��[�B�mvptE4p�Z/8��QP�yG˲�63S�T��9�N΄i�1���X����K  �ɤ�ʘ�ƒ�eA�J�8���{3�pJ6�?�����?�i ׍goZ�n#�ga+������g���{l��׿P&������wՠ�bR���(�(Z0��id'�SV.������5u����6ư��Jׅ#�ϮQ#!d(^z���{﫬�޲e˲e-�?~���-_>��3��_����վ��-���r#��+e��V��	�хx*131
,XW^Rp�H���F�m38)8vܶ��EI�Q�	TK�N�\�P��c�5�t:]N��Y
���YC�R�!e����۬��,���V�J�f�����
�1�ȑ.��Sa2d.��'�l5�0T�rf1(�Ld�
�ҙ�a�����ڱ�����܌��68mcPR�MFe8
yzM1`V�j�xk4�0hjj�w���|�G^߻7\�=k���l4�.9��u����.7��e�H��%y��P�l�mo/�_�Q�-CbFTA�a����¿{,2�w~ٔ�&M='��P '���`櫨XG�u�`#�1�U��,Ϣl��_~����6�'3>���_�ޓ�>x�wn�&c�;Wj'F`�yC�О^u����Q%�Q B�q��(���y�g{N���p����vS�����ܜ'����������p�+�k� ����>�����R�,�6���$c�6�5�]M�o������A�ܟ��m`Y�۸�,]1�&қ�� �(�B��S�4몁|8�N����wnn�!����K.��?8�����~���$C�#O=��e��Of�Q1���g������yrfn�e��<�� 	*	_*�y]0
(�ﯨ�R5�ל6wya�'��g
�i`L("~h =0ɟ$J�۶�b}=.���P�ꢋF͔M	���p?��[^:t�+T�S��u�������e�+"��Od�9 [^?���V��V��E�
o�'�(K��0<J������������Mw��r���_��J&�<�p���d��r;w�|���3��g?s{*�y�ɧ��𫯾��}xrrz��/�\�2�M_͕�����'{CN��r0v��c���������B"~����$�tLZT.��Z0:\8�(�L�����h�X�g�+���������f��j�f	%63�}h����hi(|�9ʼ|b6�i|
i�&�,�^���FɊ�r�O����|k[m&�Ke3��p�'*O�qb0BR�,������b���/���?g�\x57\d�S5�f��Q$��j��T�'e�k��JAU5(���,43?���]q10Tt� �j��b�޼�a�i���I腲��i�����<����q���{(e�8���Y��!�:���� e���gE^��l$\����3�ly�m��/t�v6����������9�7}�CSs��AX�#��'$��������`���nQ�,Vvdtxjj
KY��fvt,�m�h<��~cv��A
�J�Mcq���ҼTe -����P(�e��?44bsح��وo٤g��H�X"B���` ��ǁIEQQ1��5!)홙V = �Qس`��������sι�˫�)�'?����X�|�'�;q��q%/����~��������x"���02��x����,s��Q�/000��4�[UPk8geA2p�(]��P�bCF)�,�Ա9�,f��L�����B�e]��nw�E���5�񎎎�)SG*ے���P$2�$��B�Z�)�LѦ�J.�)SQ�T#�gd���V��Dl�����.I����z.��F7;I�� ��	�ǋ�|$�++[��`��#sY�*���$	x�$�Q��EGO�t�E����yC>K*��g�,�-_V���*����L�H�c��L����t�"/'��I���$D����K#�����-v��������k�o����, ��낟Pi��"�K:����M�@87;(����#�����A��dsm�k��Oj��rV�f���|���2:�4kp��������6�7��e�]y��\VT��X���w�y[a�-����嗫���{��k��.g.�J�l;�r�x\O����6���e�u��낓����9Dm�K1��%����"xK ��E���p��W�d
I���)XB�䒬�BPc���yaa�/^������g�2� ������r�Q�DQ���
�D��v��k����;���+�~��ٙ�_?�(���Pe�?��^}m��\|fd���J˫*j�/�o����3��#<`�1�҄\~Pr˂Y����mv�Sx��,��	��i��D�}�f'p�%d�����644���ͫV�±D��2�u	S�w�S_�m&�.���u�K�rN�)�e���X�kGb�`�e�eክX��"ȹ�C*����ˇ�v�6חEB[��?35�$���mO�8a���9K&'2���fs�,o���58���@�z��q�B]�E�*��h�;�����r��^ �p0�n����*��������{5��#1R,Cf�<�Ł?N�Y�,�zyYp:�������*�,�T���=��A��ͺ�=�#"��͂
��b谧$�ݺ������DQ�c�Y�g)Ҏ��CE@\�MC��z����x\��}�oٲ�־ 7E��eV���3��uק>����x϶-�*B��4�\A{i��7��w@�Ȃy��jji�5/��C�p����<L�t&Ǡp1��slY0P�-v����$S��f�`0��{A�՚��6�VuW(�$4�R��cc]-N�2�/�fL�X�R��0R�LEE��͛���bT �vG6���6oZnͫ����חL&=H����yXu	,��n��m7�|��6�������,�����T	uŤ�t1Q��q�@���qlRG��\*�Y���h��0�֩�ץ�j�8��$vK��8� �?b͉�0l*)�$���>./��䑇vjď~��ޞ�m[+y7�rE�F���ǟ���8�扮�~��74�{|^�RcS����K/�ֿ�J���<XbK|�sL<�(+M3�����
��<\WW�#�H 
*jm_%Ұr�?�Q��۷o�?����f���9�@$R^�I�ׇ���Y l���!QP�Di��G���fM��2�^<$��m��g�ȁ30���W�������k=nJ���ږ�� ���3���l�Y]6�w�@�m6��Pov�L�!�jY h�%Z5Pֻ��o�80�Kq8�Ըҋ]U�y�8���*+��h���6z�N"5U�x��h3�g�"	�j����pB�l�G�����q�I!DQsîe���'��R�@"s�o�U���WF���#�����������妆���yl||����iI����o뫪�������.��h䟘�TE�q,�ɨ^ִ�|��u�M ������#k׮�x���>q�m�l�&JJ#�#V �TYW����d��}�W���3��7���r,��ēpw�.�ژH��e�Xڗ/S��)��i|���'r9)���Z
���h��g�GcW(
5D9)�\����;(�͘J�x`%䀑K���������dS@=�C8�
���ኄBU5u$�M���v����x�ۍ�-��T�I�X����c�%ʥ	��be{zzz�2oH�K�:����W�d�Q�1�XE�TY�ڔ!H��� a����p5=I��v)��f��(>]�{;���԰��8��j,� ��R�9s��;�ۤ�h^jO=�d�$82>ZR�	Í|��#�l����z�Сщa��KJ}��
�s��Ej[[[)]T	2'+U�c�ݞ印0���lf~�����p8x��O��5��`Չ���Ah��
���JX����ydY��1�#��w~��n��N���'��PALq&��QHd ��[W�2�J�"��vWa��*e�0�L����꤀��2-j�Uu/������w�qǎKv��M-6m�鋗�}�-��gE�b�q��l4մb���x\H89��x���yE"��d6�Beޒ���H(����@���t'z1�����zPK���-�:V�U!/G�����vP��d��g�WP��5T,�+�������ʺ`���js��9�K�t��>��މ���7,�𺉜�0��o]�j�ݹlpp0�Ƽ��^��ǉ��!͠+��.��J�ͱ�uE�Q?X0�r������G2���a�9��;�����N���};o��׿f�9~��;V�^��\�����^�-�����t&��ިHƱ�#�u��R���X�Y-��id2����<��c����m�Z�VD E@
���LNp��*4ͱXx��GX[.i4G�3�A�g�8�":��8ඈ�hP< ���z ��LR�������c�M�z���5�[i�5_�:�Jb�{��}x���<`3��}��#����i�������ռN��/���}��3��a����&>��2���XJ�:�B5�HאNG�3T��,E0�a.:�,���#F"�h6Z-6Y0�,t�C�d��(�=�j��g��]��c�bdo�G���`bdFp��4�b!u%�XW��T*��ӟ������%����p��ov8��o�Zy8r�D?�ЫV���3O��C��ߞ�',���P�%����@󌩨XV��/QT��@�jk��W��q�!�6�wuiiis(�������f3��n߻w��᜚��'�$p�Ͻ���;�oۺ�ݻ�*+q�Ǌ��F:$��H��J�,n��̻�T�lc�s�K�5q/��&�2���鲢J=]�p�K���O<�����&��}�����W��8q��w_��뚛�"�b�:ٰ9�v����6���(b*��0��G-N%�<U�UU�<����R���D�P?���8$g�B��������Q�㣛�6���ك%���fX�@��tCj�ZY���E�5�Q�^�2ꝋ�O}lQ\T]���ޭ��B��c},k�>q|�W'''�++�v��r�t��}MW����؉� ��u�UUU�ůd���t.�M��Y�z�����U�ǅ{]�p1&If*�܀� a�t�f@��k�˿���<�s2
���r�����=��"Vgi�+�����l�]�ss�&G�[�����{��_��������o}�[��W���}g�_K���������pD�t����*K A������w(`���NЄ�'0�Cee�����Ff&��h�@SȤR啡�`�vp��`�O`�H<cv�(N<�

w~�� L��w><h�Y�eO"iٚ�:����/~9#�jj���w<���b���GҺL>��`r���<�ȣSɀ�;��^i9eSr9���r���T�,l&��҂����4�E���yF�z�N��9ppP��B�Da�*�^�6;�P�'��)��A�H|��t���QU�Td��Ϳ��Bf���;�ʽw���O������	S����b��:XF�|Vg��
|�?����>};�Ȋ$����7�.d�M�.�������O|�����Ѯ�����X���P����Ww,��ɀߕ�F��J(M�3����9�d2f��[M͍�N�P����y���r���fA��rb"��Xy�>l<�ĩ�s���#�p��[ ��D���o���b�4[h�G*��Ð�aE��x�۞j�.iETI��P�'�_(�tj��d�3�aP(�HZ+�+��g�z����>K��gn�-\�t������q��WL9��u��Y��̤�᷻]�c��uU�\~��7���)���dII�K4!�t��.%��zQa�T�R,,VJ�~՗<6���)L�P~ ��8Z4]l*{��3ګ2PP:��cG���� �D��p��oM�5,,�!>�p�7o���s��]rI�矚��7T)�N99gkg����P.���c��e��tii��+�޴�%67���}�_���^Rż�BC��,L�5��������F�T��N��WYZ��'.:k�����z�#A�&��a�����[�_mzj
>�zd�gi݆����9Iy�z0qd��u���˫� ��|.]����� Nn��l�A�ӹ�G�I���^��S�٨882J�J]E��Sy���w�!��`U�`8G���l����J�2���^��a
;��cpn����� �\N����(csee�l�ؼ� ��XBo���u���xZ
�X}!�a�X�+��_�u������s�6�HeH�y��z�S�Xך.dr^_�v"�v;8;cA�� ���k�H��݉��^	�g��1(�*47����Q�X�	��[6�𡿌��546T�}`�k.��O�������ȁ=��J�^B�}L����`ճV.{�e㺙�I)}��'I+�b~bV(J���dS���DB�
�(E"U�o46�l�����Bep�;�W�Lύ�M �K�P�z0���;���� ��AS���:�����^(����i
����<��*�� ئ�$1����m��$*�R,��T�#�����Z1�4<#Χ�A�'[�����q���W^]�^oaؑ�ټ,�jk���,��F�������h=�M66W˲�ц��C�=8M�.��ɍpF��	�l;��I.&M�oK�;u�uj�Ǡ0��h0A,n�W�zL���,4��-R̓T�bG媎�lP�������� ֊�bƆ�����w���IBea�����j��s|�����_w����W�S�V��f	��.-!�+���h�?|�\-J25!t㺡�Qf�F}I�F��< �4�iP�) ���X8�L6��I��5v��wXp�v�Y��ufz���[�����P6JmM��Pi|a&�� PRj>�I-�^�F��RUS���T�I�;^�w`�s/�X�Z��g_9p�U�y��'�)/-}�G��0Z��츀�a�u��N���X�G1O<���x��ѭ!��K�(�ʠ�V��� �F5������DJTm�f�������^���"VJ`ݨB�$/b׮]�`X�d�*���,��uk�az�y��#����l��������E;v�5W�,19o�u�=^��7?p�W��(f��u�A�������˗{�v�l��Y+x理�����I�#�����7� �?h���*K���O|�f�?`�����O�zΚS6t��Fc��_��9��_��Gf&�����G��& �Um͵�?����XYYija���Z���ƾ=`L�lJ\b}fhxll|ɭ�R"����\&#)JMm�c�=+6�b��KJJ�u��N��(�͢�L���
���驚�����ZG�
�!�N�2�6�K_�C7��*��:��I�i�#޹�fc���@��9����$��M�8�ZH E�i�Sу���nll$��S�������D���u���ڵ���9�L�����y�����vS_]��zN��������>�un>E���'�,��ӻTڙȪ>d�4�47)u�<^�|A��S�o��K^5;�.)�/d��
፥Y�n`�6Q
���"�:�����,n_��Dζ�n��F744��� �����K6[Z�K�����T<�%J��n�1ND�8�Ѥ�#J�\7}���o����5�K�	�-�����/��@��1Y��	H�t�I�]'�S6|꺭jo�e��d<�w�����m�Ӥ��g���Ғ�!o�4 �L�����j!��Jhn.��Vp,EQ����}��._����Ѹ�C�����?����j�{�s'��j����ô��׿륺ԥ�)�(d�,^�F2XV0G�� ���(�?<�[X1� R�$�ͣ�BcA ���,%Y8�X�w��\++K��)8y4y��
puw�?����γxY3��*�D���X,��ՕF-��͢\�`0V������÷�VZ�~�g�«�o�]w�����o���-�{,�}|h㦭!�(���������3@���J�4��ve3(�`���(AZ��v�� �A'/��~��?�C�V����-J����}㫩�\&6`�I��Tt�c(��&*�I�e��|�X|f6ZQQ
��n�K��v16�A�(M�>z�j#$�@��efz&���]s8l`Ԣ�(,�����$Tٴqc6�y�С-[��MN�6�MMMWUD&��+�m��6����F�==;c��Ƨ&k�&'�:��>�ԳÃc��r{9�������<:::�/���t��?�)jY��e�44���5Ծb�M7�6d��r���|x��&O46�����m����#�me�}���޿[R�K/������*���f�^��%#K�v�N�QK��A��u�UpQfC��1�	����)Ќ�1�ys������1��@�v]��t�R�&X�
�Ն���Yݴ�Z�6oEMz��\tA|a��ښ�ӟj*��{O>���U+���=��������<�u+Zn�l���L������J���~����ёk:N)5�fEAA0�p�f˔"����
�Ŧ��؂����>�i̠��$u����On����@ocmE"��J��������ܭ�#G�TVU�s��p�+ږ!WL��p���@sC=��B�.���d_�IU�5\��(��EG��@-ܽ��_����e�bN�S�L��9��`Cee��;xΖ�,,��#�5�7�N�&�Y�@����5���B��c�D�1aw�$��`���,)	�,�f��Aђ�XSU��6��,K����[�p)��)�ba�ё�g�aq���?8�_R�����pmյ���{���rZ"}�8~�m��K�ș�IǪ����;�~�L�8�;z��7h,)(�B�+�e�?<�ׯ5~X�\I��hҪq�b䔤C!�� Xj
ʠ�'f[��,�^g��2t� H��;p���y&1���?S�mPrm�%u��F�Y
�P�W����F���y�ӏ>|xvvn��<��S��3**�5�<g��f����G{����y>�H&Qz$M�J%SB�
�G]W�h�q �h4��vX�f;�֖60a��������GFG3����/�'�'N������8�J6���748����B>6"3;�[��|C�5a�!;�%�������]�L�����GgF���9)g5bx:�s��}��?b�<�듓ӳI�K_����Dg��a�zbb|rzF��^�#�=����~c�.[t٪���oTW���>�i���l�K6l,�y7a��i���^CB!f#�l@�w�\
�53�0��\V�#Y��5��e��X���f�3lGUA5/5I2��U<�rCsO�$Y�����L5(�QK�Z�� � ���g㦍�GO��IBP������Q�Iº�v�o[,F��;|�?�s>�̳`g�D�`�����{�/p;�5��X������Z�D%�^�Eȣ�KYJ����5�Q�xI�r��w�����c]G����xב��1:اHy Ocp5�����oȪ.�53�:���ȣ��������yQV����4�<����G�I��,E2����v�Y-c
�9\��<  ����V.������xt��"R�#��Ã��uUv)�C����gG�e�bp!�2�×���j�a��*B/H� �I�g�ưL&��WQ%��ZZ��^? ��j�	ڊ�UŀU�����8u�Qݍ����cǟ|������6������f�J�,B������C�P��약���?���j��肢 U����o���=Mu�ç%�q( d�>�/ͅ>3�3@�.�������Q�4*�9�hѡ��'����sQ'O��ZH:X^�Ee@]u���?��ݖ斌�>�s����ri��!
"*�p��B%���}}�`+�Fx���k�e��ь���55���5ؐbXXkII �w�!�.���oݺ%������JAJ���>>��g?{mGeMEo�`ˊ��.KVOɩXtnd�G%5<W.m�<+K��TB����WP;:ՐUc�ڳ��Z����B5�����X�?��w�b�C���p8L�5k�>r���Z7�$j˭�|��e4E�Z��'�v.R�c��U��P��vY��3�N;��Y���9d����6[�sx���
�<&dZ!,�!^Pl���C�f���:* 0����QhJ�Z� Ώr�P��2g����d,O�]^�bC��0p�撰$�&`Ӂ����< C��.GII钾��;fg�s9��{^R��4�0w�丷�rlx��vt�Y�J��o���'��Ibx��giE��sc�C �(7�xKx������o�D.J�v'g�U5��f�r��g�E���:K���;E�XnrjF�V�q:TCa(ԉ058�t9-V��KL��$�e�3���V�Z�����p���Ĝ���	�`RCZ�"/�sRV�0>�������%1Gr���T��=�?����?���\|���(�:ў<�Zu�}�b>D���$�E�輪*+	\Ĳh?8�M%z^���5UU��'rn�3R^��zE1/�*Q(�r��ɉ��\[SMSŞk�㒋vZ�$�<��뇏9涵��;���V��������ڍ���n?p�;�S_U��E"�Z�Dr~���������_����������\r��l�>-�sP����B����������Ô�}73E�^6ne^P�CՒ��t���Z"�����������Z,���z{O�O�_t��H8&��/����/���Z
+�� ���F�F��cI���9���gvnv�`b|�����H}C�k��l����h4���<yR��2ɡ=������ֺ���g=�� AXY�˦S,�i2��g�3���k��!ks}�F�Gq%���b�����ʫ���H&�P�<�4���׮^���㉇8qb�����%|,�n����7?��=�S�cnfJɋ�5/d�L\�����tyI��B�f>r�m;w�U��&�8�Ym��Ơ|M�ځ��suC�
*Q[645�65Q<SC}�4�X]%Z3hU'q�R.,C�R�(��H+�P����@`@iTA���Ψ>јI����0V�n�+�&���S��,`<:�"@���^����ٰ�t�.�q�K���s�p8��m�\�wd�Kf���r-���:|��ͼ���-n�%�H��q�ٛ�{��_��gB6�iuo����`a�.q�p���O?}���B������#������?02Z���s�%��X�,����d]U9�3U���G��4����ٜz�'���Lmm-\ɖ�F�  -��	�1����h��D�#/�~Ғ"�a�zY8���f���� F���-L�����%�#����K���a��m�Ot���^���$��U\{X�W'`� Έ�X��x,���0(˕c�������s$7���DY�����Y���,6�2Y��(�Q}���ظe&��W�<w���WӪ������9�:��_��}᳷:���x�8�?�uq׭�ݽ\��~��;9���D�i�i��.�V�U��\{�]�-/+E��:�v�s�N�Q|�xW����q��X*��jup�dnn���l�I�?e"���6o���-�8}.�?'�7�XU��0�(I� j��{a�M��\__oqX��,+-�[��,���M�Tna!VSYױ��,X>11>>>���7���ٹv�ڍ����tvdziG���c����܌��StU� 55��c=}�_��W�ng&��=�xt�2R�ٹ��{3Y�4�n{Ɋ�ҁ��e��kwܼgߞƒ�'=�\��������YӼ����쮻�����ba*���)�]�|CMUG[���|�,�3�-���Rc#l.j��sz�;��mp֑H���5�\ٱ,��UW�Sy������Eѹ�5�U�-�T�,�q�#�!��Um����e'G}%.w]8�ۼ��4��e�q�D��u�艖��bi⍓���{cld����};/,�X��R� J��!��/@Y��&;�>PH����*f����F&��E�OՁs�Eah��p��p7����>+�&�j�ON(R쩘��N�Ɂ��W^߸z�j�ϛ�e=/5�P��:2>�zY����55����۾qz!
7tz|���#}=mMM���{~����w������p-��#�s�,4�M�"�k��;���d�NO?�ӛ�py����&㱉�������uv~*	��a�3����>Ҕ�Ҳ�0����391�Ɋ�@T��N}NTp���T��jE!��	�eG�%p:y]W$!�F�N�O#	-/Z���**
ūO��?��k�JU&uTd.�$n�aꜛ�ڭ�WX���o_����B6��6o�\�`0�M'}o"c�<R�u䍑�Y���K}~���\2���KKqކ��P���"IKp7)�����f�9o�
���+��U���/8��v���_����~{��Иlg5˳ҭG��Uu����ĩ^���xoh������(���7��k�SKz�G!.�X��a�@�TE������
TPh��Ƀ�F���K��{b�����v3D���-���<��I�H"���A�0{��F!M5 )�`�bv�^�4C��\��lA
�*EU�ր˹��"�Æ�-���rN౐�YX����KJJK����R)�C�OaM:=������{_�/JRii)@|�$����.<`5}>��c��֯_E��P���6�U���JK�<8����xye� >'�۝��U4O�Ҹ2������9�!n�\�98���L�TYV�	�^��ʮ]�/ڮeSM��Ĝ�qM�]w����/�x�<�,�q�_���+�R_SWS���Kv �Bm_�p�I��v����h>7y�I���ۼIr��Z�\�(�ֵ�ɭ+��(������6Dy���̨R5����?�|��J��C<G�̮W�l8o��7]/�v"��_���O�R�R�� O�X��Z�����1�䥴�F;�.T�g�XXJC�g�v�jEF����gi����/�n;ES��p�*J�8��O��4۴jeTH�[�x$e�F*�Z����Չ�]�|��[WF�^�x���?y����R� F@��A8Y:�?��sϹk:�Y�� �S��$�h ���dΧ)8N���ļ���K�����}>�׿��۷��ץ����E�����VM���$�m���Ȳ���`�Φs�v��!N�G"��p�L��<o���gf����)ݬ�P5�~�N�뚵�������II��b18咀jz
�1���������.,, (��T*C"���f:�������j�ͮ�����$ɀ�6�&I؄l6���E[���k�	��6w>.�9ٛ���a�	�9�ߛKghƊ�p̜U�����+v����Q҉�tM�����Vⶾ���N!��O���4\����Z�7�x�[4�=6� �K�IR4h��j=�U�k`F�L�~�`h�E6%�pn"ŘƢ�&�'�/u�%���`1�:Stz}n��W�L}S��b�f���������c��䨮�����9wOO�A�Q�I		�9�l����zwY{��w���6�	c�$"#��(�49���]9|�V���^����������Luխ{�s�{�y�<b�4���Z&�9��	�480(��H���(Ȓ��h�����x*��p�v�/�sM&�H�%������1w����c2�cSIï��Ɓ��e�Kztj��m��×���G���tc}���p�<B��Yib�N��x͍7^�q"� 4�"����Q��S��]�pڊ�k6��~@t7gs2������Si�.ɰ�4��<,J �I,�J�+\{�����2���H�}IE@{m6����:�ȇ�)8��t3K�E ���c$�VY
~�)�@,DM��=MՍ�׶�-jĦ�>�Ȥ����t��%@&�2��T��(TI�㴃SĂa���E��S�H��jP
���Ɔ���03j˃
��rBb*/J|Ks�*ɲ�Ԃ4�'Ck�aP�I�k�,~��?f���##�����d��6�oߡϮݸ�yAuM9̳�!�W^��3��2���_�`d<w���s����/�G�<�ğ�uXy$��"$�Î�?f�D*ˋ2`F�
��:p���c=�֝�⌆1����/0�����G��z��
��V=����Q�����6�hV��2B���5��UU�P*�G���ʏ�]k��|�s� �O<O&�~���j	�CH� ßJM�$������\�Dj(|�������=���l\��� ~����=:>6���G���DFư�`p����נ�S�4(:�Y�H0�2���0V�����٬�hJ>����3CG\~�n�<�i�Sa�
|�����i����\)�a�=�U`&&�oO�D#m�>^�J�Z�ޚ (5���`�?y|
��aƓ�'e�=��Tf���,ЛC�#��d�(+�4�=�DnA�Po�6oެ'=3`c��ɮX��8��V�TOMM�&TE��ұh�{&�Me3B��B ���C�GPɄ�+�hw�s8���6>9><<<15�`��;v(�FR�,˰�ഓS��U��|��q��X,�����r8-�du]����m۱�M��kk�,�y�x��d��8gw�Tu�ܱDa�Y�>��c�]E{9���T���PE� �n��)
D��ǒ(Y����/ȼ����.3c��f�YU|�����TY$�د,�ˁ�������޺U+t�U]d0��{��q;]��.���΃@4�.zwF'<ွ�"��ܛ��6�ɉ6�`hǝ��ʁ��tw������գ/���'��s;FF�~���
�ȸ��;6^��/mz����>p�@��؊��+8�1��xW������ ���� N[���MMO����3�7³H'S|.����ۊD ^�ʢ�T���C�G����~��{����z���8sƋT^���I�D6/D��%���T;�.�YW[Q�g�A�в(Yfq�-�F��M���ƌY�O�NP�l��e	����~�ǁ���W�SEgdI7K!5-m3R��JS4����3-<u��dU��;�*q�o�G>�)��憙?&�p�N���Q�I������M%;�����k��1}&˩t!%�q)��X�N�������/䜜���M��qv�n��$v�곆��ww��a�+���o��bQ��� v���F�届�w��Y��K��� b8�Q[e���;h�UEi0K�`�?>�t:�n����S�=8V,<N��|p�H��"�f#hYV,���W6K�]���Ju�!4J���6�>�|�ԇ�u�>>¿�@�',;����#L�x�@��ġ���o~��}�(���]�Mo��e|d�ewF�ᆺ��[��\����y��hȶ��|:>
�.��56��3���ڹ�����6�dM&����B��
�3Oo�d�{E�k�� �qR;�/�����ov�ƭ[�mim��
�T&�)�郕�s�a����ز����ー ��d��ᑪ�ڪ��/��ٲe�(e�eťK��Ȣl����olQt�I�����IlE�7�Ǻ�}+�5�146�G��3ʫ����E0K��E��*��`�5L�a�L�4�ʀݱ��i�%�c�����Du{�L���6p0+���¼�c{��?{U��~4��6�|/<��wO.WC����Ω5����ӯ�h�N��Pdpd�s���q�С���\C>Ut:�"�n���5�V5�s�������_�v:�:��3;���lz����t�U4������8v=���:������ot�����-�'��_�u ���x�װy*�y�{q{̧�[?w͹?���e��T�z[�|y���Հ�]R[I��X���~g��Ռ�-`
/����59�t"!:=��V.�P��<0:Tw k��l �JN3��
d�%1 SZ���ʹ�(�C�d��'�I���>�?:h���? ��=w�#���H��Ydq��+�1��CIh&54K~΄��ter�@n�C=x!X;�婆�����㿆���Py����kA�0���ө������/]���t��������q��B.�p�ٌ�a�Py��-���:f���4��D���]�e3�#��Yv�����e�_��W�ޱ���7'7������`1��J5�����ښ�?�������������g�#{�f��!�fr)`	KR�T�h_  쒦�t�h.�z)�c.�?>-��,����\���X)�݅����^���-*[4���Gܔ�B�$1m��P�Z��G��?	!�O��o?H�0�V�Q�\N�EÉDQ<s�%7�pQ<�>��L�"v�_*���w��_u����w��ȑ�a ar`~�w۶�:�&��`���Kw�F9�W� �`C���w�y;��@8�l�b0o���njh�O����MML�]S�U{��ٴ����v@k�W�wI��^����	���"�Ę�����.Z2�s����ўs8���ﾷy��������ʝ��'�)�\��rc��c���KA\�2�K�W�_�����u4a�㘬!�Ѕ�Sp��D�5�Dk�L91���А�
�2��ui@��ȃU�R��Yr2�y���v�4��R+�bB��Eq�(Ѽ��M����� d���p�(0���]&78�!sz����v��؁m�WlX�7\���w�f~:�ty]��M���. �[��9N˩�.�s�i�?%S�5�	UN)/J a�'��|��Vu���G�N�Z�k:��/W���"\J�t��LiCdt��ȱ3Α���м�j>�X�Z�� 3tV�T���<%� �
p``�3���K̔K����n��8�q���1J����Pt���}��U{��p���q`��P �t�lf���b�����=�LQL9��&��?bK�m�I�,�G�GFG��d1$Kd:�����N��,5��OV)ݠU]�-����gb7M%'�4ù��J:�~oO�����g�:��ڕ�c���Fo颎ƚ��t�c�3i��4ut��[(�~��r�}^MQ8�mdh�LqCQRQ=��wNNf�`"� ag����Ww��9��;��s:�c��cSu,Wȳ��D|�Ym�����]}&E����qKRM�TSXmV��g���>�gv>��]�d���`��9{�U)kVҟ����:���S �f9�����emF��导��g,���i��k�E{e�+s�,?��fI���>48���eN.3Ɛ)���DfbHd�P�b��T��T�"����r&R��B>�����i[�ti,V�J2���qEӽϒe�k���ٌ�ƹ�n��Ų�l6G(f��b{z�8�d6_ljmj�3 ���:��(+/_�����2�|U]��S�٪�p'9%T^E��y�*��|l����zw[Gp�N,�<����ܦ����-IT$���cT��⺂�����ڌ ����z�T�9�q����$�1!;�s`:�h\ʍ
���$[dr�d!�'0���`��" �
�0���:Y kk^�p)�h��nC(bt���n��KԔ���OM�ݘ�u�x��C{�;���Sq�`�U�ُ�(J"5YT�p��v�?�V�p����p��tL��"�6_�	`}�ݻތ��6���͏��W]���%�n
m+�FQ�j����>��[�͛[=V,��Z�e<�P�sN��􍌉F,��"�Q*ʾ�	����͗Ҏ�[0Z���l�bs�Z_|��w�#W��K.��c���cөĢ��A/@���d�Ҫ�;��`�Y�$�ӯ����%���H�p�tլV?�����C Z�,f��Ç���(��.���F=�4Sm�,�&T��O%��Amtr4BP6��wpl<Q,��T���#O����<��g�k)w���N,�|�b�>�{>I�@G�6�VV�dҚ�14��m4E��>�XL�՗^y<�CG���A�����Űd�z]������]��~�w4V��X��n��l���hkkEb��*L�;�f�0k�/�����\�\���?��Ք29�Y�Z�vL�$�|R��E)��jA���3�'�������Ɵ���)�a��4�Z�����LjSMm��8������$��;�ԡq����՗6��+���H�����.���Q�������{��BNPQ
��jǺ{�,Y�/H�\s�������0C�ON���_xe~Ǽ@ �ڊr�(����(nAQ4���v�~~<��=66�)���bckۦ^F@��rNG*����������w9⍔˪t��t fN�a�C�/}�ۍ�[�|���N3�_��W��{�b�"v5|��K�Ϛ��L�Vx���,������B|V�56�5�����GOs+�@7P��ѩ��h���/r��n/jB����"x1���A�
�N����J��MU�"�#xj�AJ:����ʪ8���`�O���Y��N��_+��nkcȞ�Q8RQW���%��M B��ed8�-�\������$`�|��`|�P���T����bK,�|��s�.�U��ͥITw������4�#�g�L  Bey�q�
٧�{��������\y�剩������"����W<��S���A��ukۛ�[[�P�A�hr��ٶQvť�w���@F3����#�-�b�U��&�Cl4��@��PW���!�?�p(�c�����f��&�>���	<��{�Ca¬ރ�%1��s��ػ����v��Jp54S�+s�(J���֗^z�{;v-Y~���ĄW�dEDb��~Z8���q��Ͻq���H~�����!��788���K�g�/�ɱR��?�ۗ�Osv�8`ư"e�>���W�,�������`��P2��6�&,�y��`xtt��6	�PUݐ�ł��Z��k:��"��f�y�Ң�fWQ����jP͔��	8��-(���5�� ����v%1SG��YE�P�Qb������R�Oخ��ƌ��@�����#�O�����������`���@U[}Y���~�Y]��7��7lX7:���:��+/_pᆡ���7�u��T�u5��&�f�t����'��r�H$���x���֬��s�Ѩ��.�|___sc#,<��UTTQ�mxp������6>���)�I�TI����LK4�E�b��|���M��h�f����|<����D/=EV5w TS��	D|��4/��s�ﾝ@f����߷m���o���?w����Bb`������ښt!�F5C�������x�y�@meUc��qf*͢Ư��*��@l�v�ɞM�����`��J�l���-��ًcr8�2S�,�f]>$e��fҩI-_s�/�.�F�~��(��2�5�@����U��]q�U�V��26����;n9�k��KMH��,�����@�슄�Qe�32��2�N��Z��9�p���?�3������`;��.䊤�ػ�/K:���'MH�$�`�. �e�d�I�J�P ����/��L{~󛻷�U�_r�eN��_���������)�t���ZZ��*U����F�V�`�XoYn�ev������ps^��4i.�܄�ZȒ���4WUS�Dgmd�,������A�3 �Z��=r�{t*�`��DW�9s�M/���#�"�tuommx�����TVW �B�l!�KK��0Q�9�8�+��������{�F�fCA5E�(����ON&����x�u��t�4y��z���R��/06������ ��B>��.�Y���sx �{{ԙ�s���lN�$����ޯ+�t(J ���Z��H��)�%��X���V1�����R�(�R锃������,aw�Z�n���h��
<��m��6��ONcj6[��$U�g}��@�H1��P	A0��v���jZ=���|}�Z�3�IA�O���9��Sg���JZk�/w���v\쌕����¦go���ۘ����7_�h��t�BXe�:w0�v9iOD�e�C��|���e�P8�T��GcU^��yQ⋅BMm��nON����/�������*�I�L$5�l�n����s�[�xQ�6�`s��t��^�!םw>|�=>���o���WTTt��C����H���ݬ�WsI���ժ�p2=��'�p2~;ㆥt��u�����5����7~���/粅'�6�p�5�M����J����x	���/���|u3eצa���,�&KҪ,=��T�����Aá���=��LO0##b��`�qY)*����v�Acf�7��J�t<)E�.�ؖ���M%��L��<�5j���ښ��u�9�32:du�Gi�ބ;/�Y�A��".kv��u��.�]ҁI�0C8[4Dxg�z�܋�M2�����;p�E�?�"
�h�!i�H���X���U76P$V��NY���q��\{�������r��S|�/����(F�D`�����W�9Jcn`4Ґ����ZlU�QI� ������!�8y���q$?�34�cAS�<��|N�]��Uڼy�y6��.���^���9����xm]m8d!��FUp8e��)��&r>'���WA�6��`txt�Td�Fa� V���L������5��k}������t�,���f)��$E��L�RZN���*��r6���w !UU3�B��#����v�_�PAQ� ��w0�*�"�cJ��. ���pCC�%JGb/4��p�O<���H���<�}d����Pq�pO�����?ǭ�f��g3pq�����6I�a�^u��?�(������ڀ-�ek��6z��yN����7�.���3Vs������7]VZ�8I81v�Cѿ������O����a�0E�٘<�=���6겅�[3<}�F55Y���H�X��i�����uظ|!���Db�e�ں���h4 ֡��
`� (�)p�i�ݽg�A�m�m�`�x��v�������b��.���'L=t�9'�",'$�iJ+��u�l� �r�a9��,Nй|Q姞zj�ŧ,[4��.>9�iy)��| 6
U�F���©T������s�]{�����M��|�,rNCc�������h�]�n���?>�\"�*�p0��3%!|S㺄�3�t�0>��Z���?na!J+7�u�<jaz���u�]M��.��![0��q��1q8���pg:7��l�ω��4L1E����� Gh�v�|5k6^���w?�O����}}Sc�r^&�<�I*��6t
%��%FFs�����`����`���9��`
V��b�.�$R��v�fē)���t��.��cW)NB#!��H�y��j4-��j�	 ��F*8\1"y0�ʃ�ͯ�9~�З!���t��c7l��F3�(��������2Z��?��'ţ�z&i�J��蟐ش��=n��f�9T/�J(S�\�FcNo�(���춰�k��F�� X�e(��;����B>��c��и��T �;�P�����d`��
�~��}>����w���d�'��|��k����[�~�{��BM,��uxC#�q���Vf��>fv�4�
(�]�����f�����P yE�T���|A�ؒ��"i���:F�"�Bx6h��2�l6��xg�0����\�h��F$	L ��{`����s�[�81>�u�[�V�"hl�;#L�0�@П{��%���O|��m�}��g��M�i����9��f�~���k��s:�˦��=�a?y�����-W_$�,ɫZ�"��^b��'Jo�S ��3M\̮h���Q��K��?e6�����fi�$)ʁ�$���2ju�����D�B1�r��k�h�$	������{�Pgg��k���y���5��=1Q�DES�s(q����x�N�n]$i��a�d5�a�O&��c���B�\7�p��i����TCW�$A�����P[k#�k�t<11�OO	�)��w�r�5*ćh1�f�b.��=p��œ��P׆��k�������p����8�G?~x��λ>��P�I�e}��I���z���Z�R}4^��F��cż�(��/=�M�}~���	z��}55U���<�l��5D�M����
�B���)S	�ǡ7��*tE�*S5y�e����d���tֆ㓣�#�}}6�����AA}"��Q�� ��<�pIF���<Q�� ��ఏ���b��6΍������d¦��C�mz���r�
f	[eC���S����<�c�C+�k�ݿ���.����tb����tq4���'Y��I��U�FP�I��4I"
��Jٸ\Ȕ�b ��s�E��s$�l<���t�ĳٚ���+�Üd���l���H�R-#(���va(�m_���D^D�v�����9���ёɭ[޹d���Dr4��¹M�&666�](���/[w���JXM��k�����,�N!3�i�,s�؃ `�
��t:�*.k�Y�3 �l6kQ=�u�m.pq��ٝ0Ɗ(b$%ɪ()�T���c�+�O[�b���
��)&	E��eE�[ZZ����[�?�|�c[�y�/&gط1���"/K��5�[[�������X�@z{N�;��������h�Q��v��{"���[����/1`�b�!n�4�5��?!�{|
��7S2��'��^8�K"1�0e�%9h�1U��E���(i��^�M(d�����N��	���p:��UUr�H$R�ţc��~���L������`��p��O�xbj�sє�� f>���g�=��	��ظd�2�����v�pg���<VYV^8 �\Q��i�������vZsk���D�,*�.�?����BSs�N��575��;�d�h`�op`�q�x۵#�Reu��_xn����}�=gcY��{o~��=o���"�z�V�j �4���_�,�e����өaF-�ي�\���u�q��15�I���ݻ���zf����>1�pr�-�e���VR�.j_{Ʋ��Ӊ�窩�M$����e�M��Һz�Ҷ2-�)\C܄���HdV�.>k��uk�<�T`ɂ�*����;]�������C=������"-hW���.m��s�����=�)����zU6�x�m�Õ�}��u&�'V�=Z��:�]�Hط����L��/�K��/��������}ӳ��(�s��R�d}}=a�Z��X�t���@���h3�7�&�����?
hm7w�t 74E���.Y�`j2�ɤ�b���?*�����W���
΁�c��*d�P1���N�ұ��B.�P�;�v4444��tuϋ�7�G]�1�� �Q�\�K`�hI����< J�t�	(�����^J���갿|��U~C�R������r'�PT�`6�Bw�rR�� ���i)H��X�����H��

��n6ɂ�-��`��)X,���i���#7���9����L=�H'w�.�����r�I���EÊT����q������t���|��w�Z6tm6M���|��e/��³�<�|��;
YLyCW�,��a� n�v{���ge���c���.���T]���
�������50��'eS�:>¿� �?�Gh%f�_�&a& XR��.��c����HuXyӖ�m����uE��B}��e�'&&"e�p8:::�(���X�ܹ����p(�X�Xc����Fc�e10a����9s+*����	�iF3�ST�3UR	�(�R��9洴�|�ei��)E^ЌHM}YM���������L$G��Ag�����4֞{FE:���yj��w�,jz{˖��vG&���g���k��m6���?2��_�Lg�'��7	L��|vXv�z2�pp��Ł?]�������LN���\:�ܱ�]�0��{�
�ȃ��\u������G��rR굗��Զt��v��1��?����^�T��L�H#	�(.�蔻��'�N�!@ ��X;S�Og�|�u;B�Q�����c(��8�A�ciC��!�*�(��b�Q��*�CF�*����!��c���i���t,�	�{��G��sXec	��w�S 7�ܓ(s���´+�$�R��W%<��V:+.(5�4��e���s;榦y��WQ�����J�Y&>9�T����zeU����ө�;;����6֬Y]W[�d�O_Y(�]¡��!�F*
 H�ds�I2u5���-F 8�aV��b�h����C��6��i��`	�������(G�L����1{�"o�L�$JM�����`ʱ�Hi��pR@�$������gs�`H��C꠪%2P8.�$*�bX1E lhS�Tz`��NL3w�1Xu3�;��U4gD�NU���KQd�Oe������Fk+��b;w��b���֖�^zyٲe. ir扔�Eww<��\�v߾��;w��ҋ�/���v��
8e���f�p�#��yH���������Զ/9Mɓ�5M������R� ���3�)����^3�[h������D`��'0��lt��)��d;�ӔZ��<S�zKG���F�n��a�8��裏~�{��m��v�?51	����f{��逃7K`jf�ڿ'������������Mg�]�zv��=000w���\n�j��f�M,D_����w�~��'b���^QYUi��E/�.�����iL��U��:c�?g)N�4֝��F3�Uk�����#��=�908p��Wp����x��_���>6��f�-Sb�=!�����#O�0��Wq+�s��+Sɉ)>959��SM���%1?�;<=]`h���'&'��ϟ��O����U��S%�٧�>�3����s�6T���/?w�S�39��D����+�ܾ�^��9����"H����l��*%]�9zTS�&���5�\u�-�|����m~KC���r{�UU��iE4S���R���Qf]�٬H��,8
�>�R2�B�0�F~��pTSG�XЃU�15�Q
aGʷ:8����9 > ˲�$�`��۵��1��훕��`l�o�˷�S��K/������_�N�U�˅��&�/<�9��_zцֺ���#}�l���=
�vgeuE�8��'�/����(�_�� ��������^7�+ FҔ���}[�uA�{�ww̝g�!���&����E"�B�P)x�<G7�R�E�Bd��ʌ��[�9�7�8��g��*��bHlV�m�n���������PB)]�EB�@��j���.iPh�~�7GC�����no�Te���ég�y���+*+2�i�$�.����y��L*yŕWR	w�'�Yg��������ϫQ���:"�l�H�B�n��
ىl�wx����%M����U����o����^��h��>I!������� >��%2G����q��:a���-u����~+n�ޚ/hgm>�}As��~�-[��憩���~��?�w���?`+�5U��F���-�6I3>����T<��m����K.��N�`��` ���?����5� ��LX��ʜƙJ� ��p�w�����?�i+=>�ؤ�������ι>��+��L&WX�`њի�����=��������H,�t����}�g��8��pљ�VQх��K��@
�_�pq!1�f2I{���EL�1��-z��R���$�����<P�v��W��/����50�� �7}�&�P����H���H&��2C2�����mX�k����.Y~��&U�a�#�������io>r���w���Ӷ��������?�y]�� p��8��@?_����VECy��O� Y,�4E`N��jTeY2U��+`I1b��}������x&9�d/\�n�e!�B��܋ �)�*C��i>'Q�S�_�HZ��a�n	X����r�UW-]�,��?��_�|��A�z�������{���^qڙ�����ο�9���΃�=�����/s��H�������X�XW���t����O]V�&	�c�0i���o�������t9��x|��>��`�N���l{���ƕ+V��d|����@\5�3uS��,���c����~Be�0<n����@��D蠦S#�cG����|��G���Mh�Sǐ <��k� �@Ӵ5V�L��Y�`.j�vbUթ��,��p���Ti{V��z��SW,����$eT��~��ny�-�о��/�3Y��kin�
��(
����zՙy��Y__�w�UY��!}$��d3�^iMض��c�NLN656._��#� �����+����ߵ}�~)�Vk8���e��?A!�O��o>`eͪ�3&�s�r�J�V^lF�ʄ���-y���Z���W�ni�$J�@g@�ְz��r��������K���P	�����9U��9©J���s�Y���6!e�)v���r;].;�ᤙ8j���	���#�ǟ|rpp��h0s�`p۶����uN��=ẅ́�,y���k ��y�qM�����@�Xj��Ϣ^�6�4�|E��{׋y��"�%�{b����ٗk,��F%�����e���J1���^���rW-���[��!��;m�O]�n}��/W;w�c�l�o�|��n���=��:��śnطwwu���8�6�?Ƌ"U(r���B:!Rj6��j>o^��M�"��Ɔ�'YC⇇V��.)�(ж�(~�+���ܿ�=@���9���9��Uۿ��9ms�[������=���SN�y������P,�y^�����9K?��3��v�ޣ�������o���뗬@��j���10D���qCH���b?�*L)3e���1Ӷ^7g�Y�Bh�>:�X��T���t�_����n���|hph(u��؅��t����ʏ�Uz�#cx|�M&�8�K�wN�Ѻ*��E������$�ͦ,�H�J��X��h���u��^���+�^��?q�ͷ����6lعs�3/�x��Wm������w�vK%F��C7��@f�����SK:�gK[��jd2���z�kn����;�u:\.p��/�S�t �L�7E���<�����5O���0[A��t�
�>�)0vWe}]Q#����~������GP��m��?���I���QK6����Q�0�&����eE
3E�p徯�O�eUu8�.��U�I���k�+��vݥ뮼h�A�(�L��(?!����қu���c�&]֬m�7 >Aa�O���9H���P�����u�����K�b�%*f���$\2B'�*��f�3O?[(��x���x��J�adQB�n愦X)�#UO�朴�^��j�06��S����76���1�}^���Y�n� [\Т�7�p�왜�XsιM'�ɪ�ʊ��"9���PcT��fI㟤�b���f2^)73���j�!��j7���ض����i�U>���%�z����S߼��aYկ���]�P�`��d� ��r����\YC��~�X���F�����D�^8�a���.�����l�2_�+��P�^�K=�Me8ԹIʐ��	�� �T@~6U�	�E���+�Lǧ�T��/\��g^X���;�>�����o�r���.����g������.����G�\|-I�9��)+k��ݺw/�'�9��ғ��`u�7V�� ^3��0�	�L������H�\)���],b���1�a�O��N�l�s��}�� �"$I��L;\ɂ��KY>��L�85O%�unlRL��na��8��-d�^�)]<��Þ�1B
	^K�'w��v��������"ER_���3)��_Q]���+�HG28*���|b�̨�!9���1�`��+f��=Ţ�J�㓜h!H���y��^Z'(�g�IE��Ȉ��ڐR4j3��4�g�lNd@6��9�@uK��7�"�#@�X;G�ajH�P
o��K��60@Pp^�=9�z�'J���4ʸ��+�/Z�X�l,�2�p�0G4��e$?��t��fZ5]�.�n�(R���tKJ3�9(j�vw�O��)�U��vy�f�P�p��>��e&%y�;����+�H��c���(�0�����;P+D�VdQT����C�D���Kq.'T���}�-Wi:+H���EbDQ�N���:\�,���[j���c	q��s�E����`��¬�N&T��XΌ��Ј(����	�<V����-|�R'/r�H=��3�w��~|��܋"̞y`�~�ǚ����w�<���rӳ�U��Z��~���a��������w���+7=�xM�����-7��?�w�Tr����pg'��^~���1�b���H5�6������)k��w��0kK@�m@�EN�D��hh'|aG�ࠋ��c6^qv�f��[ߕfъ儦�ݷg�v ��ʪ�c��ƫRYe���X�w�R��4�ٱ�]y�5?��C�h䧿�9#�g.^Z!{��v����d*K�4p�P��>ه��B��@�����_P54������+N;}t8��#�^�aö�޹��;kۚ��x��CǎĢaY�r��SD�����Te�̙��W�����g)�Xee� �"o��c�(&�N�`ZR6����)��֖�X4��X}M`` �=J�������-�?�H��=��UE�ZC��v±�D�H���}�P0���������X�s�y�ٽS7$��a���*,:��Kl-S8=E#?sy�@r���70 $��R�f��+X��ֱp)�j��XW��b���fH��2�,�/D_	ςa�x"++�����d��WG�zIü�N($J�h�`�d(p �h��j:��$�K�'�0�����Q:>¿� ȿ�Y�E����&�)��	����&���fm8�	��<�l|RNLN�j�h ��
&��gr��a�����Y^Q{zz��i ����t>�F�Y��&AY�2`�s�"�p9=L>�We�/�/�T�h���$O ى{�sM�J�9yZ�in��7jQ�{Y���$��u�o;����
�D�gi���w�75����d<�˟���������Ɔ��7�>6��'?�陫V����-����/h<�p��#%�C��o���?��g(�qhd�p���$���@T�^p�2�#;ڲԁ�*D>`wy���o���ǟ�E�����-nkkDq|r�����Ҷ���"b٬+�\uO�1!�b�����׵� 5@ʿ6����{��#}ِףHri�TH݌�d�cH�Ic}�1.Ө��EdCI4���F]��|�7^��xކs�j�������*���\;���?�	�;n����+�i����������\>�d��K�-�sT�ytttdd/@�fg���K���V�7�"������$о��Q pN����^���[��ǐ�H I����Z�l����P,��ʛG���}�/ȚF�Z������s2���&'�Z tR��1� �!�D8�#�X �����Rp��I��9���~�ƶt�_�t١#�y!�$	1���5�;��Q�^��	�O8i
"���i�c9s�@L`Y�`��LWM��������E�1�e܉�Y2C�3��J�IC��M�����]D���!���*I�A�;�I�����F�S�q��,�5�&���1%�a�d(C�����L�jN��y>~s�$�?|>#-�I
案
E���ɔ��U4��u�&����L%_NP��1���WVߢ��~����M۞	Y}\�pvL��.�D�aV�<���+V��կV�����w�
V�Zec�5kN��?����ؑ�_�羯���6^Y�����On�zx����|���׏��j�^���s7�t�����dmO�����|<�֎7�\�vt`�� h�[+�k��Z7Bj�(���\��g����ݜ��}��U���߻��G{��憯�����;�]�n�S���d���m�d����'�|�����䳹l����س���)�({��O�W/ji}i�K�w�I3�"�h�zb�p���k�f$������s��_O&Bc������sK�(|����<T�������
�#?{غ
0²
�[E����)Ī��p�ծ�SSɷ��	�v����q�ށ@`����4��i]z�ރ���:��[j���ɻ����x�/d'���>���TE�����	]6ͺ�&���Z���X�������w.:��M/��4����g^`����w�;��4T�dIRX'�r�d��J� b�2�4	�R4�@���8�"��׷�?������SmueQ��07�I����N��־;[�OU`Ez��Y��-+A�=�1�Aqw	��Ob3�س+���?I
��e�z-t~M�)�کjC~R�G?�����q��h}���c\n'��&��勅�_}��w�۝n��𣢨HKWSE�8�����1�""�����G^��}�|�?���k�c��J`/�C)�zCkc�
<�9Z�e�F�G���p��9>�3eҌR�ٽ;tkƇ;_��&��C��6k��.�5ϵ�ј7��^�*�î���T"�v�y�me�x��2���&�ګ�,����
��[o�i����^{���õ!��b��~�w����];�n'�Ɂ��w�j�`���PzxX���M��5�n�l�yGG��N_���{���}����.=_Qq��-)ʱ�n�b�����;���VU;z�hEY@����.���+��s^�8ċϿp�m�;8졇?ph/���_r�����W�>o�������)�F�Ӕ��M�Y�'�������0Bu=(E
O8#f�����m�͘T+4k�ߡ���ZR��{���go�I3�
B�YPY�]d�,M���\xκ��NwJ��9n���nWG�|U�lg�����K�'�~_(d�Y��q��+��y�"V.������P1+�-.��5IDIK�lb����y\˖-����Lda�u�WF�Ǌ���+�#��ٷ��v0J$SU��d�A��_��b`yP�$��Rd�eX�f�pHYF(H�\[[I�b�A5�V���.�}��[qk�V�$�TH��<���C.�%��X�lGB�����̦k��/��LR��E�(�j&�>1�O
~
���c&�D�R�7SI��5)>��	:RU~vE��SV&�SM-5�7]�ǫ�b�_�����p�=��p _H�NSMQ�]|�P@����&IT,I`�6��f')dT�Q�2�b�C�1S�C�ٶ��p�q�N��B+��[��V��GO5��;4��C;x����tBԴ���&l~aSc}m$l���wnnn	�n�U��^c��|����sV/O������E]����v�.�^�N'��������v7�B\17>24::��ew�v�g�k�����J�j+�h�|ă���.��-��]��med�3]�+$qdj�����1
,utd(��c�u鲪������כ[Z���e�}��\z�7^�����y`�����[�]w�-7���K/�\N���f�(�d��Y�Ŋ�����b1�t�l�_T�h���ғ��-���j�z�2��M�TqK��[S���������|������H��t�s,
��=�	�!i�W^��/�ك?eB���D�sY$8�J/�h�t��(�����Æ�*��%"D�����-���)��fY�����Ɗ�:���4�<,��"ኡ��p���p$eX��r�MS��9�N�������'2 b4V�cT&��	��S�TA���i�X�-sь.R�6������$_nn��g����D�ɓ��r¯�gr�ͦK�."����,nc&7��?1
(Ԉ��G�H�-e�Xb����@�W'���L�OK�h6�#IS�����G>�S6����5�sE�/����#��xgZ�,�����ygW�H�[�?\Umk����l�mx����~_u������>t��`��y��56֎�Ooz�ѱ	p���9�̀ T7�5�cK���� -�Nc������&]�I3�D#XS��T����'e��8��b<I��:z��!M<vۏ���=������}�,� 
�M��+�����揿��/�>��3@�];���/���������_����o����:gM������>����Қ�������O���%K�m��7�16`�/�4B$�l�}�l�~ِ�l�� �z7������e[�z��M/�����ތƅ�$��o��?!My�{�9�S���ǖ�����؈�w���7��2a4z��f�!⏕V�45����Hycǜ5kE���?��+7\��+_���g�O�ϭ�޳ۿdI�w�~�/�᭖5k�H/-e�ip���&N��K7���R+�ȶ��!E��e8-��q���:j����y����3�{��"SE!�jN�$��T�P'`�NTF���^�"��H��mw:�gw=�Ǉ*K��"p<|1�n~sks[���yNO��h���(�$HBs�J������
�Έ�l�"���9� �}(
�8h-£d9�ÛL��,py,�}�ߧ�I������C�-X�jy���8x�ݿ��Ο YoX!$S��ڴ��` ��ٹr�����?���p9J8D�����k�z��n��2k}�'��DP��3
j����B�F��_Ճ�Z	��͵'��Ƹ޳Sw��V >��|z���p�=�:�s��Q�������Q\�I��o&n���
��N[�
T�2a0=1������ �����T�\��?�����ZW�qْ�pSc����=f��k�b���޾��:`7�-f;��+�ǧ�ť���X:}���G6���=�{�y��K�����SO=��뮠p���S�`��ME�meN[�"H#����L%�Ĕ��VF���2H���V0
Ri�'Bsܝ��C��*Z@�(w���.;��+7���;�;�#��*ٿg�T0����[�m��w����ǎ�5�'�S�d<��e}����3��$R�^[_(�������rg�W�r�pAc\{���ߌ��8]R&�H$2l���XA��"*Ӟ$��A��T�lk2;0���GX̩�4�,N�󂵫�f7�-��jC]��̓_hml��)M%����7\w�0��`xd0n������#CC.[?my�����H����nÚ5E59�㾓��~�:<c�)D�5�Ӛ�U�j/i�fɼ'S+��M�ɓ(�d-Uf1�$p�]�E0I*r��v6D'}69.�Se��b��S�O�gy=�щ��O�e,������*P����i6j==�9�eqƻ�֒F~�;��Y��G{F���7���`�N׶m�����ڋ/���oh������\�St��t��^�����rی����n�~���؜��7��nh�A��6���p:��x�H�Ί
e�ˊ(��-�k�TO6���i1o\�~=�7���m���qr%:T5����7��K'u���ݓ��it��=C��?WGxn���8���BN��<�r���1F3|y��e�/� �f	�~��gz��m�!Hʅ+W��W��t$H���K� ��/*�'E�����Ո�F�
�����|`��{Z:�W�^S^�*."�귬)f�w5���j	<��.cCZ��q�wd���H,0zӥ��k<P�r�)�~P�	�:T��¥B ���
O��0?��*D�
DR����ꞁ1�0��7^�J��?�p~��n�=vd��Wl\��cO������W^�t�e��S�����C�W�Zf6Y����w�8�N�ENHF"�񉖶F�!���@���� AF`%I�b'h�j!q)p��4O�t�lL��C�cq�xe��O���w��.�xcG�ܵ�V=��Ӊh�������O7|F�\S����r�W&�d<��}����c-�-p1ly���_���뮾�O>X_U�����KXj��C�jR� �$i�Lr�lͭ��C�V���&�.\BE�:y�Zf�i�.���F?�L�8c�:7����x4*�e1"'�0-���h��r|�X��Bמ�=j��
Sc�
�R.E���Ѓ= ��g���-x챇��*//�3wv(��M��a��p�o�[0w��K����>119����V��zK�����͟�\_�p�<��!!W�h)^��'����8�{�Y9w�������3�d�39T�8N[�{m�ɨP����� �Eirk\�a @)�ɦ�6[2�.��my�R���}��X�Ԋe"��ܽx��!���Ͽʥ�}��,�C�8!�5�ش��T��ჟ����
�kC#R{{��D���u�iL�'�V��H�1�	"�ӗ���de�B�<.���o�}z���b!�)��|.�<YJ�C��l H.����o���.���ڛ�:Uѱ�G!V^�n��6\|ϯ��d8�����n�epp��'��GS�،�&8K�x
J*�:A���
�R�A�����B�$�]�rb��#���ځ Ge9�xѬ�/Dj$0e^ ^�z���s�p`� /Y�3�<	��E�u��.;~��絶�����L�����ل�_�}�m�v�)����c��>{TF#U���xIH��fTX������3U4�~�~8���*�^ꮧa�b�8=q�Z�I�1Q�B`"�hW�H�E��i{��@�k6M��7I��f�1��$�t*C�4\��kǑ30�Җ���rw��s�O����i�ٵ:-�I*���?o����-�߼���]s�U�M�G{{"�`:o��Z�����ኊ���=��=~������_���X<<��O����;������ؚ��AH��F�k	(k*Mw�膅���P��'O��₅#�1�܃�V}�^��������?!��s��CD��� (No����G�Z���U�e5�+�p��%��(B���Gi)�1�T$H�DK�L�g'}��dpVG���ä���T�$Y'x�U�$pe%ő��/��'?u0��~��F2g��X7'����g �Ԧ�4&��X�)�/0����utp�*������� ڵ=��������r���,�����^�;8x��?��y665<~���`�M7}	���o�ybb�d�����BlsK��7�T\l�9��P]��O�
ˊ��fh����&��TL�b8�?l0�6��dhD#"�2>c��1�m6[}}}&�	�B�͞={��~�=��zxt��P�(�I��j�H?49y��P�d8�D����omn
�uuu���F3n3O��=��e{|-M-V���fRQ�j5�j�(Z�Ɠ�W�̝1ԫ(9�Q�+h��W_ޢ�럑Oq���tU�,�iT��9_��F�-b��c��_��� ���E��X8uڬ�M�ć��&@�J[sXAq�^l���j��>D�^eX��J���2��v�yN���+V0F����?�iSK��_����3g�Kr�������v�ڻw��W]WVZ��K�n��,f�񪫯�5�3��DB�M�/�!S�P!��)r�{���!���ƹ��7^A��	�}'�s��C��C+��{6*���`0H�l����l�	_iI��i�t���4:[[)��j�%3*ɡ>���O2�pх�-r9AϾ�/<�x��� ɢ(��hpڱ����n��y�5V��G?���L<��߰Y(�\s�E:BխH5a���`ˮ}��'��"p𘑃��^���d[]tv��S��G�`��L��i�do�)�=�&�;Hs�+��K����-_�
�b���E��~�����XGk˲�T���%���x��L&UQYj6���f�ёI�T��p~c`�Mǳ�bk2ƒ��M%&�㵕R]q��R{�/�wc��`��<c�\NWY��ᲈ|:ͦ2|�΃��o���P�޽GSI��H4&�@屌��Gw/i�>�w�o�+���c�3�?���TIII(ص�����{����ee�]~���N%����ͯ����٭�"�����5Q &�t�P��$�$�p��Li#��P����3��GK���;��S�H
Ț�a�o�Rs%��e�+�q:��#,q�h_�D起���U�o_��,GC�Ȅ�a988��P�zu��P�"�
ʥ�T�^x)2���"g���B��+�]�iUS'�=�y�&Xj��@��ǎ����/�z�;�lk卑9���J������-_����� ��X:72�P���v�7g��c��i�p�]�hl�{�Q4�+S���}{��)��YRZ�$QU1�5Ө0��[}\��z.-A �'��6�/��c�'���P�is'2@�9E���j���a�٥%5�� ��N��[L�m-��	Yv
��dKS#Tc'���^q����8)K�?.!�e�.�00 ���(0���y����BH���#�xb��EP��VWny�5xk݋;���ё��aD��hBN��<���{*�F�P�:0HًY� .��!`��ك'F��U6%ӡ`
����-C�;�;:�*s)�gϰ�f�b�$���|,����OUUTP4��1��FC)��H4��P����X$�u�X�[o�&F�[���잝J��?6۳so�=�X(�LF#"��A�!.,�z-{s{�d8���ݳ�ϙ�&����vK������'��D(uy���Œ�4�����-[6���+5�����oBIZ�-��	����zxx���ꪪ�2����C�^��B����F9��HU>�����oA�jg^��`�`h)@]o�=�5'P� ���gL�Y��B�z M;�� p�����[Y� W�����ʆ�,άk��=z�go��}wƶ��Y�C��&\V[���X.C�,��4�:k�z>�ؑd�O��]������}��{Ƨ?�1���mW]�q||���� Q���튂P[W��[��}��7��VS]�l�"����������,� ��XS[W�;�vTVV6��UU�4��jT��I�M"kY�`�����gv��|��9ExVC.(T����	�o��#�͗ �J� !\�G'}�w��{��i��������[i9��/=�';��l2�H|�?~Lcد����m�[��-rCs;�'�������t�O���׿�����7�_}�W^�ѠH/���=��kp��t��fTʊ�o�LZ+3��@��K��'H2�:>��XTnw��@��rĳ����yS�������_�x��D_S�_s�6�(�>�>�#�Ds���/}��-e֞�x6#J�l�����������YՉx�����(�G�
�X���.�o���	_�f,��n3�3ft�Ӊh,�I���t����m6U��?3�T��vo��JhHly}k2�u����
���Ǟ|~ђ���ޫ�\Ǡ�!���R��d#�)�
�Hէ�P$߸HSt{{�k�J1b�L��FQ��14�W�h���s2�p��+�`������i���w�0����k/��M��,ͤ5.~յ���6�\������s��ևLGS\"�۬F��Q�j��N&��VA&�~Ɠ6ݙ+������[A�����1�N���r����.Z�=1Q�v�����s����톐r���5�5�$g0�K&���|��`��OF��wح-Mu��j1��$�)��3��sy��`Veh8�΍�u�S�z�H;�}��T����kY�p�Q����X����Acb5o����qP(��e�]��R6����� v�����`�/"iS&������2�ɘ�G~q��2�M��^H����<���4�QG��ϝ3[�&Kݶ#{�W)J5����nOFt�j戄�N����WU�Q1D�	H���	��N���Hbʈ�G��K�uk��[��о=N������p�=:�PW�����'��&���5�o%iö��-�,���c���������a4ێ�(}�ͷ�j��X���>��s��6���7��k_�h�_�e/[�+>V��BV���*4�xE�(�2��D]S{4*M�7ܰ�d������w/�h%<��˞z��_{k��e���m�{�W�]K� � DJ��!Q��=��l
V�@�@�  j-�h"Q�L������W{e@��x�W���T��oVH��d��§8��j�VIl�l������>���.M���w�.4�oni��Un?E�2�\b�*>�id����"��MFOG=.��&+ˋy�+-.�� E`�T2���T}}ct*DTYyi0�y��tH����Lŋ��4Me�lUu��,��������p;aj������u鹁�9E�7�p6E����\JB��¡�����_�e�$��T����x��)<���Dl�N����̒j���T�KJ��A÷p�QE���D`�-M�^9��$������&!�")UT�IH�*j:�Lr��� x���%K>��6�@YݮꈤȨ�6.�8����H_�˲xf��$�
Gb�nP�����W��7��"�낕�05�%ۘh$��"\��%A�		A%ّ�QIL��o~¼�P2��(��s����#��>�:� �.\���%�W���{�7TV�l!��"�2<gޜ�I�SO�j��W�Z�N��~��/}��u�<����`���\�A+��?�����Ī������E� �;����� JT�@�Jˋx	�Y.�f��T}{������Ñ������Z�L�}�P��pz�%�?::
qG����TC�� �W(y��ER.�� x�+z���i�%�m/|]σR���T�4�����G�)��:��Tz���twϵ;=?��>�������;�������y�����%6\T�Z�[!����I
3h4\�&�(��]uE�O��jV�L5��^�!�D>+�l��?<D�$)�������|*�S0IB�d2b���%bA��hʀ�Oʔ��Y�@e0Ф�����m�ڳ]1�RUՌM)@׍k"A�F��TI^T�3���/G����q=�>=�\��
7��M8��v�~�$�s��C<׷|�QB=�-Ow�t�%���iy�, EU�J��rIު��9*5�1�Z(@��V�71����|ŠU���"2a!Z�ހ���Y�H��h(D:�YQd�|.��	T{Y�8M��VT	MVEgɿA�2Oȿ�J;P5!��jN|#�/�]e����e�	%+�B `���"��KrF�^S[YA;�#�/�~�׫�˦R��,y���<����E����̄o��������������#���#N�W-�B��3���z{[$7k׭� !�o��MW�\�����/Z��3O�&��=�:RH�X,ͱi�&�'���/�
Ĕ�mk���biI�|;�"]sf�ܹ��DSs�έۋK��y�ko��G��y�Z��ʿbB�T��Rs'��ʿi��H��t�:|dۖ��MM�?�xCC�?|⩧7l��s`����������o����9]]��P�P��d��&���<�|Ԏ%����¨<֊ZP����MT=�(�H�����3�������k&ԺI5� �(�qZ��L�7�Ү僣*���$����9ExVC*p�h�a���x��ױ�����+���_M<�(j�ot�Y3�Ժc�5[Q�NL�8��ҟ�8RMR��
�3ek)�
��_�J��,f����CZ-	�A5̯2p������,��1���u�X�Q1W/��v��
 (����T�cYM���MT-���m'y�1a�(Ƭ�a�5	���F¾��֎Y%_���o��J�����K����E��@1#ms���ޞHf��\OfGǂ���dZ-
���J�eE����x����w˼.1->���f4���j��	���Ħ��#�f��( 0'�P_]L3 HN�"!Y�İ��H�MVk4O$R7��e�U"�������z��U�u���ƓG�������=g& ��� j�(+/��n�1FX�;]=�pI�~Q�3-����u���ڱ�7_]:����40�o��ӗ]T_������ٲ~���$�t�*G*g��g���N�Wp��ti�zEûz"%�TPVSP���g��Nh��(P�I>rkcZ EK�QO���^�����p3����w�x�'*DyN~��Z��3"Z�0ځ�Nk�i�aZ���A���D�i�2�U�	��O'�)@��d\��)��TCY�m��rGy��pS����CY�nA�f�z!HR��ȍ*¯�<|�#a���pCu��
"P{��Y���7gh�p^�)cE�����I5�TL�z���P�j��"�{a{JQ���JYv��;�k���\2k���l6�HG�z[�K��Q�H�ʕ��=24:���K�{�u�7o}睝"�I�f3	Bጴ\ⲔW�n��3����T�����=������ݠ�/�w���,DC�֖�K.^�pZ~u�ccc+V������8�{����n���+.-���f�Z�fͬY�����X<�^������+�k�|��nܰT���6��� Z&Kp�h���Ar�m9�)œ��I Fb.�FD�ͪ~53����~�,��w1:6AB,�Z���ŌP�Ӡ�����3H<<��h$�r��L=�Yw�8m�^n��EmȄE-�4�����J����`��n���P�/�7�	2�_P���BMd���V��T�%��7˵��p��i|�	�;��{�$�+���P7��s��th�z
v���_��)�W���"�s�p�S�##�H	��W���I��t�A�}C��J{e�dT�4�Md�_=�b�r��B�Jj\���dysy�}��=��ͥ�m�*�L	\� ���yJ�¾z@S�y��j�㒒K��$M�%f�	��!,ϳ"H���B�FK����g�?��%���V�PZ�H*��y㺹ŦtU1cf�%1���&��.32�`���G��h�������+{��9�����>\"��,���o�[K#�ե���N�CR˴R�,�w��%hj�sO�����{���w�d*���m����~P;c�����w���s�[
Lv8hI!~��������#*/���+�mz�կ}�[)��r����C��_����Ә�0,��TP�V�ab�(���B<�����E���#I��8�y�I���K��,�&��A��)
5�Mƣ6�-����P(�����i�P���Z�h6X��%*�15e!0%q�c�)���Pj�L�Z��\U��j󺰀����/H%re��T����b�j/u�"E�U�A5;-M5IS9��9����/ r�6�����t冚�� !���	�A��@��f�Ȧ$U��*Q{(�".@��I&w�YS�k!O7�p�)#ߧ�����(>w�|1��������?S�B΋�S�����[��DA<W��ٛ�
�N61��Fw@ɹd�b'��(a��1�|����R��%Q�1��7��$H,GI���,Q����H���V�qY���$D��a��ZS�x˵�U/5�ɰlR��c�=n'|OP�Q�X��!�1�q�=i1E!�#"�X����(!%�1;�t�w�	��ȥ%2�@�bA	�+%y^�S>Q��_ti{{�_���bZq����U�4�(C� �^�n����M.0�Od'��C�����P̟�Λ�������ܻ'H
����ʛ;�9���5��#�HT1���E��|��ֶ��~����^v���d����_<>��
|6�U'J,�7}�Ⱥ1Q]Q~�o����2(Ei�t��ɲ��fI"IM�|1�(��;Be�Mg ���	u��d��'�nW08���3���E���!Ј�|��B�� ˤ �#�ޕ��B��. �@H3�rN7�d��R���g�x:�%LUhJ������<�B�	�:�vO�|�
�6%���:QP�ڮ
���&�l1�P��Zu�
��B���$Lk����s��g��1�ِ�K:m0P�T��h@}�S���C�o�٫� ?mw��H��o�nQ�4����324���*����"$�9�3I�3+XQN�YD��"�"�²	�ԚM�6j���"+���d�Y#-�#AxaPh"{�w��~.�&ߡ('��k�R&�h������2���ˋJ�C�12v��*�.�q�v�9�q(��b��b��r6"���v*2��Q_�fn���Xm'Is��d�qY�Ȇ
�9sFkS�����/X� ��rl�&���]6�!����B�T��?-�W�L�;��l��#d�о��o�9W]�d&��=�K/o�x��y�����kN��O?w�UW�[���++��1�����d�/�(���Ј�]���K <�X��o���'���(5���y����[��~�ŋ��86O@��d�>�
�0�IB�766�{�n��a��(�r����m���^o1Tp��h4A
�tw4�GS�P���|�2c�eC��¼�B"o��J�:I�yY�M���F4'|�KjR�FU��O[�/���T�+�k�4������q�0���Y�j�5��L0��	=�So#�Q����նV@��Q�����R��w����3�)8���!�s���?я�ύ|�=?��a�3��7���q�v���#�d���U�P�]�BOݹ�@O�U��p3l�~�f��('s�� �4��"�.�D���K�V�[��E U�Pi#P�&3�D� ����ϋW��q�_P��CD(�yN�Xl�9����%Q��b�߱�m��w��7�&�i�"f�pC���'������9K�hHh 8Ӝ9A��r`rO�	��>�H���V���]�Md�
!O ��h8Q��|�_���O�ӍW�l�a1�lo�8�2�Xm���e�<�4��0B�^���\�!x�AE���߾�᧏nz��C{8�����V�Xq�%�`�.�n6�$��--F7ݱ�՝�5�:��H��U�|�ͭo}��7p,0���eY�2��S sOW��Nz�F��L&�N&SP�^v�%�Xbx��s������5k***A����Լy��m���P��<���,��Q]طw��W^y�M7�TY^����p��#Pwv��As��y&I��G�V��(�S{��Ow5�d�Jh�"#�� o�D��Vt�0-�K�!r��xp���(����t5���Edp�.++��vu9�#�/�n����iD���C����D}�KK��Ȯ��4�)³'������NV�ZZT�vy(���B���%Vڦ�H��-�	��c�AE���X��p,a���.��;~38�)cyD,��>��QR�����լ_��z�P\Dc��pN�MH�w�a��&�(D�F#Q���Y�a�ˁB�x������5S���g�m���P/C��u3,fs<�ۖ�۷�߾�N4�e���~��?��{{@ﰈY�y$	�����*2� J���N��z'�L�oZ@� ���{�~�]G{����O]�G}m�Ō�C��x<��w�����Iߘ�j�fPfWU���F�d��p�ÑY�f:|#h.���:�X���Ec�q����n�����-�C_���s���B}��ܶc����W._1/v�mh�ćG�}��쥫���#_z�CI�� ��d:8M�CS������ᑱ,'�S���F#¡�[�N�#���	'��~羻�����x|����� �H|�{����_��")4�Z*�v���	Q���lz�9��;����{^{�5�����~]SS��c�UUU͝3jA��w���9�.��Ç�nwiY��[O%!d4M6��h4O��'z{��\����,M5�F�����9N��UK�T�5�SN䓖��O{LX���]�u���Ӄ7.�������l�V�@�>�p<�� �DM���v�|6���5��#/y�X�,=�&
~�
E�_��]Q�ݟ��9l%I&	R�W��yO���qN�5���G��h�K����K��x"&�Ё}pD�d�cx}}}WWMI��:��T$�i|�˚O+���4+��FI#d�m�-r�W_Z]�@�b 8��x:�2rǪ�4*R���v?N���4"��8�s� ����nE��6��겪��*Emv?ϧ3,�E>4��t��0:4b��i����b�g��'���dR�M��-[��zqj�p�Y�dk���
X��$NjMoT�T�/9˞�=�\;���*�\���)��o�?�;�?x���//q��������wfR)#��`�X�D�4����
�|-MZ�>������p���.++f�������KdLV_d��X��/�rC
�1�������]�x�Pr��mad&0pdF��vV��"��d���D�8��mF�7I8N�F��5-�q���SS�x281�)D��P  ��IDAT!	ޒb��	Y�q���،���={�����J���p���+?��{��a��X4&+��T�AQdI����P�8���_�8���O�]�v��7��k �,++��7���O�]&I��r�*�t�\�[���l&����ǡN�������V��:�4��d�$	1�	)Q�����.�*��SJ����S��� ��>��U�	�X�Wuw���5sAM�ƴ�E�ݮ�C��4�Y�����p�8�������s���@=��x4
������-[y�!h��8f6��)e�����ɧg��Z�fMum}4)*)� ��KU�V�)�R�Hp	�+q�箼�Rj��=��Fh��P2�����d�*5P-`Tȧ��B�2
�h�O-�u:�O3I����A�1���\6c2Ѝ�U�'�g�a�K�R�M�?�5z����"�	�-�u�n�p��r�]Ɣ4��V7�sMU��ULw�ͱqH�MF��H8�/�Ii�TǸ��Z��,�������-˖-;��E/����t"��n����؈?�_wɆb�'��45귫��M�������p�7��-��,֣GN8\�d2�$��8x�_Ǔ)��<������o��k�e��S&#d����z��`���wN�f����(Aӧ�t�*�5Y��@(I(|GcM������G��N$�|eU�̙�^w�֭[���;=�m��p�	Mr�4�T_w�]w7���q��q,����E�	-7=�y:Vg�[��n�kh���r;l��!v˖7��=}�7�F��,�mina��x��b¢$�/���`Jp\�� ����q?Ȱ)h�Q8A�F����d��L+[�;O�g�5��e%0W@��L�\#��Bɭj,�/	QL`�u���
X9�U�*�Su��֣��2�U[;՝�qN~,Ck�t���-�!Z���Br��8��b|P�>:Jo@��,��_��~��������Z���X̖���]�v=�{��n�xŕ+V���(�A$
�T� 7@ȿ\�oVD����������oq��us��8���)��yDφ�%�e�H'�"�d��*=���O��0q�v��?�����V��2����u�u���"�6���"�=v����i��'yl����&���>����㶅�pK�΅�Z�Wյv�d,O	��Z��Y�H�� @���
!1�)��3`�{����.ť];���5&#�������/�hdtX�XwiI"6Q E��Hi�b�&c�@`r�7=��>;8�ωlMe����c��g��{�m���(1��R�:�VW�Z/�������$W�e@6����+sy�,-��f���X,z��g�zds�2D��X�@*ѩp,<iko�[�l<<�&(���#6PRC�67Q��f�8�4�jd|�fu���VV��TU����r)�DiTg���	ȊA�a���886���t��q�xH*++w�������eu]ݻ��ݼe��%KәL:��H���<EI9��W_�U��p����<%5��N�I�"d��f�7���\Л	i�\Q��W��KJT���L��d�9]��/�b�h�s]�U�(���=Y�=�O�o��e�~r�9E�яixQ04g�#j昮$���Q��S�f�j�-���(����z���oz\Ο�������g��f�%%��]����c���_}�P(tÍ�,��4M8
Q`j�򔨁�f�$%�ɗ���GF��7o��(���h���Z�'�:ҡ��>����4�<��ȫ�߂g�p���Z)�H�,�6�B)%zv���C����j�����u�%����w�=k&�e�fm6��GF�kj�,�&�@���>��^���Tv*�]Y[Mp4(�4
u�C��z.�֖H�U�#� !��H\�(����y��h4�����E���}�3�$i#/����������%DA��7NQ���Ԅ ��f�F#Y�K�R�x|�7�b�J	�m-u/��tueu">��L��3ZYQ�n��}���8�|޲xh���fT���8.e=.E�.��%�&�1���6'Z�p"�f��l�?�5�²��2�&S��cG���JJeQ�,�q�^qm`���G:���Lf�!Օ�6��L>;	ՁS8�՞�t����T�uFQU@-������!����� �-XD���I$�P�3
�h0�����666��xb�j�`�����V��T�6�'x���.I��W-]���80�/3�>��p��b�`��w��\�`@W"H��557ih �WF٪j#jLO�TCz�!*�WW���-���6��r�*teݩ����r�]!��a*9ZF\k�t�2�O�D(���T�Mej]_�`���G��;�/�������zN�5C���*:��	M���X ��c3P��r���pI@Ѵ T]������_B���~�=(9�ˇ�Ob���ϟ�=o�/����oذ���x,�w�����/myo�/%$�٭�FƔ�,���2˼��'�h��F�W�pCd)��3I��"1��##��_��C(���2���ج%�82�U�Z����%c��ǣ�ȐB+m4�����YN2Kx�WH�-������YcL	i@������Ww�r& �@H9��"��?T�j�T�W�bG/�P��c6@��)^xa@�r;�[Z>w�U$I%���ծwv{ܞ�Y]۶n�f��A��D2��LOj�a������\y~&�>�w�l60B�3��j�/r|������I�y��
Q�p.���B���}2�q8\
R~��n�W�*	h��`�@�����nLN�,���@Kk�-���N�����dWIEEyc��c�=1w�<WU�w��Gon�<6:F���D.@��̄\_�3-�������t:���|k�~��@m��OB���)d����7e0���+PA�`I+<�ǢS��a����ÃA" 8�@	���g�qв�@�����ٸ~�7��~��}����MN���q�����4���j��9Ee�<�b�!3Q�K�ѫe�i	*���Fp��)�IE��H��z� ��s����Y��-�AD�g���L$I����� �A��KJ�L:��=��_|b��o�*�T*q�k9~���X2�t���-[�ߏ<:��C	�MepYP?�2�Q��	�bj�{G�	Úkj�p��V)m% �K�G4%�e���,"�S�@�����E�D����6���PTi=-����]���-m Q�Z��������OM����L2h$��������DMC�]"e�I�KZ����&�b�z��y�-]}�{�}��`R,���9!����s�@S_��臢:�H�?â�ҽ��,j���f6@p
?�F�G��EE�V���0/�^���h��b�t*�L���%Z��JKK_��ӵ��ȍ�5���d`���p�F�ފ�7��P�4{iC�ᣲL�� �i� � ���/�@� �p,���GA$���D�7����#G�\������R��� ʬ�Ȅaë́})<��z��;:;ο��D��x������������@Y{��+�h��NTX�z��E�?��	A!c2>�G�f����KB���on�Z-����C�p+@|����q���
M��q8�p��986��@��I��C�x�$�.��{��l���gϷ���'�t���᳽�#Ͻ�⊵�=�c�����������8�F>���ZKraƊ���"�E���Ӌ1���� z�B/��SQ��Y�\-g�8��>�qN���f|�̚8I�p}r2��X��G��o�#Գ����)\߈��P�Fhp��������/^�~��-�\}�(I���H5��8%��&B,nt�L����,��P@|q�����������9��h4l����WP独�qz8�m�sTj<��,D�V���vw7T� %�(�r��.��h�L�FF����q�ni�AҦX�-�		p��q``$�D��'���IIJc��P
���"d��O,�) e��1)��>����/�a˽	�7|���F ௨��������Y����&�����@�{O���:�V�NKYi��n++��9q���c�Fє�����Ѿ��֖���gQ�m,+dQ)X.���I@E�;�]��Kx6���8�v�޿���Ny<���㧳f�6���4u��(Ը�`(����>:8x��*)��a+�MH@f���8��@�ՙ(v5��aڃ�%��;<
���.��Q��;�c����>�d`Z`�-�}��M��U�І����h��$	&��]&��f6Rf#�۬c!&�sfΐE`�����@k�`�����H��nA[��u�7mݺueA��^��Ql�\�`���tņ�gL��q~��I��5�L��	��Y���֚>����k�F��)yz��)ApTT���?(�xʋ�谰�4Q�۵c���++�q��Y,�$1��V�7�j�j��^A��+OE.�$pb6�@=�݅��hQ��s��Ul%P��|c;*�}<�����2}	zw��ٙ��uUJ I^0"�I2�)XZ!$����_�ٓp� 
J�8����a>{ߓO����c|"���L/�֒ ���=q��~�iZ�V���L�;�x�=�`[:�xs���k.����	�G�H'� �7v�f���,��:ˈ�?���J��"+9�/-��s��t$#M(3�� ��l�I�d���5k/"H�l2����(+�͡�(F�(-^�|tth||����_}��`$��O�%�
���?c��t���m�8���;v��kbb��,Y�f���(**����X�&p��DVȦfvu���ڊ�h,�ث�,�~a�ࢍ������밚��[W/[0�{�}�,��\=p	�4TV6V������{�w���D&�5�V���o����i�5�U����vR>pA��|v��P7�d��EQ޹cWcS�N�%I���h��\ãW������������&�n����]�v�|�����w��)�@BUF�APЦ�1�L�����`?��3�I� ��b�w����~�G?���'�7���ۆ����s���
\�Zw_=A4O5z�R��K��\ߤ�6S�v
gY�`0�Ri�@5�cc=�C���aH��r7�B@�M�,�M$R� @�!$��w�N	�b~��'��g�}��e���\���/W�R2�p9v/�_�!�y�m��C��&<����d�G��4<��C�]��h4j�g"�_�z��
6-�P{����v��F���#��
2�=�����j��x�@ҷ���X "z�$��Mgw��,m�hN���<��g	g1���'�yuO��DR�m1�T�f\�&��=v~{-�$Ds�	������mj몫�E%�p���j�m76�RA�O<u?��Zʍ?�PŊ�"��Uo����9�_��>ϟP��)�d2��� ��8��C�F��Uf�Y��ʪZ���X��9����d*Hӫo�]]]{��+C��`,M�3�gf�� �����`x��t��Ng[�'��(r{��C�:�N�o4����� Vv*c$0ZQH�#������%t�鈄'I�����*���-��ap8�dD e=�p8h
�l"�&ҙ��b֜�r�謇f,
�g�6�W���n�[�jw��F�����N83PX,�.�u֮]��'I�{������]�"�nj
��̥�͕���{�V�e��/���=�x[cSMy%�ٝ��:�,��C��4�z/��*�C�c�,�<�)o����;v���555�=.�������~I�=�事�i&�F��vC�N>�;��z����v�&���qN��(\�g�G���O��2��X��䤯��??�g��]]3mf�+��q��z�e�����>��-)-����K�P�7�e�{���=}aNf��Z&��?f�"c���8�C|*z��D^�Z�1v[Z"���U���x(�D��p�R�L 7@�g��Hj���Fwu��5�>͸V�d΅^�b�
�A� �L�i��APCh���/�<22�v�G��k��?e��>裸g���k��OO��8I�OP��q���T�GXo�!���JyQ �Κ�k��g��8����6(ʓ�L{W3��s&c6�A+��H$��x�Xc���=G-��Љ��������,$�KdYkS�@�A`�B��̌��xZa9ZR��Q�trޢeļ�N���*�E1����H�n�����e��+��l�*+.ѺWb�>)��D,��+)+��#��eZbI~�����'B+�h�8���w)��'I��n��[�r9�Rt��J�M��DG|12|��Z�m��m{�d���e�ȋQ6�5�m�M��tf�έ6�e��֎Vo[�UO?�����ƍ���"q)�QRJ���L�Ug3r=��k�:5��c$��O"�뮻eIY8w��_�|iiY41��/�L��o۶�?��Ύ�7���mmm6�5��F�-W ��2X�����K����N�a�����F�t�M��FR^���A�S{]�����hu��T�
+�$�i���t�*��,Mw���P�_N`����%��(��F���o�q���8!)j�2�6�d���� <V������𸻸��gR""Xp �d���1+Ⱦ� �F%Ɣ��	����;����\�Pg`�DI}\!Y�4T�Y��c�(�K5.�+�	PΪ^#%�H@i6��b�3�)Z��$���3������Q�Rm��8#/e�\�e�Q�!z��@��b�yK�'��N��d�x2�X�8��?������V�k4���?�ڿ|��=�Q�8K��Ȱ�葁���]�v���\�E��@Y��d �D^��d���(�i�n�����I%�H�J����1
��h�f�X2[�p 3��dDT8��@�M��y��iq�`(�r8�-D^P�� ���d&1���B=�X��h��\x�,gMBlz >x#j��v%���d2�كo��
�"C���v^�*�t�C�2A���"%��P�ѡ�&I�ٔ�Cý�.^1���� )�I+���v:�J�l���4!_u�\&��9§��TcH����1�6'ROL��꭯�_���{8���\|�^n��4]]�Q�,Kr�-�nl6-8�y��K�I�f��1`�[��*���4��;�������ϝѸ��~�6��F3��{���[�*�Z!�t<������R���lhhhoi=��U/���ƍ��O�ŧ�������y�w��=�I��~�������׽M)����Qg�WN-ٶk���BP�]����ʚ�g"�����g�N��I���ئ�#��3>��*ޖn�{�kg�V��O4ϰ�Y�E��
��yj��لfQ 1�k �}^���a�D�1h�f�ް��3=�{�E�Z*z#!`9�IU�H�y�2%J�b�d���>v��gt5�\e��'����P�H-�>��n~fӉ�t);"�y[��`�%X�d���Ͻ|�9�X)�Y���/��(��0`C��^�����X�2�mz<���֪��|ӵ,x��8�����v�O'��rN����������M�n9 R�?�ԧn���uG G��4�V���o��\�b��N�룊%��#��T�����{tӖk6\$J��Y�����}��u��.[ҽl��H0�J��!�h�6u]�n�`��C���A��׵���s�zઑp��n�&�#�6��8����`�(�B�Z,�vN�ȁ�� ���cR�Dw����{F8Nt(F5-�RU�x�t�COk8����J����.|�P�Y-�pU��5R/pc�D"�/��4^ Z?D���D���kht$����o����/���y�}Ӟdعm��>��p��*��9�%���JV��NJ3�Z�4i���3���i;8o�,o�F2��d@M�����sϮZu��ŋ���A\ g���X�SU����kV��>��_����|�x�6���R�jҘ��z_7�gaw�S���pX��Kz,�#���K�k��6c�v;I3�ۤo3��_fƇ$�O�!�x�,�����wX������5�u��l����+��X"�=qx��tp��M������L�n�ZtIxč��oIx���w �ؚ�/K�&2]��cdHW���fx�p�9�]���rDF0hh�p
<9��i��t�+�2��O(s�HpHY�����Ĭ[���Mq4�F{������{�̛����֦ :gUl]�G��<y�C[&�t�� )�D`~��0c��ǎHZ��R�?�L:�{��1E�D1���?r0}�T/]����j-b���k����T�e��]k%%���B��Xa$��V�t�Y��նm�Hc#�$�%����~���+f���:�� �c=�De��_�tJ)��p�֮=��Og^���7ܸ�k�(�ccc�`��>�뺦)�n,����,����0]7li�g�L�0��/"�L�p�,^F�P �*�E�ZD�f8Ӏ�d�^9�6��b�F���q�i�.;�+��NJF��	����#knnƄ�4X�w��]+�xk���Dc�F3M�f�,���.�d�OY����nhSƂ�x�s��X�id`�I����VK��e�cU�HX����-Sz��N�$�Qm�|�����V�Xa����ڈ�w��B���o��;��^���KyL
������[�愐l�Mr�n97l>�Rn��~*�D>�I�i\�L���a�4�p ʽh�0g;�	c")a�^>���͂}�b�'��+�g��u�C���u�9n�mЮ5�l�x��;b�O��M6 ���;��75yH�Э�$3�s?f*@J�y��_0t�P(�������"/��9v�w��b�}E1B���/�=��1w�� �g!s������,���*ڽ|��;zGF�/�;19�Ħ'm��e]�lX�����9�Ι��o}zO��9�p����tF�n�YI�(��2E�� �h�eh�n��e���~�A���^w���Y�)e���Ξ�9E��,dZ�����@�����vm9�c�6�e��!��ItJ8��X�x�/��pC����Ԏ�6)͕��<�j����0�ߜo���y$n���@VR��{I�iW;�V�����t���l�Z�yFI��gc�Q��1���9&��b�I��I�bJ*�ud��������'D��wtK�8��2���x��EX���i�'ZcT�R�u��D�BDF7P�CEF��@]�^�f���&;����0<C�[�@Q����d؂82��d�c����V�O�f�g=�IN��m��$������x�׆c*ʸ���rz��]��S��'!��KtDI�T7�3W�����c���k�b>O$.�`U �H����G?���}�+.�����Dh��X���cׄvݎ|l=O\>��NNN�Ò��v4N}4�PI�pD�:��c��Yx�2oDkg'vG1���i |Wk���w�f�_�FY�8�)�-:��j}��ܶ[|�m<,� �������68�sl�ۀH���\�hj��,R������Κ5�����T��A���4܊�|!/�REU$�_�Ď���O �U���ǎ~��;8f�ep���eY�m]tV[�L��}�c'F�MZF�UMU��Z���;��b�U׬�t��O�{u��G��w�X���*+�GOL��F��T-�X/G�LB)0('�ع��0��s��W8��Y�y�$�����l��6��l� �z�)�	��˙.[pi9��cc�S�+j��M��t�hv�c8�cy�y�2@X��2�d9�T�bI1��d��r�{~������̙����������ą�9r䡇���]s�o��#Gut��<c��/)�R�T�d��j���=��ug�I��Y_*_��̖]�{�[N,��𼳗t-ھ��Ï�ah������]ueKcC�**Dм���	Ծ��m�y:�A��N��xPӊB�t�UC����ZZZ,,}J�1���TS/so;��;�qLvbL�"n;�l�9o��� �+L��ܰv��D�2�tt
���Y3��M{�z�3n�f#/�t�@0��g�G�j�v��6rG?R���H���Ƴ�=��?n:t�������.zk��&�m���J���ym��.3FL������wèh�
�7��'��@������"�fI��rے ����9|�)�����֨��[�5���]�7�f�#$��<5�5�e��4� ytb��%jY
������G�jٌG�Y1Lv�WT��8N�����U�,ǤL�(�˲����h����)�qE@(,�O1���R)���	�Z���n��t��� �X)���b�R^�-�RL�TP^|�wt2��" ���� ���-���G�e-;c��|NѬh0\1P��}��_xʒ��! 'Gm�>n�)}�k=��'?~�ڦ�wI�m��{K�ܶc��prV��l���š��5���"�(�x�$�JѦE}�G?͔�pSg��&��
�s���r������/�Cck������}4�c�
y�y��/�Ab��#H`�7S�J�� ��^91�����PX��	H�x'2c1U�4�@�e1oƍy|(fEI���JeѼ�zߕ�{��?>�o��Zg����4�#�R��W�b��Ww�8�TJ�D.�N?���S��/���'�x�ч^�d��\��{���[��1��h ��#������^�����w� ��3W�ɉ8(�c *�����j��8|�g����֭/����\{ݵ��V)[��>���{/�Tt��f`'�c�ba���o�ޝ�XW_�Ή̌��[�L�_!��d'b/ʹ,�!�i�%@�T6s�W���pv��`)��;�02�b�7-�NJ���,���qKX��2hW���Z��MD��`�MQS�]K:���������S��ҕi�=�;Q1��T*��Xo�[��zI�������t�զ#�j|'�0�Z��X���+V�;�Z�7�j�����I������PQ�}�g
�xd���j�X
|��O����xz2��u�|5�g&�'�����M������c�洵-_�M;����v�)y f�s�2������O.��Zo�urb�O6����}蕟l��6{N�Yga�U(U~wߣ�_w��aZfՏ��g�|�����}��b��Z[�f��\���1�o�G�^L�u�Yb�=_0�����
�X_~ϔ@��Gɹ?�0�e:�,
�Dr2�Fb1�����G�#�}�Ű8���t����Ybx��!Eՙp}Š��ECD%��z����$q<OX X.G�6�`k+:5189�ˇ�.�X�b��١�.[~N������G����I�|f��8ײ�d�I|a�P�KV)�����vM�COn���}�^�61����}�߸�hq�
��i��#5�ո�]���
vDę��Xdg�S��3o2NrY���R|�������D�W*�$��	 �6,�o �������<�@sSۭ�/�8	��(�E���l�A��u���L��F �h8.2,��뮽n��=@5�ٌ�X������i~���ܐ�&<2���eE�5Nbie��Z6�F�E󽉉��g���З�������^���u~��̪���0LM3������>���/���9�����Ο�7d�,��bk�K7�2�#�]#��}n�MWTF��4�8��9��#]H�Uq  �[������O"����=55ަN�O�I�z���	8s�"s�(�;��>0�$����ޢ���R<��e�9s�8t����y{F*z����_C��HHض����|{��v��{zw�9���Ҏ�_�����wՕ���˯��^�^���%R�{~qo4$]z�z8���;���l�����.Xť�i��"+�Ӝo�[@|E�h�O������@���L��?ГK�s�mݼ���/Z;oa�K[�{��>�ћs���Ç+e�S��d���k�k;>x���(𺷭1>zlpbbܥy��l�`/�U-��|^�ss�K��������R�x�X���拲�+H20�o$�2248��[)":���(�#JB6g���ʶ�-m���d*W��C�(e���z�\#�MZ�&P$�A��o���?�Y}��˙���:?}y}S�����ܸ���Jn�D����/i���8%����=���(Ա��������ݏ�aÆ�Y�艾�d�5`��x+q�{���;��D�|m��ۥ�٨�Գ��ݹp�ˠ��m�2e��ScZx����H��VZ7t��eop|b�?��AlQQ��,z׵��7��442!�o~��?�%��j� ������&�ɖYq0=���%�־���/論ʀC�L6��G�G���9>1�� C*�I��ǸA;~?JM�=��UMy�1�UK�ӕ�Y��6�v�3���e�~Yr,��8��)�*�u�j-m�.�x�c�W�*���Չ��Gv���x�-w&�%I!�a�=��EQ��j�Z�.���+�*��F`�����Ӄ��L�r`�2�X�\��f�]�#�睚�=]�������*�BC�M��GHZG�7%�?�wF��qC�,�Ө6�	�>�U�,|�[�I<9^��rm/��cNs�ˣ��3
m�B� 
'����Ϳ��m9g�*9��;z���6S*h�*���-ϝ��,��ޗ�T~���O���w�,k��J��������\����]��G6o~����g9���HdIM)�{3ã�S芩���:����H���L#b�T��M�^}�M�^��Dfss�}��gxx8�b����}�%�]f!�a�\ˡ����1�K掾�����������Y��vM0�z�ߤMC*�Y<~�E����쑓c�JH��K�@����t{�4����냃��1����gxd��������)ӵ&��8�]�B�ԓ+(���㛷��kO�#���2k�n��4��4H�@���}C���Α�nXw�\��[{�+��<�g��Ez��p���xD?1����X���ༀ^(�����X�D��� ��."<�ƽ�!�5GB;O��`}CO��a�9�>�֪��Le�H��D�Nۚ@���N����]�y��g,�B���89_y^,V��k�����0L�ڎ�=���E�����c�G����o=r�����:���3iY�R�X�㙅<[*�.���J��5"���E���,q��w/Yx��^��UU��,������ph�ڵѺ�H(�����_������A�o��k�w����B��ހ�,�2��
���N]7֭=g���'zz���B0�ʂhۆ�Q6RH��6 )���ɤ�V��n�={v*�
C�"�P��L,��� N��"%��kQM��M��M��4	�Ƌq�b���QoӇ�g���(���cz����x��4n��.�?L�g�U�Sע�4�V�Ǐ,Y8oú��`Q��p^�7��M!�P�X	D���կ���7?G!A����v�G>46��P����}7�_x�9�6>�p�R�%^�D���>�Z	��/�5�}�i ����FG	�s��2��h���Lv����bS��?�[�jap``���{x�Ý���\��+�2�şݴ%(I��N��(ȍE�69�sj����NЌ��=��[6���1��q<'�B���E�K�H�����&3i��[�x�
$yHk�A����V̾4<4k��@q�q�c	����ʶ��(�V5���7ͦӹL��!z$F��n����]�y+4*�k}Ќ$�:t2�=��+.^h�h�Yuqׂ�&G+ӎELMf�1n��UW]���U(��7�����7J��#�'O��	*�ԧ��Ych�L]�0��/^����+�,�	pJ�"�e{ZOҙR���n�m 
:z�Z���~��腔/(���%,�{m��P3������o\ؽ��(���_xɥ�+Ƌ�{��k��D��͛6=�w�-S+-[�lx@NM��?��f۴�V�x<��8 h!��L$݄�˟x�cE�_�hQ����"�0���^"���f5�v�s���?u�_|j���@��nݺf��O�ze*�TՖD�44�6Ik�������G{V�X������g�gw��L1�.�|�x]�ڲt]�q�em�jU��m� �����>{MO�*����X@�q�˚|&�� �V��D�7)얄�5'��u*!HO��N��"�E��?���_��՜Z�IL3+h�vM�R�$=�a666�'~����&߉�x���Z�_�[��SWw7��eEi��^G�~f��K3<'W�<�����"�b��斂A��'$���O}�_��/<��+e�O�lG[[K[��m�Vh���*���G�B�Pp5i����8�7| |����@��,r�;iѴ6K�X��2UU������J:Z�MQ>ϒ%]�فx��3ޏ�Ǵ��FG�{�n��|GW��2-��ju r�gRC�O�I�S��������Ԑa���T*���D���[��,K�L>�կX��_�
��r�
ࡃCOڡ�"�<�9�;�����^1��Ȣ�M�� !EtېZ6T�3h�0���m����mw�p���ߪp�����H<���3�<���xΊy�r5-15�B�N�]z=~CE���>z|tx��W�uuu�㓲(�N�t]��f�0��et�F�;��x�p�����,c�ڍ����@h�#���I9���bVJ����r7n$$�ey��14�V�n�,{}��/,�K��7>{Ɗ�m-�����.\^�\��l��mj�J\�GoQK�\>_-U�>���4�׿�ҋ�M�8��б�MYſ*�l�h�9��$��Z�	ep�m{m�������׷�\�u���a&Xt�O~�������.	�"J���X.�L��'�z��o$)�� (�C`�Ȝi��n���L&�Q*U���_E��`�{{{7\p�L�X�~c��Vzf�`'��pe�\/~7��ަ��D�hҌ��o���ߵ�*E���Q�/Y�TWT^�(���/@>�� J�,�`:::0��wғ�I��4Q������CA//��1��?P�2�'���7�	瞷��G��7or��K�pR�Ұ�C�n�Ŏ0PC�{=X�{*6C��I�*��S=�ӗ���X;����4��,+y.�=�3oq3� ���c��G-Cw��6��'�����ක�v���brr��
�4�􂿫�����������f[�И�� F��L&[�吅U}�7��mܸ��k�ojiUT�Kthr ��׮El|���є�;X�4U������q�VdG�m�P���í]6`�^�t3YX֒�������F���1,�x�]������M!�G/U	�֜V��0��?�ȳ�Ͷ���SY��[8M������ã	��j�ĺj�c�"�f��GƇ��$�P@D!��8� �1��:�HM^�� 7�ԕL
M��JR��q���%]��W5U�ʦ��Y���<��i���.�d��w��/w��W<�?�kVK��S,�>vh�E~��m���l(��.��ܻ��gO�w��	|�_Z0w~�\Z<o^8��|Ã}�R�Z-L�B�����Ǻ�s��eW\�M�����������8ֽp�矛ϖ;�Z#�0/JUc�S��,xp���8ǲ�x8��� �
������b7#��ʥR�T�dRe��D�8O*�Ȫ��a�;�)z��pHS*����Ȩ���h���z9���6CrŰ7pJ�rjU����f B���f��N�+F�ƍ�
� #�!gM!h
ɟ�F$��\�7�iѵ�k��շ�!�[�["�V���l!��.��!G$O��yU��d���[�x��4��9�e���x.��hF��Y�7��̑c��f�w����o���h>���՗oH�������ܑ�t���Ö­5���Xw�XO�9��ͪ�F�A�7iXڊ�����n���u�k���Ƅ
� ��м(���nݺ�k��A8�sx�k/�w��$�t�yg��/�h�n�F��o�p���H	ܛ7�i���nddDU�X,�I`Y�i����jUQ�UY�}~?�ݚfT5]U���'�������qu	���'�Z�t-l[��m� ��_VYd��Fô#p8�c�ł㔚LĂ~8��1���z`piK���ȝ5�ƈXb��.�	�m�P��R�`����P\��$<���mW�R�����X�EB��`;��X�1�����OK4n>ú���8)j�!^Ko�SJ�#p��z��K�TݠdbQB8��acߙ��h�Rt5�AS5��ڬ�]w֜�p2�J��#��P��c���Ө��	���s�o#=>4�ד���I��믻��ي_�`�"�� U�> ����K;��e9��t&���[�����b�Zx�	 �L�\c}����C;h*T�xe鲋.P;^�O�kJjbT��7_)�
X�U���$�Ŕ�yp����3,��q����
��s������:�,PfZ���Nhq��S�Z��J�������"�����[��vN'�kDv� hZ�y�ЮA�e���\!&�����1�<@F�%-�M�a��@��ɣY�O�S�a�t}C���8�-��w�4Y�b�6ð��2�<�5���.}�r+ql�z=��dCc��u�~��_t/�7�/m��/jo����YM=�VM�ƫ���T�Gn�!8U�Q���y��O���J��}�^:�ܳp��}��S�ܨ��F�a&�~O&<�����a�,+�M
�CR�0z�
�W]u�Ï>�կ�oe��s�[=n B8�M�/]� &Kg�ݷkm���0�c1��\��7�o���ñ��L$��ͩT
g�ި�B0�^?X:�\�V�Mf�t��7���ˤ�����<� �
�(�7�/<�¥�_ٵd�c=�@����m��p�����vJ�c�^�^�:C1.�R�-�pċ�j�|p��n�a�!�D8�mϛV!��ś���>u���1l�LE�1O#=f���m&�y���`�&F�2�L)ӄ�[�/f�<�� @࿈�E�f�2�/�=w�3/<̧�zE�K]z%�-Ui_����J�-Q?����mi�&P��*��$�"��x����[J����U]	����u�<-�T!�	���~�=��4���%>����容b=�q���P�_�㋀������I&�N�O�W�������JE9ٗJ�O��,����z^���	����� f�nCG��{t-�h~z?
<��V.��u��^�i�,�DH-��c�Եr����ݚZV.�Y�d9Kq��	��S*U��W�o�1�̇O<o��=�,���֡p<��z��R�N2���dXf��3f56;�,�ˑH�&���Hw�M[4��#��t���&M�$fIk��Ű�3��Eb��ã#�Xwg�����:`�B
i��g
|��H���eh�TٍӱM�ߌ�"b���)�񐦪��9Q�DQ�-�����\.��w�B�8`�RI��&��Y��w��65>�V��eܱv�P*�
�e�������Ƈ���Ƭ������������~{8.�n�m�W{�a\��?�+�Џ��;noG;S|���rٜW�<Z�jel´v!QnB3�)e���?}����E� �3pv����G�^��P�
V��+��~�i�.q�$q��1�y-=4��{�Ot�Oݶe��wlݞ��_�1��V�Z�9{~����e��!M�dI�S�n.�Z.Ѷ14�<:���zY$
�������TF'�o��V<�-_��J�s���B�_):U�j&���b�T� ��+�rn�t��&�ओ?���,M�����_��q$��D�g�Iǵ���T� ̐�2�^�2�tG�h<��1�iT�z�ek�Q�|��m��8x�����ޱd������٣���� �X�q��Ap�5� �8�j��&�6g��ΈΘ�by4{p��U��[��3q��%�3��Bv�c�B6UĖі%���m	X��v�m9'mX�_�;c��;X�|
���F���7=���y�,{áP�hC�����ͱUU=t�\�ѣG����O^ T�r��^au���z$ H�TK�O�6�p�m��j����6�س���޿c��ÇO�#\Z�FH�~�	gϞ}�ȱh�>WȢ7�F�=����8��E������?B��ħ>���3�To�,�uߒlE�b��\6i��3�aCQ����:cUw6�H>79t8�_>�1I�֨�o�J�lZ���HM�ܟ�ee`�K�	G*���P\���ؼy���8�<r#�2dҤA��׻�����Q��]|iCc}&�v!vZg�d��g6��
m���}ve4,�|�r��Glim������˟.��#GN9���L$�=^��R�hpK�U�ma}�%�]���FѬ���MO��7��V�](��u�Ӌ��<[�����8��MO�}���֖���ўc�j�X,f�L��*`�Y
����M��+�F���B����T-,\U�K����Ϝ�]s�/8d8���/\� K�7\,��\�4SK^	5�<��]z��Q>�o�V�L������������Ɇ�f�]H|e���[��vd!��t��lV
M���E�`�5�8Cb���<4�b]�q�2	��Y��%L׭����QF��dj��"�*������*J����zeA
��c7���~�+�J��y����h�-L /C}��Ǖ����Ձ�\^�RZ&ki��۔�(��O 5�XO57y�����������իW{���O�"WRK�ñ�=��$
��D$����RS5��G�����c���Lu���i���@����;_�X�KU����M��t�ȉ@�t&�2��
ƚ�E:x	�1jǤ�L"VW{|��Zk<<��,"⍾����?:9���3�$x0����4����dk{ !	��A�<5CQ����T8�H����554\��xn�6]kb!�Y�S�rxiHǓV�.�g�����Le����q��cMM>/w�� \Ƃ�-�C��p=��ς�P,V�e�ǲq�܍�2��s��Ę��g*q��8 B��}QޅJ�Ҏ;uC�*U�#�.���ȕ�Я�e�` 4L=�˫juddH�~�C2���	�+|�����|��M��1/��^���::;i�R�$c�����Jr��C��7
�M�x́��4���� ���ԥ���9m�<�����1�^z�u6	e9nD�-�}���@��,�&��"X�(��9��?>fe���J�w~��?��ѣ�񘗡e�$���㓩ys���+/=?�?yr��fN��|<��4�P�l���xbҴ�Ɔ��b��>8i.���g !\C��,[����������y��᧞|:_*�%1ϙ�����~e�k�֜\΅�,�֚�n#ɌZ�!US��;u�i��sJ��&d��.b�lW���ʪ�3�i���}�,�v�&R55p���iY�)6<�}Y�M�X�e<c�C���*�m����R�ů~����g����_��u�s�b%g8�(U��f�A���ٷ�F�6
��BJ{��d�>�
~�020������{����^��ږ�R�&)�9֐E�a��"�A�+m�p��������i����}���hO���oX�|9ЩJ�:1:l���`�+6�w�#K�����p]<����BՄ�Ŷ�!t��j:��*^�/O��>`�8�Fc��܊]k5�Z���z��- x>�W�ews��G�:,��z$�H&�33g�+�74�~
����L]�Ȃ#���.B�k��a�!�,��h�\���}��:P.ⓓɉW��`���(+����w���/��{�	��i�>| ~�`���~�7-_�M��1��(��J����U����a��L  $��6�5�s�]W�B`��Á`]}<�|�P��D)C�Kl"(�+�:��͏�sK�5�'J"EM�J%�W�\ܶ̙��H��x}r�'��	��u��J�-J8I���ߵc;ˋs;��N��r����������ΙQ�^Tڞ�N�Z3�o�!� �r2�����[QJ�XСUi��-�'A�?���F�9ټ��>V��ah���Ҟ�{��s����w/�:�v�\6>?�4�P<��;��}�n���tS����i��������h�B#&�[ZA���+I�Ϙ�PU�_(�ps���d2��^��{��t:m�0
�� 2n��Ӏ�)eY2�\vA9<P���MѢ��#5ՙ��J=7G�ҧ��G@��f���e��ju�X4w�d���L�d�׵���\A	x$�R������K/-?s��ٳ���h�����? �?������쇯�<Y�����y٦8�l�j�@q<˺Rt�RU������0�ܸH��b�������|���j��ö��b(
x N/�<~�'��Bح��1��:�΃{c�ȶ,R����k��Y�Vu�3�}�����P>��U�\|��˙t>����/T�fc��ϋQ-ֺ �A|jǁ��L��y�h*��8K7�l>�v�₁#�>!P��U�R�G�9��;w��E���W_}��Y���G>|��x��;w�OU*e�'N���
���+M�:��c��r<ǃ#EJU�;_�7�pNO�4�j���O������r�o�od0�8��?�
�Rm|��/|�A%��}׮��o�������J�b��xb|ђ.�0���Ax���'�o|���&�����{�Ǯ(7�p����'K$K���,sb``M���wU��N�Շ�y�/���`_�󯽼x��h2L�[�F9����� c-�].ep��L7,�1p�ਪ��8��i����r��Iu�^�AY�`Kp
,'0@�����	W�̑L"q��{���*����&�U�G\�f����~z��cG&Y���AUѼK1�Ɍ@3pY2���b�����(ӌ��b>	eJjo�@���}N���J!���ＷB����?�hW-{���;�n���{O�<�U��9r��/R�VO�qG��ym��9N�Џ���$�}��r�e"�K�p���z�L��j��� �P�,�*pа}��L�SIK7|���HX��F�u����G�������G�u��d�e*U�T�Jn	�T$+U�p���^۝�FX�^/�])U�岦T��p&�Ťg��A�^3a�f��Qo�'�Ʌs�s�ㄒi�H�328��R��d�T���KE�f�&˖.�8��4+��X�gS�p�ol�ܖ��رcǶ��IT�>V�����2x41 �hbP�
<?Ԥ�*�ɯ8w)c�����������^p������s�������<�w����-���u����7�՜���JnނE8&Ffo���?�Mf��-����o�Ysֺ�{������5����ż��*��􈞆h�>&]}���]�x��Y�q�@�E��c<�,<������P�#pX��uL<{^W5���Û��f���g����nX�nM�����/X
�Ӄ���1F#���r�V�odh�$k��e�`o�?�(���|�--sfwtvvΛ? �P�%�p�ʗ�;�^}& \<�zpY�\��ཇ��=w� 	T����ڞbx�0��ٝ�HDp"Z >�ɱ�����p0#�+)�=�y��[>�}�k@�O���jR��hb�&�8%�N��:�opmg�˛���rh,`o�x�+Fv��O�;@+@Me��S��ߏ$1����%��X^�YJ�����s�\&���rH�I;
Kat��v���:nҥ�� ���;��g���pFr��jQ�ph|l����ҥ]�q:�N�\33o,�BD��r�!GG��ж�b��?l�4`u@,�8��kWQ��ة�i�4�{r9k����^"��Ea�"<5�����'�Kr�P���8�� i��7�iN1`��Emx����m�b�ho�чzd"Y*9Hdxw`�C3..C�j%��X&�t�G� �>�?-��h��G�Y�r��C��M�'�'���Y�W1tMj�����d���e���yl"�+h��?|���Pj1��`EQ�T��Vf2}�����[�`2���T�,�e2�E�Dc�L.�������ګ�����~��<�5Ѡ(��+/>n�˻��e���14�O�ƙi|<e������Y��y���'�wr����nt0�dI���y0�p���_�p��`����F�X�x'V�K�rC���H-�v6�:�F< �yVhߑ�CG���o/
�'�,_eVK+�����y������͙ϱ�!�<�bO3Y��Z�, hрNQSs)t�С3�\	�<B��R^)W���k���)����狳�jo�@��2kV-�壷������` P(�d�{��utt���h,���F��@�����Q1�����+E��E��,YZ_�ݾ~����v����$�%K�]u��{�`�ED�/�*�b��o���g��^6A�'GV.[���1���~oSS=\L6_`,=p��t25�Evx>���rҀ��pٜ��x�Ąݯ�Gj��O���Դe���3=�b�I��I`�q���ه,WR�$��Z����<k:�X�TQM�fJ�o��p�<gZG�H�!w�M���Wlkp<!����O`YV�8����@���70�79�0\v(�}����f��;�լ&	�$:�*�G5pQYEu~�D�do����zo��@�g.W���:6�鴨:���6�FLSC����㓙,�#*K��7h	x��E���9x)�&���P(�*��Gy<.h�;��XO<֐�ꜷ�椪�<�����9���u2�ЎI�Kf2���^�xt���]���@�Tˇ%?��ʦu�xˊ!(m��}�X��R�Cd�:����8?����w����`�o�حs��9�wϡC�zO����:.�ZH쎫�HO�"�N���6����0ry).X1�����@�7�l�j")�����"8��i&S)��k�Z��O|*�o۾���ζ��#g&�#+��)v��m��gJ��@9d��E�H:Ӳ��b׼��]������ӵ����тyK�����h������d:cY�\&���d&��`ֲ�ɦ�:�����QE)��X�;D�dM�ѭZJ�'��X.]N���]��5h&�=�~6��:�w|$9
�!���/T1����]~�_*k'F`?��������]�����)�4(�f�$��s�;���󵴵�:�[%�0@�u�>��G}���O�3��]��k��f��=�����5��#�O��' ��j�`���P%^X�|ygG�{:.��2��)��c�.��`���,x[�������>��N�� ����I�S��Q�W_� H2��H$�E�Պ؈(��;P P��}{�.ZLj�l��Ɍ>���D����Д�k�oDd�QM̴6�	�����fO7\�ib��(x��L�E��Xșf��m�21�@�3���=�����T������i�b~�?��m��u�%��$8�-�L��8x0�J�@��R�ع� 
;����ۀ�$2��cׁe='\EU�e�q,��7^��i���?��� ��i |Wk�Q�Y���4�{p�9�A�y��̓�UՋ�B2-��@s��w��ɧY�і�<Z�v� �NXMÝkʗʹRi�a�h( [/�Z��ǹQ'��|��g�{��+.����{aG�e����_���;��ϗ�`�D[d	�6�a8t�h���!ґe�C�u���)���{pP��X,<204^$��ح���j^2�;v��韾��ܴy�_��뻿|Ƿ_��* !���~�
�7���p�$��6j�6k�U-Ÿh�c��MMM�����g�^{'0����@H��fw�W��-�H����׿������}���Oߎ��٦m	*H^���_��{����������g�d"Y�g��xM��NcCtvG;�D%�6}�� �V,�����O<x��6�ŷn�����I�L�Ӕ������Q@|w!y�'�~rŊ3�uM�Lz"���V���q)���-���q9%���g������]?���~71R��m��lu���ʗ�v�e	<��O~q���Ζ恡��xý���C��b��|�������}�T+�RM�/�?���)�J!<,�lhn+�`ơَٝ�BIѬGN�8���C���o���o�<����䫙���M&R�B���aV{9�� `�7���3��M�p(�����<�]q�5W^y���S �Ai�m��U�V�������_�=7 @ �����X�!��ܺ|>��wr����Y��c����M�_WU�s֭��s����w_��_/����=4S�T����2�8�����ǰ�Í�cOm*���wÑ�T�އ��'�M�L��X]�(��e����Y1�V�Lf�����	�R�p(K��c"���<��b��rjŲ��*�N���Y���MYV�@���d:$1"�h���{���:/ЄR��p�LDL<��Y�Q.���RV��J��,@HJ�$N<�̳������*��4�K�oZ����\�S�T�@4��=���ߞ*$ƕJ����t�zx�,(��h�t1X��&�ֈ��C0���[�A~��!�#b��.��g�M��viגw���I��tM��Ui����ށ�D2%�HE�f���d&�>%/
x��H��ܶ=4�5Js4�{���Eqhx�����6�sU�r ���TZ��W��-[�L��8F۞Q��]��驶�#��tX���dӓ�>�ybtL�T��F�E�LA���xSc�T�~��[2��K[���ͳ�+.�!�655�;�{�L��LbM��5R�c���,+abif�� ~8XM�~}�s����?pY,���\�\.Wȗpo##���?=���A�x0�в�k١�eٓNe&��E�xA��Ϋ����B|�88R����O=���^{��?��@�g�ڕ��;���g��m�\^+�QUeVC3��tV��w�}��'��W�H�w`�2l�8��<�g�[�67�77�y=�X,������&3�C��y=�c=�p�^|a+'J��w|��!J�-7��*<UC�nna�L�uJ�C.X`]���{CA��'q�;b	Qx\E���c١���;w���̮L.[Ջ���ؽ���'a7��,	2.�tXW�F��P���V�f�v/IL�),��tuu}��[�Ѩ���$2RC|y�2�຀�~͙+/��x0�c�\c��������z�i����I�4C8�:b��mV�UI������A" 6�q" a�ݸȝ)�Γw�/hj�B�;M�g��+w���'ҩ"��Yu��,K�I�p/�Ò��0(��)���;��A��e��kj5�$�<Ⴉ�|���W�������]��:��j��`LOx�h"tL��W\u�O��jz�.�J&���q�dʛ_��۵V�Z���:�b����_41�0<C�A���C��6n~m�ο��/�ʥ�G��őN�+�������~�����9ŵ���~��L�B�^h�m�C�T���X����!�]-G"]��v���ۇ��.���ϗL�{v�~��u��`;�,�;����㡚���A��6S}���6�5^�pA:�ٷ��-[�dғ�Ba���g�~��$YOLn{�u��Lf�Pյk��hS�e�"��9�\ �޽%Ж��
a���d"#{}�p؋��j�L$Hq��XS�[���y�����bف�{_|�ɾ��@����Ʉes�N��O7�4`��x}Ӊ����E3Z�]�H(`�Trr�sq��7}���f5��L���7>����[o��%/�|r���9Q��#(��:����_����n��v�ǉ�	UU�Xȴ���8<��{v�����.]�1gn,+��
BX��R}�m�,��r��d*_X�f1�k�^ߣ�Z�qUȝ��Ra��&Tk�!���	��s�"�tA�ka��;��"rxU1�[[�&�,g�N$�����'�J(��d�̙�	����UUCX��aaö��o�,��;�(����K��?g&� �s�iiUS۲<�[�R*ئ��nu<�K�aƏ������B��a��6�����I؃��P���D�tē_o-2�J
� 	�ں͵���Q`1�^��M�hjy:,�F-�E�:;S�e�A�ݱx���i�NE}�w�cn�6G�D߱���4�:����ڽv�J�:���=�N៹Hh��e�6,�tIʒ~�]��i�j��w�\�y7~n�3wz�^�Zu�P$��D �)��N��%�6���K^;N�7�c�q7����K4u��w�E�w�Ͻs��yι�Z��7�|�3���r�9O�_D��֨����@��k͢���x�)������q�R1y!�,�F�l���Y�m6o���/�u�MM�C��&�=�X}]�mY�J^�������	ʴ���*���as�����J%YV�ꛁ񘪭�#�M-����ϿjêR�.�5k/\���MOo���_\s��i��^�]�^ޞ���C�50��~Y���_��g��~fd4���@���B��d:ŋ�UW�>�䳷}�z�*����H�p���)��s��:ٙo�pdۮ��	��{��I� P���N �ޓ.�Y��`-�`1���&�~c����������o��� 뭾���ڶd�ylx$L�#���Œ����wz.w�)�,�4u��;�뇆K��;$9��fa�����P."��8�pA�9��HV�s�26N��#y��gm�̙����u/�;�c�p
N�ܼ�M5͝{ޥ��EB���D� �X*�6��E���x��M-��{����=|���'����Ǆؔ�V�R�C�Ƅ�up�`�!�[���ga��h�loE�a��$�W]��ZKk��7_o�6m`����f�8�JN�'�RWW����]'Ouvt�&B:fA® E����g���|�׼�3͊�˚��IF�c�</�dJ��i��3�
G�:���U>�/d�{�$�e��~�?�Q��&
���b���T����-$PEL�2C�Q�w�6e����C�l�>�5-�P���#Ԃ&:.l$!�(U6��]B�d�i�
�#Lls��eNBg���שr���[�ى�.Z�s»��r�_���:���	��zK/Ofv��9W7ÑX���=�4T��4d���тcw�$�kQGAk!A,�ܱ���l[��,�{M
�b-!]]���՗^�}�`���$��2��R0v�G�uH�<g��d����M���8��HL$�o���w�����KJ���Z�T,��-]ڢ�5P)�w�����/5����R��籂;Χ���e�����a�@�2�0,`���'?��z�u7�B"]WkYN���gcc�� .]�C�ܜ��A>rS)�т�����IH\�(�0|˦�%�h�EPue���`>Iij@)r�l���UU�]�(ꀀ�ȊN��h�0����KW��Ϛ1}dpT��}x���������<������[����j�Fcc��^�윝˖0_�����F6o9NZq+��`�+,��F�`H���z�g?�i_O�,
_��g\�D�
�n��ƛ��Ľ��{���t��NٱcG9^Z�f,���03�;���?2h�*�X���jp��O��cT�vA����&k�H)��Kl�D"�#�u�,z����X]�C�x>�POm��tc����C���ޖ��&�Q��^j�qsf-�7wq0�BZ��£��ct�k6Po��K���X��߾���O���n�6��_�;�v}�����%�����/���/��;�}����x1o)AY����L&�s����B��P߰�⋯��2�rĀ�����aV���/�!����Pyl|����p�9�)����v~�5�hP�)�-c�r�x����d*�,8@&Ƴ��eY�h���AE6��%W)�l��W.�`���[&El$(��R	�f[t����L<��8,�D"��ea�cz�)s*��\
�`�ƀ���� (]۫�3���V��9E��&�
��y���Ǽ���~��+�V1ʆ����S�i$�I���<כ��G��++bű�+ V2ٌ$8���)��׶�ɿ~��hD�@4�C���ᔀ�e��o��\�*u����*$B����$��Ш�VlL3d�\�XW_��c�����p%�.� 5/����HѨ`��X�P��n�Z���YX�z�ϸ���	ey�oDWh��D,& ?�����Dl���.��\��F�J����l�=?�6�9sg�_qE����JHVC0��ˊ[	F�$C �wGdT����SN05	~[KS{1���<h�x2Eh��l�2�J��-�����<�}�wv�D��fl� ��t/^�č�
Żr('�»%���F�H��$���D9*`h/Q����?��Î�̚;kт����_�w�����f�\��8sz'�E���}*+��� ��:օׂQ����X2u۬N�h:+b��O��z	l�28��BZ��84�!j  K�Y~�rU�{"94��� }�[����G���ƒ�Ǖ�-��T;qa� V��듧�*��"~.q\�
��Q=�/�LB��%��9�yz�����%B���M<���p�?}��\��3w-,���?x�7��=�]1(�`BuL�ڮ#��\:���w|�s�M�e���/��i]�d��}��[�����9���&C�;���9�֡�J�
\�*c7��k� �X�,�I!�����D,�E4�<�g�K��4�$W_W?�-�~��R$+pt$[#r��_�p���H&3+v����A�w	f��KKQ�b��2eb���Nk��^΢J�A��7����.SxN��A�<��]޵<��'w��d�
bB���ACCI�/�f��U�N����;" �d��b�@�����Y�I[�Uu���M�u�Y��Y���2[*�bɆ��(��^D�M�.�J�u	��21/c�lAN�P�X؃�����s˗-��ʖ|!�h���f�*�Ȓ��57TJy���
)f�kS�u�W>�_w���U��>e�/g����7��}��Y�b24jģti�Rp@��f	�y�(�X�U�iZ�����
��+/Y�J���(i��x�q�N<����%�lڶ$���4\�`�(r�#�P_��մ���
�(��ؿ���lp��� 3\�2KR ĝ���?��ab�G���|����R�rA'�����';OX��p��F�X~��׾��/��R�X��/?��CXX�����K47S��Ǒ�M$U���2E�E�tMS�T��d���
)EU�0?�زY�6O�������b��-��b@���BIx&�'�.+a����&A�yVG�򘚝����x:ܲ�ʁ��K:��0ϼ�S�>V�`�> �tq�6YV�U],�<�%�������v:5�xњ�jk���C��._���9�կ~���oXc#�H�{S&e���M��4Q�U��G.�p�s��8{�̎�f�w����39��������[j?t��u�1n>�������N�Ӭ��S����S.���/O��{����`��m6��D��+����bE�f&@�1�kH|�
g��5�(O��d`w�`U���o�n�*b0�' Q��e�>".L��?8�"|��g�-����<¥�������\�ֽ��
�̋�W��C�?��@@n��_����S�&��l"�#� �t�^hqr��t���DPc!d7@g��B822���w����Ͷ'�I��wܚ�����0����BXF�t��i�-!-�^�ݑ����jZwO��=��kVJ�hkj��9�(����T8,e�%LiVsK�����.B(�ZM�L`2�����
b
(�bѯ݀y�E�������P2s�b��Y������ֹ-�
b��Wt������g̜�����Бc]]] OBZllp���v���n�vI��G��p$��8R<�ʁ���W�[r �2������%L���`�Mv��8PZ
����F&U�d%vH�C�I~b��6�JFW,k)VH� �m���6�吥\4���b8�!m$�#f�K͠°�S$��9~��ї^y}����io�\�pq[۴����\�J����pKK��K/-��ݻa~`6Z[Z֬Y�k�+[���mJ4�����wZ�Oѳ�\�f������ɮ�MBMY7_-Krȫ�� ���M�yUK��3�SB)o)Kil!7���W^����[K��W_3�sڲ�+��P A��e�G��S)R,"����X�SHmcC�E�
��p<>�g7'��o\���o�O�I��n��y]�����7�����7�3��1��R^�Jolh��n��ԍ��v(���[<>_,1�)�!>���r z��W%��p[{����x�w��;1�V�Q%d:ĺ$mn�(��"`���k�a���b�R���JS��'C��qN��1���a�q�'tT.�r#�ŤHiij��������Q�$����b��&4̤!c!�Nb�HL�:�rBPV,�eZ�G�U-��c7�J��JA����T�J8k2��
,m�<��s�y��a���XzP��$��v��%~����`�b�Œ5������S�Z��>uP��='�Zhbd0Y%�̍�V��w�6����D��{/�&�k�U��0�؍N	��uɚ#�n��E?e>'��?���\*�(n5�
���]a�[%d� -@��\
�[`6������	�����|������ׁG����ƶ���O}��9::R�S����?p�U����<����<v�W�Q�/Yq�����l��6Z���r��[�j�U�$NU0���*�#�-[������=ڿ'cG)]J�	���8�*V=�����M�:t�0"X�[���+��Bmm�Ç0�
bѥ�8f��G�I*:e�4LP*84�#ÉfϚ��[L��|�Gl��O�����ck׮3$�L��O/��M-m555�t�?���w���[��?��������'&�_��T*E�P(���ރ�9vt�:xd��K_�b\���h�&�F	��*�4��i�?^�1tM�"2�V#>2�˚:�����8̩��oݾ}�3tz��{�����;X�;P�:�5�jx<CBa���^�~�M�LB�H}�et�$�ddhd����K� 	�"��̈́��^q��u�C����?2�W��e)�	`ը�Wa�$E��E���؜� �CC�h�R7�a��r�ڥ�G�hX+zNH���bٲ\��P@���>��ҼpѢD"1:2�ۋ��e��DM��3~�exth����9��/��FR�F8=v'����~"Sh�eX@�|5R�0z��)��3`i(�Ϙ� n��Q�E�rof|�+/Ϛ=wI0��fs��8�z�D1ArK2J:�c@b �fϙ�˶��|__�,��0�"���j����IFC�d�"��M�O0Nt�O�S�2���V�㰱@}F����[�[���]�"�����b2��%5
U���e)֦��b�s)�6(g^1�����Е�pD�dd_�>ȵl��	9�W~�9Bo����>���U�ȳ����I�6;S�4Q�\I�h�0A!%(AN	6W	�2����#'������.g���ۺ}G{Gg]CS��k���-��ف���)���|͚���X����}������q��D�Y��Q��:�b�]g�{���ǛeO΀;��ܫ��ĶJ�����+�@,oKb0����!�Hb�OX_��NQ���\��BI�N)-�7���+v۴��n�1�)�j�?��?z���Pմ��K�,��6����-B����%K֬]+�2�F�_�uQ�A/Μ=+�i�D�����5]h���2~���!ό�4�4DY
${��Քh�#_��`�/�6����j��̚��u8�:�ψ���M=���#f	v����/]�j������֛n�����Ȟ]����8qb�����[o�lq�زyΜ9=}]�l~��K��'��z����%��؏~��r��v/�ө���{�4M���B�ޢ�R�lZz�L��o����7�%��9�������bŖ9
�I:jVR���&gc����.���w����׿~��m��rnuu��=��W�X���ݽ`���o����ݳ�S�z��i���`u�4%GȀ�|��8�����}���O'r���;vH�t�]_�j��J>{͆+3��eWR5�\��	Һq�����;;�����>��}���4��3S/�㴠ZFA���&��#�����=�c�b.k���Z�s
%�ֳ���+�`C2~J/V����tp!�(ʙ\�l�X�&t:��-�LEV*(@��};�R1�
�F^t�Y�P̵46QT �-G ��ʰ=��3ֽ��C9·FI_����$��r��S&�Q��N�G���
�D_QRԈ�?qA8בZ�(��!�y�gB����p��u-M���S808r���p8ZP���,F�H�ol�>��m���`2+g�O��f��i[�;	�)���0�)�)���h)��h�_�w�1���5+gu��H���v�����,��{\�N��&)��ɾճ<SӶ�zO?��9]���:�u�(%_�8|�X̿�<�Vsss0�h�O<�d��{�����^��P($��ݻwoߵ���ϱ*�-�M/]V,���'2c�U�^eI
h*eD&�ٻ<΢�<�7L>u���a��Py�a���s���}�T�Z?�?5��������o?�&��kׯY2��ӧ�o��GҐ�녛R1#kMo�:u�ț;�̞��ԼbA�P��
|GC�k����L_{��O<����ֵ�Vԧ�AY��M'#p�̽���9B˵hωCSn�b���N�l�`w.r8R>�I���ڞ���J��QqR��B�X<v�,�d*�Q�,�4MKi��iţ���F�1-�CÃ��_��аsǞ���l6֒Z2䞩���u���h�S��m��G��s6�'��ё��_���f�9I� =@¿T���`,����d�17�,�5�u���yEI��� )����+����!@����d��z~콳��k��ao6��Ro_��x�����7�s�*X��
���L������Z�+�]�O���������a:���d@>�͞=��>��7p���X��[���U+}��	εLY���$?������Ӆ�����V)z�')�}��&���JI�<!U:=�+!N�8��$9�HRm:~�mz��M��~,�	7\y%��.��{�/U%��!"~�#�͌��/����9}�U6���Q��ɼ�kd�e�;S��;ܸ���qF)rL��qi}EQ75�#��u)Q%�d
$.C��0��M�eQ�w2��NSQ��o<�7�u��Hi�֭�Q.]�-�˙|���)c����e�k�:r�G?�g�ҥ��GǶ�O�46ׅ#���r^	�&��a$4h2��֐%�-��헳N�4s'i��a�-��j�é~��T��T%O���G?q�MXl�I��cF��o��Wr�� ���ZdŜ�M��Tp��t��<VN�d���r���ᎎ����	�H�2#�T��f��nQ�����:�]�׭¡#�a��ĉ�P0 ��t������<�0<�#A`���$J�J�1���,���L#��#!6�	OD���>Y�tڤ������ԩS/m�4c�,�q��T7`�󄬽V
� �_�`ww�a���$��^M'a�c�+�V*�x4�tuxN��q&Ne��i�4渐��el���"8Z��������G9��m9v '̡]	�i����g�|<B	�t]5(�
U�=:6�E="=��Ӡ 9�f4|�U�q �N
�Q��(k�ͯw��}���~����2��H���sx��Dċ(a�n:����y������}��g�?�����'_���Ƣ!-�����/�Tש]�G����u��k�
m�ļ�@��*e��}S����W�a������ǆ�Ug�,ܦ���|b`��*�������CW	2ܨ�D�-S([��IĒ]4���^���������޶m�#�>:o���e\��+/vM�1�0G{E58sƌt�t^k��ox��'k���FG�B!�l�MA��c���(��h�;���`���c���+`+7�(o�[��qŁ�-��ƺ�N�=�w�(����5J�X�Z�i񎿆=6��a)
� ⺻O���/���������=v��e�K�$��۸����L�eTFGG��\w��3��_�n��}<��ͯlv�����Ȓ\*�\:�Ȱ�Mq]/�=#��E�`�����JX���$"�`a���E��uy�Jj�˖@�*���1IUښ#�e�|��r�L���;6fUm��Q	%e�Hk�x�� ?�&4�o�GHcTF[I0�!�pyS�^�2�.j:zyخ�x�1\�먉b�����̄`�Y����D��s�R�T*��5���U��NX,��w���1ږ���Xy��K����J�p�TW���,3��]�K&c���`��������vP�p45pU��o��J^fb�@�-�X,}�߬o��"��W�P���ǥy	�ʮo�zg���m�����{&,�@�u�4�mâ QQ�XN�9��\>�G,���*-�-؄"�~$��A:P{�.;0�^~�e��Ʉ^փ�@�T�� e��|D%��`L�U�A(�2�,�r�j6��-^2G�(�<yC�R(�q,�FQa���)�z4_q��%K.H�4������8��H�`<����Js���[F�ƍ�n������A��E]�a�q%̕a�K�,|E�JV���)y%�۝�I�^�G�]$��IP�]��]a��[a�-պ��mOp=�b������g%Q��D4���S���`���mji���m\�tn<��x �j��i--M�!�40��M{!�����E;��x�Q-�]t�2^PYZӿG�lҮ�w�>�?���(��ܱ�'Gr��y9h�f"U�8��^L����2�*�}v��CO���B5�4B�s6��O���~�������ukׂ���>Q__
+�������멧��!D���O��7��=��O����p8�OaE
��dì��&`8��,�N~x��cZrh�0MP���j6p�0���F��T*�w_Oss+��=I�E2��K����3���X�)a����ؑ�Z8���[��!���h��J��5�=�)Mp���	+G�t]x"p��9JXJq!<ڹ@�z����-���ѩ��� /�>"� Ie�|Rc�9�l��S�\�}��5ʞr�^���1iW�a�V/&H^8�����{��1a覍&��b��(��[F�|1�s�����HLX��e��@D?? �=NW���Bć��Ai�JF��KA]PtP��!���Ѳr���F3h�;'���"ɔeFN;Z1�j(
DB�ϫ .h�T;�f+��/e�=hXN8TW,>��?p��sRu�ǻ�������
j��͕"��Ķ��Z�h��͡��(k$���u�M	Y7�;B[ygᎲYi6��Z��"��S� �i���¡�J��m�I�׍��i��n�ɏ����}�����fϪM&����o"��E����92|�\����Ob�y�q5/�������B	�f`�V�Z��W�ʹ�ҋ妠�g�po���?8�mx�U�.��XI�D,+�m��n\wA0V'F��E�h��W)z��c�Ű���
��Z�{&I蒮 �X/.�9��gvv��ʖ�. s��^=�oo"�g��Y�>�g���W��������'	���_�~��Eؗ{���GFFdI
��-]_0#��M�R%��t�H�B��K��,����=��	`VZ��da�eѡ1���{M�����9�wϮ�7^9��V�m�(�5�$	HJ�G�=V@��	���U!U�Ue�&�7i{M5e$Lg�iJ���VV��ٚpʃ��t+z	LO�$�!��=\R�WԎ*+��Y�w�%�Ƈf��Q�(������8'`��6~T#B3�66�➰=�j�)��E]�D
H��]�GA���.�G��uпe�S��m`)����<Z�ǡ�g�BD�]�.��T�4�Y�<��'�L�}�LU5^T<���S��-	h�i�b��y1_��W�݀�.S+.�66��ӄ7�qQ��eݰ�y����M�&W�L��i�e�N��`)ܓ'�/��3�D��������r�������5�~hU^'�Y�%�6-�D�'����e7	�?�|۠jҭ9�gP���p��^��8��lj�`��Gr� r̃���@�F{�-�9=0�&�7�`Tv�=t����W\tksmJ�믺b��ݽ#�Q����/�e�����LC�U�6�`�1hoL�d�T��g>����=}�a꟩��I`���I�=����&���?[����bα̠*6��j[��ͮ��^�;�緣�S��T��F��̫粊T熍ׂA,$u"��C7^�a����'����,�PW��T��s����_�ҁ����C�H"�p����w����ւDnjl�lnL� �?���w�ݻt�<W��:�bXi�s2�{OPM�ޢ��{�D|u,U�9dD�p�S�V|AU}쉞��b�H֤�͙��a�͝1������4�1�#m�<���7�36x��j����]��+k���rğIERo۱<Q�dn�e �0 ��M��AD)�k�E@5�FB|��j���~?)�+G��q(�����a�
!O��`�&��8ΰp�h9��!���b�l�`I؅��LL�U1@1(+�#�o����J�|��9E��ŏ@^o�y^�xC��]��״X�<�;�AƂrA(�hD���l���~T�;E	L�gaM��rc�&����!1�������5_�_����NS�>K� 	�����h��p0P�h<V6�l&g�F{��=ݜ��̔�#Ȝ�~�e�/����'�xj��ś�x������a�YK�u�ٽ�wW��&�s}�^.7"��JC4/�1 "��{����?P���"�6�-�3�ٰ�]㓟��O���,Y ظ����q��W��>s�7��o��7�~g(�J�*H����~������#�虫��_:.�(���(���R����2��lP��= ��W_M�j�{���T6\8��+��I_�J|�;V��;�����U3�����J�=O2K�U��ʏJ"��W��<�-QAQPϪ����5%��'RlU ;&V�eWh{�Cy��H���%�W�n	k��h����.��ea`�c" ��`YV2��*r�,j ��*ϟ�I��N���iN{+�z���cq�4*��)?�|zSqt��~�Bu�x����O�<՘J��	��a�E�GB��}���<t#��7Ln}d��/~���~o���~��X��%��t����i|�Lv\�­IN�3I���av#s ��X�g�I�φw+��
��Ȉ��?"G�Y��E�y���wmG�d�I�R�R��c�;T�����"�� a���J2H��1�6��#�R���6���a��]�H2�n���>��M���B���n�׭�Yt�� �9E�����2��%+L�fc9"�	^9�����.�Ѩ!b�8�����y��m%���,�ã���(-�_ZA�[`�����6�����3��BWn����+���5��0L�T2�ɔ���X�e�R��E�h�&܃
V�EYm��K��� b��"�9�mgm�G~}�5׾��S����N�ޱo���-��J.���b<�PN%�r��yQz'q���2��ߤc�Y4x�駟\q�����L��)r�yI�&%��8�D���+N(o�V��{���so�*\�P
����ѝ�?�i3��)1A�{J�W�D��	X�&�5�Pk�jI�6iSif���}P⪞A�x��|DZ�@�����zu0 -JM��S<Bf�;���s ��'K�����-���D��g��G�Ke+o�7թ�s6x�V��YN �%�plV|HB��gn���U�M$�G
E�g��q��2�Dg��	l��, �W0���aS�n
`U��Dɥu�.�#��Y(�=�d|@���k��^�1��8�i.Wܹmǲ���l6�ߝ��J%Kg
f[���|�k������GF{{���Ru	^���QEN��I�-�j�6K��S��Gg�n��{�T'�-�p���챣,����T����K��A�*�I�3U�ޔ� �g"'�vu����t,���Ňo�=Q�+�ax�b�(�~e����X�GTW�B�bb��� j�G�?YQ�"��� �T,�������<�)��9<	%j �#��jT4U	"s��3�c�˧��oab`�������؂iVL�\1�)04E���X��ñ��:���"*B����7�kol{c��c'����`������5�P6���a�0D
ȁ��ʒ*�JJ�c�����/L�B�J��^s��񱱺���������[o����"��IGK�"��|^�eZ(�R2�Zh���l�����q\y� �2�٢�q�-�V��%�-T\����x&{���Ν;�����wht�c�l�X9~����˟�ÀY�-�,��_��!ͣG_N�G��y�J� �aN!���q©F`ǡ8Tu<m���L���HT���\5jM��$.�΢,����/Ղ<�µ��K�*��_�N��ʼ�`4�srz.�Cj!N�u&GBJy���#C�9k!���d2��Qm����`�b�4TX;�]��e��"b8��Bj���p	��h0�A��b]�{zʎ �H"���8��'ߛ(�3��|�������n�6Ծ�_?���Z��QdZ��e@�M�Q��G�Y��+!�S���

-1��UT/�/E;	($�ˠ\y$0���:|5z�����wpg2'(�C�[� �jd�8��)N	Y._�ؚi�S7*T�1���� 3j12�sh���<}�Ox�l������Tc����A�@q�0���
U3]��z�M�y$�)��@ �}]��꭫�K$��b�(�s9Brn��1IV�0Λ,m4�8 �$*��4��W���XB'
��Q1xj�ۖͩX I]G<���L���3��N��斖>tñ��e}||����F�P��jN��`(,I<5	y&l��֯�l+rV�j�N�����t6��Z��B1�
�$���h�|�4��@�uttФ�Y���zKx��1��-�����r5EA�1��q�}�ͪ��0]�B�h�rs岋�ᕻ���Q3��� ���M�;u�m�)�Onz��H�*��K�h/���d���l�0����UAȰ�O���\B%Gy�y����BU���������K�;�y���yV��x"�ʳ�>[__��ٞn��f�v3M���ifgg���TOo!��x�**�]�؇Qc���l�כ���v����El)p����A@�B�O�f��L;��^�(��pZ'�YT�n��_����+Ko������4��j�P:���T$x��\�ǶDMe��c�?����pח�����%����,(���A��;JF.�o�����U���(���0jk
���#lrʣ�F��� 
��y�a�K�hԮɃ��T<�d��Iٴ�FjPs�pa�\ˮ҅җ��`�}��1[��ѕ �Z,d�Rي�26����P������!�3B�P��I�V*�5A��#����m$�4'{ə��ۺb�G�s��]nR������!`���O4/�Fo��O~u��2�|8"czšȉ��	Vl��ƝL��i�%g#,�ðpu������@X�J]���O646q��N'-CG�_���_Ǉ����v�k�x�i�	�P�6-��2bY�g�R)�~� xK�� �#C��#�9�D����>�M��g"#�{I��
����XOhؖN�Y���U0SF�):>뜛J��'��R�u�ŦI�pOpM�����m<,ءr>�h$�z��PO� �
�/z�@�7uP� Q�ǵ\�W3��*)���1L��"h�"���7���`��i,%H�"pa�*U�H�]1���Zb�s�b�o������hѢ�'�b��H&�������P(|�����R.�|���Wo89<t��'��?�y�������/��hm?v�P۴��Z���rșV�j=����7��m�汤�K(��,�b�<�r��`�Zw��O|Ӂg�~�F��l#�]`uO1�O���u��D���p�Lfbͥk.���.��&Ϥ�?αf���m�����z�1��{OD=���j/�=�{�h<!H
��o����ݻ�_�b��E�\�x���k�t���m����s������O��,�K~����~���Wtuw������rY�@�}�e���'���B�TW��������p��
�,/����9��84ie)�M�b�.	"Ek�D ���M����(Ȥ(�8sb�����#����8x�]���֚I&�~)05�(�7��"m%�,�(ꕊUS��x�i�"�xMMH��T����#*�urF�s�������B��Q��2�K��NP���b)�N�Ĳ������3�$<�f8�@��SG�4*Ua���E�R�tTӂ.��p�0D����Ks�rl�3gμ��y|����D4��헥�e<�kyG�ǔ�c)�� Zw�a]��񾨧�c�������.1���3���	�#����M2
�uJ+x�6lΊegF��55�az-f#��)��Y2�1��B�b�.��N�&�qMQ�l1o��ΈA8[eݳE�Ҩo��H5�+B?���LZ5�'�\�4�l��>�p3a94ݢKYYA!�[,��8Ź�|��ZIT�G��̳�)��LÑ;Z�D�\��"�y���Å_�!y���7^��=���?��ϊ���1=��nm����_e�=on�}8_�Su���t0�z@�hm��x��jviP��@Sǝ��bQ���<���V>��p�>&�_1D�6}�h=��.�>MLdk��񑑾�S��l�R+
���eT��F�=�[�Xْ�z�Q�V?������Oߴ�m���Z���[��U�o��j�5\�����n��rY&[^:��M/��]7��?���˞޼�Wv&tE��"���%+o��c�������o��K�X���/o޲�T��Z�X�����zR��d˓�G�8��r�%��z	���Pjc����3]R]<d��Eg#D�>��δŋ{w<Y43�c����l%��Bޅ"�d���X&��������6xg||BE�	u1K6����N���?�)��=�*�G�/]I��}���ٴ�cGO�3%X�4�4�"\�{�<�{��*��^��E�����%'Щ�w��I�,�Ȼ�X�g�]4����Y��A`Me�ܹ`�64�:t���@}��zm��W˴�B�D�~0�~H@�'����O��E]�3��ci�3�����+��`�0ٰ�O��4-��iZT���-[-��#�iQ�ڸ���
S��_t޳[��"	���v�>g��D":T\�.��r$�:����^����5-o�j��^�3��a	*t)8�2j.�CgHp�%�C�6iVd�S���W���"_�������JP�9kܦ�G��j��`���#I�i�M͍I��`��J �/Y}q�#y}����5�5v����L������Ӧ�	�����$V#[g��<���(�[*��!���&��x+�[��`����P2�ho����[���:$����R��?�˺
��c���lI�i�#����{��1&���wO�+I�]a֜����ށ��3/�pcc��h*u�1{�:c���<�<襁	�q��/�խ_����f��"��^�l�Ek��	�!3ϋ؂����uV_}��;n�B(��8dǞǺz��;N���"h�����+
BPU%ζ4Y�J*c���/��ᡑ�3ς�RR&��`&�xh�X�T>0ҝ+s�d
%P}B4��u"k�~��[زHyOX�Uu_��Ү0D̾����8����Y��LB�c���$�x;�G�Y�Z;�&�@�����1y�D��8x��$ɠ*���C���X�����9ZP�DI�
]��k�*��h�8z)H�#J�Ӧoܸq�+[�o����3lf�9���dSSS2��7)�5� Z'A�\9_�_��+hS6Go�%�iE(�R�@"S��mW��@��m��J�G$ѳ��>���Ys:g�21%g�%J5��s��٫n}�w�r4������1���jQ���J*"|ͲQ48׊+��:D�ky���QpΔn.Z��	�j�75�"��؈��΀Ƞ�������h�,2��!rc��i�"a�!؉ N!>���.�}��}CÃ��aē鶶�dM��odxlt`hd��W��o�ٛ�l�7o��i����"��W���ǎ=t���P��ԫF����{�p����?���Nz�UB����Y�X�i5�U�<�,��v����e��K.<y���;�^�l�Y�e�27L#(K��@�sl
*ɼ�^���_�f��o_��'WT\)LH��޲qy��Ŵ��GO|�;���'�,�-�m���U؃�(1-28L����x&߯�F��z�+��;g��������=Mjjȩn����D�a�ːֶV�qG���zx�E�7:2PM<��lNX�1�H2�"�-������$T�l�/$~�-&0L�5u˗/?,��H<�!�J�rr�"�gX��X?%�g�h��kU��&���1���-��nQ`~���}����9E���d�AU�����g~��52��M���݃��a��̘e:�&.�eZ��i�c���A�`L���ml|D�e�%�/�����t G�W�QOPD���1�V���kr(����.^R(����(m��I�x.�AQq��C������u9�G�iq6=�X¿��,���?Y���Z��O?˫�k�e
�UJA���*�&��޾�a^Q`�c[�<��Y�dʉd�C5� �qܑ-/�'54���M���f�$5-�N����So����]w�ɊF�ct�6S�7,Y��f�����}��S'��z���*z,JD5�.��dA��R%�1��p�1�@� ��WJ�7�����÷�@7*f*�P%Y/��P��ĉ�ǎ����6<<̇�M��6�ky�5~��~�˟��l6�n�q�Ȯ�{�/]R)�/�����ݿ{��Gk8��M��@���4E�)�l�8��������eF�SX�Ĥc��,G����iG:���w]Z���~	�����o�)�����GOn�Ճ������C]��;�o۽}[ �|��G/]�<_�66��:=R��1�����2�ŏk���<�vm}���7\.`������z˟~����E�\���K��p�S=|��{�cZ�����ǯ��
�<�����Z���ii2���io�nL֎���y_�ͶH]�������	M>}��KG��Yˏ�x+��a��aU^�ԀH��E�pv��tzy��h� {�೨��7Vpf���Ӈ�퉄��v(|��� ؑӧ��̧?K��_޼e�,L>e����QaiZp�eko�妣'�?���Ͽ��i#�"�L��؀T�q�
�_�<L�^5E�?z�S����b?7�=�`��^z�\�������_>40��o|c��� ('ǐm]d�X�ڢ���c������?�O���ӱ��0'J�Y�ҥW]�c�>�2��k��UǠ�0��`s�G�y�-�n�108��߯�
S�[�:{��\�HPS�5kDIB{�(i�*� ��#�A����$�ϻ�!��E�;k_�������@`$S5�BA�+=�'�8�E@⣧�~4���ᆆ�H8Pm`�[<��hF��/�h衐f�*}�G���L���L]M�őYD�v]�mЎM�m١��g�5��x
Ͽ�e(�_qՆD,�.i1�� �=ѥ%J�{l|�׏g��'*���ܱkgsKۺ����Jp܂QY�beSs���$U��֌���cq8Ij4�I�ҕ+���\MM��y�f͞5myb�[���_Λ�_~��7wʢx���,�H9�H�,D���g���b8��Tbj��[Vf\][��³2!B�.�!aS�8yT(NM\��G��G�R������v��/�{ｫ�^�hlI�O�>::~ӍgN��o�k���K/��H9G�������~���R8�?qbՒů����m;�����M�o�pն�w���Es:fL'�Ҍ��տ����]�����:r�)e^x��冫�,��ES2Z���d��mZ@zᙧ��̌���x�!��jD�B�R�\$�hɒc��%�b�[mƠ��NyeuG�7�j����,J�v����TP68��(����B���\��ݭK��
̖�H�a���"�pY�4m��Νu;�)|y�k�^�N`���)���~�#�p�9E��m����&���خݯu�mi��D�_"����v��a�-�x��mf�1}�Z�hO�a�7n"��>u����m�`K��5�,�M�|-�h`R���ɄwF����o�_���q�x.7����.c&�(<�}Dc����h4
{���:6i�O@;����a'��=Ƅ��������3=��Q��L����n���h@�;�P�%I�	H��="�*rT�L15"������)ƃb�uLư4%�L��\�ԍ�111
Յ4ͱܦ��6��r�>7��Q��(O�_(Vm������x&����{��h�ʫ.[+K�׶�D�TDy�׿��H�\0wx�x�s;_��M/�z�̎��|X�"���O=V�N�/=ݕ�S�'N�ػwhh��p$fX���x�Te)OΜ?Z]������G�1���&�)����(���H�X MYv��tܱ@�ج:y������D鬼��Zy�}K��z�I�t6'�����v����t|��%�r�@�E�X��-��Dj��6NRkR��P���M��������/�w�N�N�� �c��x�´�����n�3�$�ĸ���MϿ��T�`"]����΋G��6�����k��J����Ĝ�ƈH�$"����}�w�G��Y�t��]�B�"����ɠ���u�Uk[`�K$"yѠ�x�L�1P�<�s��|ES�!���ѱ�cM7&�s�;�$��2��L��X�����w�T�ea�*�����]]�^ٲ��s��ŋ[ZZ
�h��ژ<J�M[@�*�򩞞}o�5wN}]M}]]��7Է�bqQhc����"|_ȱv��Y��i`��˅�[^H�`�ɒZ*�������|8,#��>��Mo��X�C�/䯉'b�b�T �ѕ$��\�cY�K/��)!%��"a�e�2S���^�""�=��4�H8�ɨ���!v�\����D�`��`��.�i��"�߃�fȣ%AL,V�	i�Ǽ,t=Y�����!7�����5aF$�!��</DD�7�b��MDc��x˂�\ �슁n p�b���R���y�Qv��Jmlt4V1���U RE��|XX�
)�󙉉�o�]Şz�ɯ|�o������;0���������W���Gl{k}cC���(-�3db�3�Ѳ��?��(J�h�4�bU~0BpTCh\�uX,�O����x����ȡc��ž���X�l�Q*�v��?�я�ۛ���y��7-Z0WU��DV���#��P#����]Xm����s�۳�Ã{�7B8�>��PG�k�d	3U�Lh?|^V��m��у{߄G��O�Y�Ti���_!��>7���o��gV<�8��I�6^���5�͓T=Y�h���Zx�`]e�|N������e��:3��7cN���\��.X8�������{�M�ޱhִd*�NDt�2t]�������ϛ��er��mi���X����DD���!K���Rq�	�(�Rg{���m��L�%�x��-�9�j=R#S��WX�w�HR��DG�1�A���������'>�Ț�/	�B�lN�9~���
��p;��{w���8ƖW���d'8^�$��Y?�h��8����Xc�]�s/xZcG�Q�����أ�=zh|t$�pv����ol.J��_�{z����o5���ۻo"f%-N#�B�Ų,���6G5���^r\��&�&��kO�&}�����qr�����g�L�;;���*H�H`LG`��_�bǱ;���B�u�$�'n`;����	!���Z�v��^�������yfV+�������}�X�߲;;s��������T�8.���;�f9N"�47��aZ`�d�1v}�!ٜ��&��|����2Y�XQoh�5�~�@8������p��+"LZ�c5!����$�k�d����_��g�9��ͷ�z�Gd���n�����u��mڴ)�ݫ(����w^x�W8ǰh9�n�oS�J�O$�lI���%ݒ/�ڪ1=3t2��8O*�AQsd8f(�L����P5�ds��0+V��Y�?2<�����C{q�a͊U�x�2��m�X�lzn�豑w\�剻^J*�UuF-�e�=�J�g��LF.��HX�y"l�����ko;6�|�/�������%�׾�S������j����G�����w���������Ю�_Ϟ��i��,�Om�fv�:��®��l�����XG���a�����ރ/��:�+��݀��u"
��kM��_QN�8����s�ڥUW���+�����]-d����<2�ٽ�����1���=���=���TZ5�@~�35�"��e[��ǘ	�Ҽ���4�Kےp�V�"B��T�"0ހV���2$[�6
N���J2�q�OG���F$����"GH�C#X':3`�I]mÁ@����F�Bb�2*<1^t��	�ډ��A/�7�WSM�C=�
'�H����С ��m�4�l~l�����--���ш��f�IP5sշO���{PL��8�������@�v߽��K�MGM.����Qu��'6�4-����^�4*e6��/�>�Mq� �����T�3�ʎ���c�cc�gՊe7�u�o~n�\"	�y������~�鵫�X�I(��Q�3f6XY��g�~�p8D,[n��Y��jd��qh�x2�b����Pp;<��CV�:���:���O۰�FO�o,����BV�UM�������Hpnn��:Y��ɺn��c����l�]�s2��w2/g	�h������	��}�\vy�`ᑌO�>��S�l��W�2J���i�-�5�F) �%�Q5�P'�~'5%X�.���(�*��ƚDg8�?ztdt4
2�>>�������j�9r���z(�����23۟{���a�����5��+��(������rioL�Np-b���������B>��x������PE�%K�7�k��#ǎ}�[�L'���Oy��ʚ���35>1>1s�s�_��_�#glb`lvb����x�:�18W����w��hu#��=M�H`Ǒ�F֡ܿ	|��g�TF����{VM��d��1^IT���ڄ+�G�����R�@���#�ۛ���sXdqe��D߆Z0eFG>���AF�E; �-�i�#8��8w �%�\l�n<���Å���I#��/r�7���=N;·t8��� �qGy X��]��7`�������h$	�7���� ͩJ���\�r��D.O��Ε���a1�a�;W��RN���J����CGןe�!�a4F�՜]�nkI��rR��ug�����Ke�2<2��f}��xI��t,��o��*^_��$AΆ�p,G/�� ���sa2�D��hӌ�\���� ) 
P�G ��r-*l�*M�ޔUӅ�G���4�S)ȟ����e��WkE'*:|��7a-l2b��&\u�=҃�)[L�Sr�9��S������ly֡�/��#'3���5B�RѴ���mw��Pђ�����_v�f^��(�M�JU��-V5tN��A��2{��$����vO釳��2\XS�9NB�r)W-檥��W#a�����O=٥W��~Œ��o~�V�Z�������}�xر���I�0G���8����R�z����G��68�}G�@�@$��ŉ"��b�Q�p*�D��̃�0uU���N��H]�#m>w��7ް{�.��Yc6[R~�n{_z�3V�rC�@$$E����c��]�׽2p�ҍ�"��^��P��M+���GH*������9�� �.�z�)���ڐ�̹����1�O)��8��j���6��bWlrX�'��u=��\�a k�Y�kps��ʾ6;;K�HA!�$�S�7��"�]p`�s�Œ#I"h1A�)��?��?������ӎ��=8Jf�_4Ǩ�Dq	��h!q�nK5�bB�8���B�����cZ��*D^���U�ŬV�t�5�#]�#ui-8�af
e^VV�� I� s���k����Գbuk����y||��'�M�T2���}+�hN���J7
�n(��ed�/&�`��r7�0=;�BQ���� ^�>WN.�!Y����(�kr�Փ�1*��5v��Q�Y&�܌ԫ��R{AH��|.�����d�븶��5]�S�U!��*ѳ�L���%�(�k�/9�Ik��>_#n���$O��[Qk�Z.5�<S�����,�6U D,s
�#��g�~����̞���J��l�'S{��Z�$��\.��j��k��BÇ����3�Py���QGH���n��uJY��F�����СG�olb����U��y��W����W��Ls����?u�{��81
!�\�T+1�,	��M:A���Kp�:ơ��K�u(�!�dI���N�q�7�J�|���Փ�U�`F�|g[[1?_��/��輣[�a�U�G��+��x"zb�ئ�7 C@�������3�ͮ>�BEV�y�����2��sJ$�-��ͳ	s&N�:�r��Ȓ �ALH!ܴ�lb�E���
E	O�Wp�,rq����3Kfٱ��	8���4!,��G�b,ĲH�H� R��9��2S��qhbhe�q�'��8�O��蒐�Jf(�����U�qbݞ��4�'_D����3���D�pH��Y�M��iG�� 1Y)\#/tȦ����Na/�T�_����B���4�e<2�FF0&�k�¢��BV�R���F�¼�3K���P�ϋ�D�ȱ�?��/J�JSSr����{���~<�J~�sn��7�	���/n���H\a�\�V3,[F)��a�����5�Z�-�;��V4Bu؝j�fYرrP���p&]�`5�d����Vd+5���/������g]�|�;7��4u�?]ч�u�+��������:{du�෫�n`9an>�n4*ֹ^�<:��͇ҭS�®�w���v���@N��PW	������k�[��"o�������_Ҟ�X�E�"���&��q;ǋD��'Y'_���BD���5��C�?����}��m�=���m�T3���s�Xt*�D�f^}�˄X�2C��X�W̢���;Y�t�����ݛ�����=�<��Lf����/>��xN.f~z���^��ӝ���k�{����~�`�!��7�dpI"�'�t<գ]�@F�E� Nz�m��+ᣥ����Y�j(4�:yuma|��pҌP�������b�Z���Vk�h[���}�Ħ.����cg�_�XYl���8*��޾}�_�E^�P4�?����\�Vcm�@�龟��9��xkj&3��Z���|��
N|�&�-�A��%A��ɲHm��y������' ��N ��p�[���*���d�2��7-G��j<�17���T*u����V��u�� +��-�7tSǘ����-��S�q���,� ��
v�1[D�v*��aE$������[��0� �(�Z v4�1�$���z���b�U��f��c��o!I�h�fa.SU�K.�Z�j�8���I���8���cA7nAU�~�������$R)�\��%ˀq���*~�E�
)�4$�~?#a}��%ڇy�h�P/>3��]q�e�۠���4���%�d|������*5c��;^�S5���D:��9Ϊ�Z�j&"$x�0�q�KW�+:��dzn>�Z����2l(0�(�
V�8I���1"?�k#*�ÜB�ڭ����p�wԷrU:���'6,��۷�[�� ���S���١��2�\:�?�Qz�Y�zmUS���ڡѱ˺ߙf��m������᧞�[�� �"{��(;D��rM�1��@�c��
����QSSbvv6
	��#	����4�\&�x�֖�Z�R,��B�p9A𢧑ם!CxP���꧞�)��W`Z�S��W�{��h4�L����>)�';��r����m���e��L'۫�3$�=E���5�jjN�B��ӓ��5�8��ڟ|�fp�F$²��]�8��X`%/i�bR.�|i����J�<���P=�[4Cb�D��~4)F%��3�����٭��wq�Lg�O�mX��|��X,LMO����]&��<��#]]]=�K��N=Ԅ���x����eA�XIcX���������/k�95���i_�dA�M��b�l!pv���cQB��;�?8S�{�t9���G���YV������`s���LZH��+)�PI]onn��;��8��狲�_�Ȍ��p63g5��l]��t�&�t��-$�fhR^�V�J�����Rw�ב�p�M,��MMM���A`�6��\��\��P��H�M�B�,�"뜖abNo�XTZ��c�z��>��y�޾e�l�6`V�L�yt�-���-�n��4�Ѩ�`�$,$��#���N=^U'>���ގ���%�q�D�=6zbpp�曯��Gеʊ�ݏ<|�Ι���	z�
���8Tf#�K_�����g*`G�ȪU�>�>��#����?��s������յ��>p�aEBS�$�&:�Hwc<����>������nH��}�o��P��}e�����2j�r2����^�p������'?��n8}�V����&��`��V��wg����,׵IE�"a2�� �̦�����d��bp������_pn,��b���������]��<�ry�y[������Y�Y6}��H��!�3"+VTu||����睳f��O��\n�s�)����ɋ�*���\�X8�#�t���U1�(�!%Dw:�Vd����B�B#
�#��������o�;6�"i��		,��I���uK`�ѬӼ-�,!G��~�P2�=��P`/�U�5��9'���rɚt����8ѓ��*�ˁ,�����ߤ[����b�XK��ltK,C8�Y~R-��2�����'���&m1:b�H��*� ,M=��? nMV���<l;ӵ����ࡎ�������@O_��W^���-W��3���7>��cL}~��%�V�l�=0^,ɦd67��+V����aY�Óյ�}�hʱ��M�U�V�Εl���+H���?�oҏu�@mPg�!��l�ei���|N��R�8v��K���#�$�'MG�X��H�ن-bF�j�j0ȔK1n�U��>	��Ts
�^�	�;�ok_x���[A�x<�h�ʭ[y�as�J�Dƶ�i)A�yS9���#���)d�D���5-,�h����\��C0�L&#�ȥ�^��'.gfFO��/��/��;[�~���rV/�cG�@�`�:�Z�#����\uvwo�/�կ~}����C��v��s��,cJ��+����o�t�����Ň��&Ijb�b���O�E�w�?��Y5��u%�e��U�`Cʒ/���8��D���>�TUr���	�VU�f���_���;������!�a����#ȅAM�E�3�S�����W|��?p���K~����C�Z��=�P:�r͵�._�[*d�x���}f����+�R�BP�q�h�m�p��m/���t�Cc.�䒻yN~]�-��'�lNm۹��Ǐ���s�Z�>��u,*E�6αᤰ͉��%�����b����K�n���08���_�G#����Ts[[�j�jM�i�L�I ��u ��_	�G�ׇ�Ɂ.�ʚs삦|c=��(�p�����%^'6!���]�76�	�3|46�ޠ�C�B�OO����<����U�+6n:7�͔˕��)He�EE㶶�\F��$�`�����9o�?dH���~��p�,����t� P!  �Pe����z�ѧ>�g����{j��-��g��|�884����\��s/7�=\GW��}j���UxSG�ڼ�/z�o��Xj������O|�zA��*Ss�b!3�-���e#�ؖ<��b��$��6�C\4Bf8���p�Y[�Ť�&8�\��Ǎ�j$H�� .�j�Iд���튤��U��M�#K����8Ҵ���q:�I�#��6\z��#|K�B9t��E��by�ME�y,
�:����?�Vⱸ*���8�����b0}Cl+���`Dʷ�B��/z��j9_�V�x�]�%-�~�&���VD�`}�_���]�Ńtj6[+�p����BČX�e���2GG'���<�2Ξ�-1��|�����L��������%lNu��ͳ�J����,��/�9.��[���ئ���޽����]w�=�Z�������X(�E�cYe�����K�u�Xc��z���1]�Y.���i$|�D�ɺZ�wiO/d(��K^�ՠ�G哈q������"@�T�%�V�;���0-��p�������;��=k��!�P���o�E"`I% �:�?GY2�����񑋯�a>c4E��/]��Ù��7h���d�c}g����>��e���)�r�I���$���b*�A��2'a��F�2{w�Y�nݹ�n���ܳ㥗w�Dk�-��B�����󛚙<:x�W���&����3k�m8ޠB�1� wY���P��]
�X�уaٔ��x�§����V�[��;�r���$�3�,���<ұ��ϋ�h�j^ѿj��V��h[���OG�	A�	��
�8�O�h������={$�����֞���Mv�*������(�lF�KpSC�h&��*UH� �Ta����+ŚҝKW}������_�O���~��n:>ڹ��K�}�f3������S_{�7n\�r/0�1&Sa|�x�m�M7��M�M0��o���u]Ue&O0_��>��GamUU�P��m��W�X	�	_�#8NбA�m(��!��qs����.[�jx籝{��}
WWn1uӖ$��E7�"q1g��-�!���%��QId�C��h����(;�H�.?��p<��v�����#_�C,�������ż��b��`�R�զH`�;�A�N��^��naE�Z�3zb}��y9��LI#=����#�c�q� ����K��N�٣I(bצ�h$��y�Y2M����R�\���k���믐����c���a9� X�VI	��1��c8Q�DA��Kj���o�M��U]�͍��=��- �6���E��qL|���GV��!"���^�^$��mLX�L]D��~G�����d��Lr�T��J�[|�@7OI�:a c/���FY5��B v��Cr8���3�h������ᮾ^�f��3;|�H*�
�PеC~�|����\���#p�S�x�矟�Q�>q� �< n���*�l_�~����h�X)�B���ڵ;�+��]�Ԫ<2���\�T�xO %1�Ɓ��9�+C���|(A�>�$Eg��y�	����@<Yc��8y���
)����I�>�a=��W����A����T���� �F�盞�����d2�z��`�Ph<0|��G�Jһ�;ڳs�Í����rp`tC4�(�No/�l���%��l~p�X�y����O}D��x|�����ɗ!5c*J�˃�{+���^���w�&޹��3Y���+�m	嚫/,f��F'sGV�y�/G����Q�F��=���3D�,-��[+�e!��K���}<#��9&&�d>�Rޑ� ^ :JI��ײ\��L��bDb��$�`HM7�G�^���e����f�:��Ff�bI4��/N��#���k%���i�b�ZQm���e��Ήt �$��Ō�q�v�o�X�sᕺ�Ü�<;b/X��t��x��&K�$Y�j�� �^�|!����0uÇ4;�+���pSY��Rs�~.����U1,��*XvC	Y�}a��݅�&�<t�

�eY]����;	R~����ŗ^���q��W�X����g_�y[�M;v��ݱdjj*�'Ƨj�jj�2�\"��S��h�m�c�������1?��]�)�4�F���Q��
�����wࢋ�����������N5XFOL5�a�9Z=��2�i�����N���4C��*�	�� `p�6�y��/~��_lI�E�oM�!�8�/�5G��>�ϒ!��?
�=K,M����ۃ��������S��?����5kV��Mz=��?��������pwo�E�S�щl����EKQ��x�0���Xٲ&8��!� �Gx�F���QM���'���I2?�Bh����(0��
�AF�b�RN�N�����K���yl�)p����i��≦B�HN��`_ V�����������N������~ �[����7��t��()�t��d�p\�>ųdɒ��֝/�n�r��ǟ`8%\�X�|;�yx����~�+��h��$N�k�8Z�d�fA���k��
˩L��ߍ�C�G����%�U\#$yB2c�Y�\@�p�ћ�[ТE���[�d'uL�^]�6�}q�$Jp�J�g�(C��@d�v&S�����P.�j��8.�L��[��#!#���j6ϸ>�<2:˸���J��R���! {�����X�_aQ����M8�С���qH�l���������7�l��U��T����#
#{�H$�l��c|61��`aY�@�R�(�NË��f��Q,����0�'�T+E�vA*`8���E�eg���K.���w���뻟}����5��|ֺ�D�7���P[�`*��VB$
��n@<`׊R(N7�>��S͡���;�"�rD�}t%�x�8�R����	��ʩ�n��bS޴N�g	C$ku1EJ���WE����RV��#�g��Bq鋞I5-xv�w�� {d#��)�ih��V-]����S'��Z�r���j�Y�ss�Q�86|d�U=�5��`�i����8~��WvZ�`��={>���|�u�dI!d��gi?��S�W��ͻr{K�б�~�@6[,U��-m��'�>vv�rۏ�g��S�����!�J77���\��`�-��#e�=Ӊ�\��X�.Pג32�Ct�0��as�\����Nˑ�q����-6����]�v�<^�Մ��1����H(�럾�-����UK�y�,[xAv~���`ooo�.�HFXe}Ͼ6Oor��)+�%B�>i��>���W\}-�k��geg��������������GnX�
%�u/�_���+�L-�6G����M7�76��E�Z��ג��o�R��\�lM��+��K�"0�_R$H��j�X�f-*I�5�Ql=$�Lʂ�y�ɩ��dHR��ܜVgO�*%:x�3�����y���C�/�8|d �;�Q���,e���>?�G��TS$N$;v��e��hRR,\¿CC�}�GO;·t��2BZΤH�Ż^75p�3{_�=9>�~��htvz
�i�������h��������t�M�o۶�T*e2xM,-�5Á�,www�j��z�͠���f����BW�X�TL�#�Id4��.t�8��Ѵ]��f���@��7!��+n�:���ŗ_xig"��[����_]*d׾��'(�7�R>6!�w��C]Kvy���W��U��?�+1L8	Z�1�������,ײ�L(&�~'�-i>v���}rz����1��L��y��eZ�x�`1�j\=��D-.%ehÐd���ʮk""��i<Db�I��2��2�;E��"T	��f�bі����p!?/�n3=ݝ�]��>~���ȱS�d�m�*�x^�l���.ym�eK���Np��:��=V�f�(U`�K&S�K��s�}��1vtQ A:84
F��dP���Z"�<>:��Ž�7���3���߿x~���~���v��L�X���GSm=���ͷ����=�ҹ��[!J����k׬U5C� ��cO>���k��i$�`�����_�߾��hnn&Y���n����ۯ����YU/��ëV���S�8@|k3g�D�G�1Ve�Lbx}�JM�/JNH�VUkC�G�������R�ooo_�v=�#�ѷ$��Z&��L�N����\|j�Pl�tX��r-���lX��˟� >��U-V�����#�w�_/2��ܟ��~2Էԓ�}n��˾T����]��2;;[�4&C�	����5G,�7�ZU�u��B�*������#��=B�D������B5��X7�=9�UDn^�=�M�R�5`C��1b� B�pϯ���X<�e��#�HD��>�O���G<�}�(����gW�XV+W��������;v�p�W����Y�zVg�sp����O;�?�x3�=\:��,J�Ra~v�%��z�7�p=����O?�����8���O(z�6nذa�سg�V�4kZ<��p�-_1\p�S��aoΊ�=�AD<Quqi��^`D$$��-P��^�����J��{䵀�bu���j�cxE�ܕ��7' ����I�Wl���7m�Z.��fi����@"��|�]q����<�5�%6W(���.+l{~�$�-_�b8f0�?th�g��7%7lX���>�1�«�
�II �M&#�^s�����.d�Fs�(�q��i�yC�5&�ؓ/B����	_�s\tc�y�����3�m�
��V;|tr�K{>�ћ������+���r�ŗ&R����s���$��%��ɇh����c��[�8p<�]~������_��d�^��=� �����D�;N���麷��x�W��,=�l�	/��
�Õ�Js"|b|��{����\�j�J��'�z��^\{�Ɵ�⎉�)_0'S-/��<�����C�/�y���!S��WoM7�>����|�� ѴV�l��̺5��C�p�Xpt"�>��K��\6�����4R<�A$Q�Fc�v��<�`U[�����7�LMH���*M���@�z�Zxg�?٩���v��G�7]{�m�S$ጥmA���מS�� �ήL��l�zC�
�\v���I�l�w�גj7N�^N�7��FY�jj�+���1`B-LQ��Hk@��I`�lNdj�!��:ڎ��P��Fɟ��d��#��}�33��a���J59����M�Tk�C_�_�T]ٌac.��j�
�977���*pl$�l��J5��WU�$�v��o����iG���S��$��{Jx�ܹ�$�hCb	�Y�����"��I+>�P�L?>1,�Z��Ϗ��� J5�p��c��tF�Щ8tͥUG�]����#p���؏?��ޮ�D�mϮ�_��J��%�:�=��L���jj�X��!Ty�N��qE�S��ɩ��~��[6�j:+r橧����l���CZ�5	�4mtl�a�ٙ�H$��������>��}�JE7���V��}{z����mS����?�H��O�S��կ�j2�D�� 0���Ps8l���d�O[�r��{oT�DWH�!��C��d�4'&&v�~�뮳-������;w^s啝��������G�t��]/�}9�����m���/��R�8������y�>�����{��z�֭W�������a$�TW���������}�UG�e�]-s�q!�(��Wd]�ھ��}m&;���vtv���֩�)�Z�	,���\t�e�Ǜ/�&���>gs,�\���/�-[s������36�	�rrn�_��]�ڊ�pvn*;[,�*�����=~|�R��eԖ���� R�_�%�
�n6%R�S38?H�� �<z�-��<�=�5�JE�&�3%�ڐ���^x���lUq�)[oo��WYş�`��$D��,�]��{�s����+��Z�X�����Ҳ�e	�ب�iH"�{,"$N��4i��+.�-�x��O��Ĵ4d]RH2��Вq�I����(d���iX�aS5��',]��@pb|43;����Rk��s�[���ۻ��7��C܉�HH���jX�_ B�\�$�x�'�f�������-+���T5¶�C�Ǚ��q���v�'�U*EV�%�4�6����޽��������p�V��	[�[tS� -�}���G��b�X����U ������)�r�2>>���K��~�뒪����x�:@ω,������}��m�.�C`&��e]M��[��|�]��Nc�����+���D_w���\$mI%,�-��^2q���B?�\.�������K���%����?37ud�={vW2�T��9_�T�*��
!��	��ٱ󅫮�*M�A|;ŧM?rx ��;/�H�C�긇�755�.�~���w6���Ԋ�)N���p��sl��-�0����E,o,�U� y��
��.mx���2���b�5���6��<���W�tݦ7�������7�"U&�{��C o��>��O�u�YǏ���s���;�Ļ::K5]����oAp���׺��c��)?ï~�ɫ���F����,�i���|y�S�FfP��@����n��[�f�V ���K��~�ֿ;ph� έ�z�{*55�/z��XS��LN�Ӻ(\x4nJ�Vjw�����B>X����-��]h���A|��.[F��ay�������)�K&�b=+��45�T�]R�6^tu��.\�>8T\�2
�����y����j�ٺ�Vs�\
Db�>�V�DI�l�Z��=�9Qp��t8���&�pTFB�q�R�M]$"�Ɠ%+\�y��^Y��%�uPm�<�L6�& ޅ#�EZE�^���i��a��%�uJs�e�j���i��L�j�m�����������C�KZ��&G����CU���1Yx�����߷��=��rć�>����x�S{�o��#|K�R�R�(fX������  @.k:$=���w������u�ZNF]1�YB5H;^��8�O�jƛXW��f��k���|>7�+�W�'�~jxx���t*�я~�����~__�9�΁���c��#��t�w��H1��y���R� Ҕxv~f�����t�P[�s� �߭ZvM��oʰ`���v���(�J��#2.5��7L�]8YK�
&�^)E���U�C����T���}�)-˝���h��.+��O>����}\�Ճ�D!AnP�HM�$D�6ϧU5��'Y�A���Ę�K �DE�%��.ͭ)Z��A�?;22�Uk�	f���9�&���M��Sqzp�5u�,"t�<5p�Ĭ]���_����_��G\��t�׿ڱ&�P���f�!�����lMD��h5&O�sOϠ��iGTnD�4<�v��ğ~��m���G��D�9d�W����+������g>��(��W>������|_tIGw׻�����/.9o�(�K��/��ay��f�_bL���䎾@�/Kw��Ͽ�W_�����V�I���Z������/~Y*� �����#���C�&f���_�3KVw������"���w��˟�	���ݴyu"����68�M���u\t�K��p���ĢQ�T9�"Gx��1�$�¾L>|��Su��Y�Rͫ��������я�K�>���GF�fJƧ���?��Ͼ���p�vC�YV y L�6�OW�ș �L[2
/UK�z��$5I 9!���l�HE�>R?��'Kh�]J�M�Ԩ�����ly�`��,�x���E�W?�#�]}���Y�Aa.чqjj�#	�pڶ��	,���L6[�(���X�v�:���M��Z�539E��H.�E���I�������:z����7)#���KYE�$2N�6u%���X^X���0���9�J�:�uWWrgH��4\���X��YT��e��ڡ�=��ʫ�����Bp���~�]�9����M�Z;Z�S���ubb�p���>���g�޿�����W��)���C���C�W-�6y��U�H�,y}�t*�ɇ��\����J�r�VUu̔� �M�ġ�$5���L���Y��Lڌrŕ����׮=cnh���Ll9dT�d
,�����I8yӱ��j���۷���v{�P����#ת50���VU�$�q��Ա��7ȩ/��z���Nv�
sc��嘵a�
Q�����$�G�W�Z\�4�\(Ou��_�X���8�裿{��>P)�lav6���3�j2��I6%5	-IWH5�,�O���+�������* �>:4D�-8���)p6+>:���8��CJ�9z���vvt�-E���s�-��_~��@ ��~��J�Z�^ARK%�� 2�QD�{��7=����}����s��b�e�]9��C��ٜw�������x����9��@*ڦD��ਮ����� ��H�
�1΃3�P���1;r��z<RoooKK��/����	��8�fT$sɌ)|��1��.���a�bGW��S��V���|���f�d���B����Lv_�]X+�$P�0Ѧ>� =6}�=�a�T���N�V�1�aحtv�JQ��H�K���p0Fk �ٓ��2'�g��G��;�V�ũ����Bh�0�`@�I]w�.*�	����F��:��R��m�y{��}P�Q�u�	��$�);�\.�*�R0��g3½0M�
�Dđ�!����rp���:�,��9�̋2���hY�w�����w�������tk�0_0>=3���[��{�<�W|��������l�ܚnjK7����
.Χ�/K��x8O(tb��	��+����fYӦ ��s:::^��d�V+�
�*�(B�{*
\��KfgfG'w/]�����ޱ$�@��ds3�C����_B^gS��d[[-)�7=���X�]�v�[����.[���[���ɧ�z�T�����g��Ts*�����7���E��K�����PH�I�*���L��8;H�H('���p���`�e˥�t�S��N��o�@
�2`g�i��w�~���^���+z�Y�|�g>���dx���c=�����Jf���1+ '�P$�+��;oa��-�'^�e�Z�������ٙ)ݴ:�@��:�lvb2}��kjj��u~z�\��=2�fUkc#Ӝ�A��Z�[��F�Y�P����r�9;^xq��σQ<cM�"����e���^�����+�;^|6ښ�����L`7����|~����a��@T}�\�e^��)6:����
8�b;��#.�Œ	H�4Xۄ#���8�
�:�����u%��q�_����y�i �z8\�����7�B�zr��x
��?\�b���P�Q�] TD���l8�:����a�D��8( H�*��7��I�%%&,h`u����X��~B���!�@��m/n6�Dy���E�x۲1|�A��T�	g�׷�q���w�
)�m��w���|9�65����r\ѵ�-�
�@;d�8��9R>dt��uXк����]����8����d��ѱ����B��\�
N���ӿ���b)�*�.3���ٙq�Q�|'��W_yy�ʕZ��֊`&k��\�8�so�Z��,H�HW,�j�T�w��aX(� y ��ȼ9��Ƞm²0��<c��o�4��=��ru�#559q�[��� ��Z�45�+�J��U	�I�y �={��r�_�{j�Z0���L����#�c��3�n�������V+�6e���ʥ.$���&�,h��|^u�=�,�Lg�F��4
b6�������o��jQ��jժ$�x�AG���X-�l���;��/}i�ƥQ�2s�[+��-C�ߨ����.�qV#�ǎ#�IP�748016>����+�⇤9��|���۬k�&���$�������BU�@�b C��:V:��뙟��M�\�����u�:�2�-���mO��~Co{�&A�D�����36�K��ၡ�V���]ほ�n�Gh��5��urn�Z��j2������6r|��p�Ñk��k�M���	
���$H<�"QA�%�G�R�� ��m�dlF"ٵ����Fo}���d���#��G�B�[��H�d���f��c�i��&8�*�W��Go�W�S�@Vڐ�!�#ȳ����	ȷ#�i�(�� b��o�L|���eͥLJ49�ig��h�t��(��UcQ����a.^��j�$���2@k'����$A�FpSE�Y:��Yýͽ s���cS�#$���?�fG�z�*�J�#���D"�jN�G�c�]Œ�(zHe��p�c'�Ŧ�NaT��8���#��bB�lI$�!��uɒTs�a��b>�JA
����إ�]\��B���/���~s�ޗC���yY���<K���{�/~�l�.��&��ߧ\p�k�W�? ��90�z��-����C��O���A��"�s���W��M05՞U|��t�3�R�!ɫ�{9��J�`���[�x!P@d+f$Ιg��
�
lJ1)z�%�8��g3�C�'�'�� ���yxgD��?S� � �~�L�v����!��[�Gp2"��Y�h}sn�%�c�^�Emi�]�a�7����/�x�������z�m�&�O�S���-��կ��+u��w<p�m��-_�]����w��:H��U�.ǵ����B�����B\491	.&xu�(I�Ө����hSS��/	����q���l��x��m�!b�*�H$>77G�-�d��^�?,; �LB�)U�c^��U�P-�DI-���nܰ���mE��0���yk�n������m����1���C�� ���|ȱ�R9S�W�\������臟��UM��,y#�)U�:��$=2�c������;�E--J�yT�B�����w��j�,'����.z�e���#�����̧?�Y�F���?���@���kw��R*�tl\�i�9�<��9[6��Z!!&�T��P�y���3�t�἞�%�cKe��Eӣ����y]�	�\D�TU����O���p+ �mq�~EnZ����fp�qX��cA,�ذ�r��c�B�hfz��o2o	ր�۪Z3L��W +q��#�rS:�9=ˆ�2�T�˵
�>&b��G�:)< "�e �d][R|� K��g\��g�`�E��Lo��#���?�`	�GQ:;���g ��MV�X���'	ȵ&��+��;ĩ�"y��E20�"�Q!�����y�]$8����@WW��۟?w�o�~���/~�R�p*�h���u�Y��#>�h�ʪjE�*0"��Q]#z��@�u��Xs���%-K��"D��@������,K���d:*��^�Վ"�lN�I���"��b�G��E`�Z?(G@߇PT�U�v��!ѫD⩮���]/��AE	X�e�Vw�N�bq8甉���p�4WO�t�!ѵ��k5��m��BmW�<$�� Ɉ�"}�{��v���t��t{WkWd]�X��֬|��n���  ��IDATB�;���߭����%��ۖ�Z>�rb�eWIDc�Ba~nf��~x�\>+IbsSʩ����|�'�A�DΔs���0'�g�s�lH�OV|�G�V�������L׉,!T%"\$_���#CI�h[������=�^.�IH)�I���������6o��V�j��<nא3�S:25�T����J�����Q�f�ʡ��CC�D��zB��Wa.Y�r����t�Z��6j��O¼��-���Y�f]<.~⓷._~f(�z�W�ڑ�����ŭ������}񋿅;��c"aߵ��:9|�on���ο�y�x�la.!��l�� �R���:�j�W��v�GN@�|u��3���R��P![�F�Ev��ˊ���&��l���S ���3��C4����m]�w�ɼ9l<,�|>[�V�4��ID�)~?O�uL�uѫ�ϾY!�P�������sQ�󂿹���q�����u�v����v��αB�G"��k�x�m����>CS��P��ѩ\*�s��y:DK�h�\Qf.�F>k�
����J5��[�z��۟y��h4R-���O������&����x��'9�Դ2D�H�IS8�w���C�)��t�V�������!�DBH�FCn��
�E�1�s���[�~���a:�k��8�J�VQ��%V�����N+��0�P�C�[ҫH^��LQb������!d`���Ҕ�>FIh7�������i8�f@�utph���H�<P�0="/655m�rk�b�W��|&�
�(#>޴�3�Z�����M+]�$z:�.��P2�	�}S���?�\èUJ�|�3�]�h8�ժ�ԇ���qMQ�A�f@�"�?<ppp�X�Tj�|.���i:������br���]7��>Fr�gg���:C�q�|>�lzi��T<v��w?|�}G�miN���/	"AXB������������2�����"��B}+Kp,Ի�yT��B�!��c#>ހ�3;;e �q�P%�\�|D�0�ְuW���ǎ�@*�)f9C5�0��2�ѣ�;1={|d��Z����1s���g���.k��,S�d8B��]�X	F�W���%��oS��L��#���>Y��-�=4��2_�-[~ѕ�^Y���Η�^����R�y�ŗr���ug��7��[8him޲y���φ�Z*���*��!67Y� .@ѿ#�-��v���?��0� �]t�E�T�_6A�̧mV�J�vbј�Y�B��B�]#!!�e��J�d�|\<��:�єJ��j�UM7�j����A�R�TK3捜*���HW�6;N;�?�@kM39ǭ7�)�L@6���NȨdIpL���RU}�ԚxR�t�!����ۆ�Z� p}]�g��T*M�lX�!��}4��z-���ut<O�P�		��(2 �Tb>����J&��pN�����$�۱I y���o!x$
O� 
�t	��^9۠P$��Цq	$�A�U�6?O�R�A}CI=)d�δ���I�a�.s�k��:��L[3�r���cO���˗�Zc�[T˓q���,'�X�_�VYA�%�Y�B<,���ucǴT2/��H|n���q	����b��af~�'�c�@fw���Sɧ�x�[�o+V$��f��X��z�Ųa��=+������ӻ���w����_�391�U<��X�e���+��+���aU�C�x����%/���/�[տ�24I��������Tb�/�LmdhlժU��>{}?����"�����,����٭��'�-1z���/|2����{4�A��X*hX(BBe�kX�n�(O�M�����q7+jI�@�����ٿ��q}<��=�x���������8�B$��LM�2���}�����5W �/X�m�&��8oq6��e{+ek��������}�4�y�����y��o|�Ž��
Wo8��U����J؆ojiy������K;~�ۻZZ�`}��r���.)�:T"��<1(Z�2���31d���T��6-u���&C:P�P���2��I��D�y�,1�H��Ȭ��s���D03�u�)WU���P�,גd��J�I=H�Ǽ�ӎ�-�P���Q��?�'��ǣh�a��g����<299+��֠Hf�ZrL\�"'�y�8�:�>��c�s��H�	�90<��D%ܒ����"�aE�*�5P,/�f��a皎V��*�#9��z%��1q"/�"�3�Lww7l���Vx��w��E'�&�"�{h	���G��[Moٓ�dq�G @?�?�{YA͝��aH ��������Ŋ�$�Ba��R���^��#G�#�c��B1�4#�0�y�s�e�Y��j� ��i3;_z���c˖.�#�\Q���X��[�j�l&���|�zzz_��.�R9xHpm�������`\���ת52��;��Ud�߯�Q;�]�&<z�w5_*��!���}w�\Wu��ez�^���e�]�L�qÅbS`:!!_��1|@��wl����.ْ,[V�J����޼��s�ٕe9�?����h4;���=��~z(�N�YU*�Ac��mo���׫�����e��`����F��/��r��e�W��_��tv�3ψ%h��:�F}��������Qt�
�45�ʲ`�殗��t�&�]�����H�R����Ʉ��	�3�2�sp�������頲��Ϟz��o��m[6o��o~])�M�S8�,F�����D�XϨ�;}�ۺ�;v����{� �15�}�P�*�
�5�5UM�YD���/�^�vI{gWkG�G?��O~�s��r[�6��K.s,n���}��W�����4�f��wƆ��[,V]�{��g.��}��5ɼ���@�2�΃#����W_���;Z���]pA{*=X0�XKo�7��o}��|��b�fT�P1�/���g����GG�M�Hg2u�`럏v�9�
maY6���*��T~��l�3y�k�/��b岉�������X4�'Il��<0^�@��h��W�/�!߱fT-*{����w��B!������K����Ո��kM�"U��g�VJ�B�T�	������s�:��i��U$�8dA>Rb�!�̠u��k�F� ��d2����*�m�5U���;�d�2�Y��`��*��H���x9I�bf���!�8B�[�d�s��e#~3n��i��OfQ��W@L�[ż4����!�f�D,� ��9����00�����D�X�c�Ӎ���!�8=��95K��!�9bz��F�G���T*��?y�����O4������������ʦg����Ү=�]~E"���.�
O�UXwѤ�D
����aY��"�@�E"�D2ძ^G��Jծ�MpC���ڧJ���{)�Q�J�9�σ �u0e��,֣��Cc�xQ���8��s����*Ȼ�J�-MԸ��k��y���8�dl�̴����w���5D���O�NLJ��Ѯ�]�-%`��S�#2_r��#$o���Ξ�~��琢^+W;Z�4E���R� x�q��bѽ��z�;](��g�r��j��c����/z������M��-�^y��w=��Cn8ʴpJ8^�&3��Ț�T}ؖJ���ʂ�$S�5�-ۼ��;����n��w��^~���}&h����s�;���[,� ���K�L���guEG#�w��P�sN���UyN-��vݮs����Ȥ�ߒeo�Y�駝�����LN�MOeJUn3�� �UՊ�46��Oœ��h
F����><�"6��������f����������~��{��¸8�.pׁ1]���LLNN���B�(���!����`o����j\GG̬���PEJ4�-�^��"<�1���!XY�<w�~ig.���4�-:�+����UW�E��͠���^��#�r��x���c`p���4�r�hX���d�#�4��)�n��m8�H��X��(m9��$�:����#n4P�~�TJ!�W:���e3���ր ,1@vy�/�)�����XfՅ���
cA�m�3�S��a���[ZZYkzD%[ڦ��!�}�׀$����1� q	�j|}*��[.�78(J����z��Ζ�]{w����^�&�c�K�XBWBGL�I�Z�R��U뜃�aF5WCB���VAak�	�/<�??]ӕ.p-%	sJ�+UJ���y�/��RE��$%��Rӿ��K��s�����:k���YV�z{ܲm��+�瞃ã�X���z��lΊ��RQGS}b�r9�i��G�����ƚ�j;w�X�hW8̗��eX�h,�v�Z�t�z�n��)�ܾ}��>�9�Nģ�޾>�0�-�E�@N9�U=vuu�Y�fa�����M�=��ũ�;%F�Q5��Z$b�_o[��u����ۇ�{�,�J�X*_�����5�"��6g�NT���v�T$ᙧI��*�^Q,̨J�t�l1RTIh���@��H8��5��%c�:��瞳� �ӟ�-	w�H�_����/�5�n�Zp��[3�.�e#D8�`�䲓ph1FD(����CK�e֫U�'��R$���A^����(	���y|M�ꮌ�8o��B� VP8>�%].���#�Ia۞q�`������}:;��,Z����|�	++scXW>c�(�g��)�9����45�����f�}����Lo'l�B1��@��l�X�M���j�9x� �]�>A��\�P�5���������}t� ���)�Y�^:��`���j���z�p]��F�RS�S%j#Pӄa����P�0(ŀA+69W���=�/S�p�.(hI�Ռ2���
���ONL: ?�٪Ukp�/���+o��Ͱ� R9���ܣ���,�ڄ�	����`|�a��r�/_90���42<63�S@GI�%��b{��M�i�Q�Z���]y��m���C�m���7ؿ����?�7o�ʕ��[:~�{����n�j�럷j��y���_����Fd�SD�b���dv���xt�$����v7�X)�E;��u�h���/��7��帡H$�nu�'����؂`cu��H����sX'��Ω��S����`�KN>�Ļ��]Gg{>
܏��^�󛚚��h��'�&h��s[w���o����?R�<�{kK�;���+W�����5�Y���o�떭S5�+Wkj�.�M4�+uߪ��lڱ��v��**/)�,+��"�Pwg��χ55����%Ӵ:2[�@��������;w�| �AU���n��Q���5���$�NZs���2�3}Y3s^n|�U���Iճ:2�[.8���ݝ���s���>�i�ء��c�YC�z��������̵�^����N>@,B�K�)���f�,�)--��:�T�X,Z�j�5�\s�y��ᡇn��J�b��`�S�	��K!l�ޮ�\t�x_�s��_��w����� �S^{��Np��Q��4��B �����[��r����sw:����������y�7�r�- �4M7j�'S��."���%��O~�3=�������?G<*߳jU��J��e˖���_�=u�"E,�����kb���G�L:�C����0��9�x��C��]���@R����������F�Y�����"��0�����(G}[���H	������$b�Gy$�L\}��m�����W�t`��U�W_~�K-T�P"����7#��YW$���9����
P�* Q�"ZH�'�|.�hᒥKc�"��<��!� ���<IT�9j��TuJ�j"�Bv���7>>|h���� �8;w�y��'D>4p��dv�q�.8�|۱��ޛ���>�^�m!H��EK�c�p�^b�Tհ�H���k�>���i����ŞV��=��'�y���O�xA�T�,�q�z�u@UÇ�'�
��*�����W\�����`��|ݗJ\�&��kE�����~����Z%��;SR"<��C(�v���j{g�/��P\��b�r��\y���a����#�L�����e�����#�g�ӧ�z&l��9��s�#Ɏ>ӵ˓.���17~�?�۶}���<K�L�Պ^���O�u��sH�;{N�ѩ�x8$ F�P�@,X��V��ڷwlb�g`��5���H�8�r��a��>�%��r��N���S7����ln�������|�i'��f�W�֯Y��r��TH<u�?�OƊ����o�fr�U�eN�ĕ�����ǧ'`g��8�(1l6�J65�7����$0�$�Gp�7mڤ�`�Y�@�ⶶf���v�x�s�Z�v�7��5���0uja��P�V��J�|4�^�z�/y��L���B�bO����W�ȯ)���zS��y�Z�X��u�|0#dF,�#��G��n��|������L\���h��F��Z�ӓ� �TY�l��s��:�Ȱ��\���j���,�9�8��G~�O��k7���D��T,��L�qT�$�导x���W[XJ>����]����h����H7����H�R�e���x���)��hn8VԈp�/_��8.(�#���=B�
��q�\���(lY&ǩ�3��fPf�p,�e����������5����{�tgO7�:I�衇��ܳk׭�EB�SA�B���邬x֭E��@�'�§�*�������#��,�E�*���k0�����j�7��gG�X������i Cc�,8y�?mî�n�D�IK��Ϯ�/�ٻߡN�z�Rw�G�ܼy�!Lw(�-��
wċ��(�_k��s>42�7_,�,���8��r����QV.?�R���ة���́dkr
R�!�i�����y�U0�d2���mY��N�%]�����Z���l��=r���o��񱱐$�������^�0w0�7�-���~��\�G�$q�m*2���HQ8��e�9��w��PD?��C�
�K�7�\N�uWrbl<m�4��)22�kP�$0�'&Ƈ���.��+ϠH�b�ί����m�K;�����;������x�>l!���M$<�u9�)£��/^F6�B����mK��2�����CÇ����E���4��<4
B�7Y7�O.?�oߞ��v�njmm���)P?����)����xݨʟ0K�#R#s��#��H�^	��^��o(B8��$!n�H�a�|�t��W ٛ���Ŕ��}{��F"!ͮ�Uw�H�hd�"ɰt`����Q(�y�?剁�gT�`Q���p��+�Nc�9�2�1�t1@%v�S".�
���#(-l� %�8 e�D<���iZn{{f���[�m�5������rK#[���=�i2�]>h�}��Y0!�������QyI��!�����Q�5g��v��d�$ �jU���G��6��]*v�����b8[��G��*�J�j5<FP^�#!F�g��yD�059	7��fBAF��p����B�:
���鸈��cڋl ,>EK$ �c	Dge܇l��	'�/X�s�vB�`���K��1����z}�/t�O9e�eمBIB
EӤJ.��N!����k���0�uw��,��j��Z�S7K99F�S�>�݆�q�a�=�H��] ����f�&�zE��-#�#$<l��F�F��D�t�얫��.R֠��
�7<�B��w��k��6�f]�Ux�pB����l�r\[��Q���-�l�n���ߵu�V�M��R����r�|��!ۡ 9��_�8��[c.�.Kϱ�{z����C�>�q�ӛ6<�+pt��q\����Q	�r}��k����Id�3�b��ѡC��7����x��^��)��0(bo8O)o�0��r*[�F0�e��c�1�����
e<�͞@)wt��xT�϶c�Q�q#P�K0O�'#���<��� ����/r�ꩍOL$	�;p�¡��U+��	��2�&M�L55Ā��=��ʎ����`��� ��
�������9 L��Z�H�Ea*��9��Y�&�|�n�Pc��Q��O�Z.V���qM�:,�s<��M��+|�!t`�r"�a�_U�'��8���]�ރ�/��E$����x3�d� �5Oғ��Α��b�\E��:ܻ�"�yc�:���Ţ|,\�e�
�G�[ϳy�L�T�����0( ��`Ɓ�� �j	G��ry���l���Օ��TrH�{2鶎.�ld=�B�V�������Ɗ��F§�$�8v,���7P�-�Uc�#=���
�B����� K��ʥ"|�iHV]�N�\e|�j��q!0&�1M�����@$R��@<Z��(��V#��NZ�+8�U��Ba�%��������"L+Z!u���5�"�:�kVl���U:��,[ w���s��q��a�h�R������Me�L98<�h�È9_��Pv��=xL���x�".��<;w���r6���R��Ȫ��1�B���O�q��wЖE:m"j1�#h���y���*�3���!��Kk[���e���Wlx�t�) 2��mR���=���&�I��bE��b�0� �Q���"�Zq<�\��A��4��p{ln����v���x!��W_�l�����K.Q%��G�ztt���{��Ȗ-[6oz�Fl	�>�*��x^ۦ!JRDI�⑜�tm�Y��M �ee8!���WU�*�f}:�b�6�0��c���g,P��ؙ�����.��9$�0�b�R����������o�Q�Z@r���'��
N�rv�ҥ/=��s�����c� ��>�R/Y���9l���) *�R)�\�ެ#�H�"�ֶ]p�Lk{[����;0�,�m��bK��(�IB�Egg�������I����������]]�c�?Z�T�bZ�f�V8~8.���Ikr��,N�����aK#�4�(�x<N�1��Ĥ֧��@��=�p�Zuj5?���9���GR=r�i����m�C�D)����mH�P(��B5��^嚹�?[����rm�ڊX��I�����u�h����v�;;.x�n`�>8S�l��"�^ڎ��[7}+u�>�`���'`^`���`�S�TI`�BPkM��Ɠ����`?�W�'� 𚩩)��󹼪��v��?7�CDU���Z�{2��ip�]N1�b,���nf
�m��ax���"����U{�s8���`�����(�a;�*49:̨Q:�#�	,Wi���3�MB�����`�G|g��4]78�����,.���W�)Q�M���ͱ5^ F�J������yi��9���Y��~;8{o8�4p
��/z���ƍ�J5�/���tvvLMNMOg���ww�K�h���߷<���e^#ۨ�e�@����WL'�I��Ɠ)p�Y�G`	�`����R��<1v_��HH���A�ޮ��?��9���}וW^�ם =�}����Yڶ�����O~��I��L&+5�Q.�Զ-0��Urx����^�DN�#Z4���Ĵ�8��ʫ���y+aݱӑ��޲Ƶ������퉉	t��Jr]KRu�yu���AY*�Ъ�9~a��-V$��s�x����F��-d�2��	Z[d��l^֣�L�Vd�b%��-x���#� M �.ܯ"k�"����|}j2�F�?�U�,�Hf�|F���#��s��g$[>E��$f�g��Ϗ �7:O��T�L�Gx0�*"���di.'+�
" اB@��{��)�������|�=	#�H�Riz�H�~�jB���M�ԿH-�3UYA�h#}� 
�\ȗsN@p4g"�b�יlaq��g"��&�+Ү�1���!x��;����1E���z��ѐ=gNq�n)���N�@�!у�`~�󱮓�69v��I��}1�s�����Gs��BFV�DJ#� l�;�D@�F�(���¡z��N���csG�����뢕*SL��M3W�5T���Յ�7KJ�M�u�g,Z�xj:�L$N<��h"���	�3�L�
:?o��*8&E̚�tl�'@G4��7��%���`��#T;�l����E��@�7�������hT0]�CEӨ�������Ɵx�ᡃA��t��oz������۟��������Z�������k����O;���,���e�h���lǱ�u���1_;���
���T�(uW,���I����J�t�xI{��K��e������ƹ#�!���7��pծ�*����rN�9�udIb������˖´��Ʊ7}�4��N@;�g#�rk[�ƪc=�FQt�>��`5��uYnձ�xR�'�����*�O+V.uܲ����E��#�n.�2�h_	�m9�H��`2c`U�,:2��9>�e��Ұ/)0��K����0�(��>1s}�i����'��$ P��ܣ1���p��[
��b��W	v$�7+�
��R�Ƃ���p�4P1S�[�V�Ч�����rs����ϻ�a�"|m��� b�/9.�⑁�fp�,#%V QYP�ﳆ�p�`
&�<�
��gf�z2��z�9��J#�֥�s�ȍ��Y�0���ُ69�������pA����t�O��Xn���T�@e ��sO-���Ue��Q�IR"����ˎ�˵ {1��=x�sc��p������ۊ$��H��U��S��l~�Pi�s8�	E�#
a��̞*�d!�t�rF�n��ֱw�^ê����64���;�~	e��F�Uǎ��'����������+/�P��Z�V��Amź.+���DQ|�����S����Wj��Y3V�_�k�����U/�� �n��vP:���)>���v/]��u��xp��������� 9����׊�֎5�V��j�\g+"���!d0EW�e��]��mp��̚���l �U䪅5���l�p}7k����902>9]�۵j6��Jz�z[<�P}	��FӣA0���0*B��l�N1]T�鶎�vMs\�R�I���e�a^Cc�U���`��d
���>�6AcE�[�R�	vCa��3ĉF���	�6�ҁL?�3+2E�5F�5X��>�QQF
b_�*)L)"��y:��ŕ%�n�Jvz2Ӗ�Si�H4�uLd1��Ü?͟�B�<�*�N(�4j�xP�K2�2�5��G'0����pdy��m�ɤÎ�Ȳ��d��`�� /^�r}C��j�j������1ExT�)�qW�H��5/��=�\d��%VeP�U#��h2<51nX��#��@.W.�Ҕ��"�^&s�0�dg0�2��b�D�r�5�fZá`	rXjA4��ڢ|.��w��̥�r����h!�o`��`�c� �Q�!�σ��.`'��C���T�#��!�X��R#�f�`�S��n�1Y��A��2�n�Ī�a�5��LN.\|������L�u&��Ñ0i"
(o��u7k�Z�%W��f]Pc��<'����ΐ����#�E�\�s$�Sd�q�-۞E�J'���pI��M��ܮ*�`��F,�w�^^��^�[1��\7�+�p�"u�oۙ���~�	���LIò�V=O��������G�\q��ub�s�	
՚YػWjM\x�e�|�Z������N���l	9ԃ��:��<��,#,	f1/��⇸-��	c�@J1�E]�ڸ7���p�N%���v+�� &�t��6�<���EVH:���ǷX�mf-_,�b��N��G���T"
�! �l��]�+��x��\[��&z�W�Z����Pخ�u����d�\3C6�<�,�l��ޘ��ͩ�l6��r,߳��ښ��X��!bI�LqU����J3�@'7z�Qյj�����[ڵRIT%�����T�)��a�0��h������c9$�����P�%n:���+���GD�2,���R�@)����=���I4k%ۊq�,�B�_"��J�J�<�P,pc;;��B4���EPhN"�*�J�lS�F9�y[6H8�H�-!�'G�q��c�����˕t{k� �ԯ��](�Ī�Q�h��@K�/��<�c�UQ��<6i�P	Y>�}^<��3����Z�)8�j���� �G���v/�G�
(-��%���L�%��ԣE�h��_�C˩�à(,2T��R�3T0��~)��yX4ذ�H
Y�:���	���Ec/p��F/�1���($�P=qXj���|}��֐��M�bW��R4M�� ^w����	���'ԑ�J�܏\����Zǥh:�驂�	ER�Tg("{X���Ǡvd�S��ׯFgg{�Zmo�XX�&!�G��f�ȼ��9&��)��	�?�+D�P"*;V_RTO�����B����Y)�b�y��P��o !|�!�sp��#��V5�t��H"!K1�D��f�3�*GC���V���t2��f��#�8��>��4r���v������
��h݄$T9��X��YC���%��[b�|�r�_�E��-$��t=麦��U���{���[K��C+(�EP���Y����ۓhoM妦c��B��ü��Hc�|tY*�$�%ݽ�p�����Q����"�l�{��O?�����_w��a�����_���$�۹o�����|�^I���X��Gސ�����+���hL��B�������J6g�:��_��Л/8�%��S��ɖ+R�X@��9aR_`�������d5Zl"MVS;�=��	ǭ�`4�)!Ma���ט�-����fF�b�bX5gYh�:�t���]DV��T�٩���x��}Y��Cጪ�����$jQ`T858ԋ�*����8��+�a[bM�� �5�wٲe�my&��NM��y�j��i�,�B�ЋG�ḶŲ>u&`�D$�wj���U�*x��1L߲J!-��Z<��K6!�Y=�� )%?^nh��eLRA��G��V�Y�q�݊-�@�|�/Mh`j��pXR���HLY62vA�zC�s�a���z��*U�<��Ѯ��ƒY,��/�N�Yq05O�$:�/��p���R2F.�"D�a��@qMi<��J���j&_�5�����p�,�Fh�!vR�b�D�|2�t���(K��VŌd1x<K�¿����+����ݻw�T����a;��H���#`�?�������=T-�9π  �䫢׽��#�������$<���J�@"�(�	NLl!Uu�w��7�j>8rr�����M	���|��A��E˒2-�uӯa��VTp�������	sQT
����]֙�!�4f��F�n��Ź���[��:d��K� ���bv�� ��	�!�6!��M��2V\����w{�-;�w����o�_����m������"P�l~�G����W\���-��q/��淿���]��7�q�+G尮]��/TK�_��W_����������{�ƧK�>�+_��m�\
�����6�"%ڿ��##� :�"�w]˷�s6��Nh�R�\�C�Ԏ���������=��s��͉�xpxX���h\���\�U�Y�]����b�&-q-8\�b:T�-yc��BE�.����8kF����h&;]c�W�u�4Ω�8��r���э9�/L�Ɋ�a�Β�K�<1��Z15]-�1>�/A*"@Q"P6���Ű>1n��@!:8b�^K�%Y
��
�µBI�G�o�Y+1��c9�H��&L�,4J��gci8LA+�}�"e�H+>�ڏ?����DN�%�	�Fd��D=6�F�4��N�C��oٺ�s�039311V(da*v� ��ի.��h����?���Xs��󖮌$U=��Br0xK�,O$�����t\��(�Ԭ�1g�{y{�ò��,��`
�gJ������ �vU�x��Q]/��$B����!��n�]]��X�C��\6��X,�L�VL��|�E�a��A4���N�fh2vk�!�.�7�v�l{kK�n��v�\��b�%M88ExT�W���лkU���Q�� �HkG�V�� :�[ʭ�U��J�~�Vsk�ȎDMEe,Q��n�r	~J�����`��=���j�GvE-�r�(����&i�Zl�z`9�E;]�!�5��ˆ@�h��l���[ܿ����k��r�����u�eg���s��{���3�.�3��v����?��?|qp�u��e���.^b����[�!s����g>��\{O�_}��?��O�U�J�5�^�xѼ���h�VO����b5��9߀��D"�v�i	�IB�QD��H��sr�bٚ����:���y���}���f[��,\������1G��80+��Q�+2����[,ZX���VS��\]�i���~�@�tÑB�Y�R�ǰF����b�w��B��cpd�	������S�72<�a���ԍGy,���(�(�'�aP�n� ���EBMT<�W1xDZ,�Z����-��Ov���(���F�� �B�Y׵]G���K�;�i�g��99{ �De�P²f
�	,��(�#b�&�Ѧ�8�GX}Vn.4Iw^��U�,q�)����v��11:>r�YZ��f��m�w��;p�3������e�'�����nZ�r��"�a���l���u}bl~Q��X4�LĊ��m� 
 ��@gVY��F���r�%�Ku��5-۵s�U5x��~�j޶&V���Kᙬ!�rg7���ɉ�q�=]�޾8�Tb�j��$����R� �0�(, ���	n�h��w����g�y�W��%�ȆQ^�`��3�jmi��e�}�ёCp��b��kE"!*���8"�"���40�xb��W����[�u�_N�h�j�4k���|�Y��]��B<�%����?�p�wn��O��2\���noo9�����T殻��ēA�}�3�2�
�mm�a�Pv8V��	�rEO+�����`	��q���n0���+�|ԣ��F�XM�/:�ן��<����؋]tђZW��<]���-�̏�x�	u��F�������%ԛD����G>��Ï��8<鶴��"3������+�.�H$�"�̭^5���7m|lc*����%"�<�r>�*��&���u�P�O�G��=j20����'R�l6w��'ܶgk����'�Ο���MFv�g�[�l�bj������h��WY}+G6�F��:53�(r8�U~o|t�w�����a�-��r��^G��+�c��5Vm̔�컘?��t�Ŷj�]�U�Q��q������|�`ϐ���
岁�l�u,[��阶�aO��y>M���㱖D"���J�}�e�#���P��wy�Ě�)8x���$������r�j�4�{"���T�H�F����E���\P�B�c����՜�΀'��;����]ʾ���ꛊg)�O;�԰�X�B��,^�������U#������=穀J���/~�ɏ~4��ص�[n��u���B5�A1���
XBЂ~ȓӦ�߿���_dǬ��_���$���lm��A�F�B�����>xp��p_w����;�o�O5w�Xp����(��/]aغ��c����%K�\�p����>���?v���~Z�p�O<�ß��=׼+�iE��Ig�3#�U	<\	B������!��&R��O'�w���x�ӂ�H�B��v����ŋ����G?��80�o�kם8<r��?��ǯ�hKKzjb�<j��/�8Rf~i��.1(͐Y#<"�4��~4���l���]�n��=�'o��_���dgG��#).��L��=������w����-O���[;RW��b`�.��~�q��T�d;/'&&�Z������g���^z�I'�ٿ�ܾ}�2�֎�.�G���X`�b����T(�5���u�Ql^�;�g2;~p��sOm�d�kr⬂�U*�����2��
¤�[[[k�191����nkkx��D�p�8�����/	�h�h[�T�����T�����L�:::	��u�<rS�G5fYgU�́B���,�Qvlkll�����L��u�6y�( 8��7Р�S.��C8::#W$�
v]��貮ˊ608X*����F6�h2T�1���a�M�Q������#�Nи�8*z�(Yu&:d��V�dFԚP5AH��&�a𬬤�#������(���M�)s�ˋ�B=��T�%-hɾ/4@`A��C�����rnh�z�ݏt�[������*��ηˆ�H��q���󞒚����;Ɔ�-_�E�F(3b�bMk,�ǔ"��zH���H�*~�{7�i�3R*#J|T�x��'*	
V�"~��n�y˽��W��[Zi���C��Lb`���N�gp$6Q!�I��ź�2���ٮ��pp.}��u�������`��ܽ���tAKK��D�V��H�V�j֭����9�A,��&�`�"u ��.d.?��
��i5X�Ӗ����W\�ޑy�Ƿ������tv�o����{��6�r�ͥb%�˥1d6J�c� ��9�=�c
��l}|���K�t!{����n�뎓�7-^�D��z�D2P{7o]��ꌱ�G�{�٧��w���.>���߻���{���� c���T,���|���㸕��^ ��B>�7���::,��d�0i�n��	n��)�� ��A���PC����a5ّJ��?�����}ۿ����B5���Ё1�D3����B�m�b�lo_�^F����w���B��D�f!�F�f-�l]�r��������'����_�5c���+"UY3�F,�jrP7"J��v�_�8�_� ��{�GH�4kc�6m~F�˗^z鼾�}��?���CC�E�4�sʩ!
!��ǽ�>�O,Y�h�c6<��ѱ�\V5$kҵ)"�������d"�s��0��5�8� S��؏ %Єb����0�N��� �@U<��} �xD�P���,��X��X����zs|���!d)�-]�^����m��~����A�S'��0ϢG��ka)�b��{6Njء�ծ�{>���S38-�����QQ���3ð::��֩��+���'?���n�d�<���XB��y�h�1����K?/T:�;���/8��Er�!�8q�/(�G�y���{lM��^�΋�.����yF�%ٸٹ=��F��5!�Xy!���\�X�46<�X�P�](������}�lzf�c8��O^?33�[q\���	"+м̠	(��<es=�?A�`E�^&�or�8bJ�U\��0jN�p,�P��� B@��l>��d�/\P��G��s��ۖL���S�"��X&�>(�cP��C�ZD�@��q]��8T�o$�Xsm�)a��)���3~��S�=���~��o���3�8c�����3n�����������y�Q�Z6�%�p�z���/��W�8�R�o}k*��u�?����OãS'�t�ǯ��S�V��cd��z�3W_u��~��`#.^23ڷ(?׵S�0�Pp�lBŉ�2��ϞO���az�K^�W)�n:�\�jI�K�RD���Trf&[���G�|8c�c�l�Z����k:Ɯ��N-���Q)gH��;��=�Z�I�nx�R͉|x��M��&�?�.Ϳ�qL՘SiO&�G�>��]��oVk7����W;��N=u��˧��� �����*�E�</�) .�N8i5��eodt?��"����Bsr�}{���(���-�l.؂،(���U$aK�9�WlS���PX�p-���LU_eN��P�\�r<=�ְ�
GIEO%jv�[�1Zܶ=*9s}*hD���!���1�eh�f ��!Y��[��Q[(��-}}}~��?�X��V�5��=S���5<>
c|d脓N��W+L�M�8�'��Ɔ�/��������+o���w���������R=���CY�J ��5%*EI��Ԥ���[���܎��؅筸�dAE��'<��Z�~����u���>�wׯ;��R��#y�T�9��>Q�9�\�5�l@ʁ�t<b~�9E�-ӎD¢(Lgs0Up�{ۭ�H8;=��Ѿ~�ɢ�EB^���������7���HH��jk:��<Ƶ8Jc{(���b����
��eA�H����s_pE�G��HP���nۮgXu���}/n�?���T��#��ի���7mzV䮎���̾��Ko-�"�eq�đ�D"!��X(B���S$]Ġ�H�
�;���@B�1������!2����#�3�Oɞs�)�.Z�n��l1�	�]v�{ٛ�b#�N�Z��?�ֳ
�e"�7���.ف�J��K׮�'Z)�u�P�~���r���yg�?���0_Ò�PX��_V�L&��຦ab'k(�,fl>��+����'�Çƿ�ůTl\���;�:i�?|��N�@��j�$I޼yS�>�����H���g�Z��C�T*19�"1/-�@U��m�&G��8�F�����+׬L'�Uc���\���D�R.&�js5��~����k^S����š�g�(\>���3�����y��@6yC��|>[�˗,�7�S>��q��;�/td Hs�P�eAt�$^�8��bAecP��r�wK��H�eE	�Z�V�5��H*���Mh!�����6͛׫HT{҈��8؃gH�.�)��t����Z��5��G0h�˗,�±�t�f���)��]qb&?�˻����bU��hhͲ��S��m�6��|/�L�t��u�m�k=�q��@�qk��<���c�&�l�gsn0�ò�ɡ<�s�HWϼS��y�@�Vs���� �[Y=3>Q�p�R/��]�]]����h��!�9�;���k� �A\���bQ�;p��6�j$F5�;�.�\���\P��"�hφ􎶋�����U/��n�V)�"/"C#/I�u#�����4$0^B�n�%����#�;	Gm2[�\����ԏFC�K��=�-�J�h�����SO?y޹�]~�^���G����}]�7�$�ex=�3J!I����!��om������P��r���ׂz�5q�����d�ȭ!���DCp,,s�?6�&��Z��r��R\�;��v@�P$_��o<�:�GQ�eU��3�p�=8 ԛ���<��I�,�J�3N����ki����y��s�XV�T�ݪ���e��.�V�8���1<<�}���C�`)kA'�rϊD]'���o�e��gS�T�`���#05U��k�>�1ExT�ykrb�Q� ����9����=n�1�`�D��wm�2x�wS��G?�tj���*�P"�!Op��n�P���t[ж��=�	��̂>����\���H��P♍O����֮蟷m۶e�V�C�H2	G$�g�1=�=phh��='���%��)��]�}��bBe�j&w䕏��=����d2��s����4̤l��<����IٳwH��u�jI��u����������z��g�4?���mͨS�/���|��ז˅r��e��$d7`��?���$!�{a���Ν�Lz��U}})��)H{KX4�N�f<�������kV�KG�z������z<�(j�,�,<A2>�^@d�*�0L��u�Ϳ~�g.Y�ܔ��.�,˼�l�`{k*HS���������]�e����*3�������2���,r�,���İ+��0��X�(*'yA*Oz�����ħ?�����LX�"�����,pmtc8��`^�Q+���t����T"�yOě�ݙA\3�����u[`-(�g1��Ř3(���xY4���L�-.h�e �C�e�9Ojڇ�3\ �N�B�B�`&(�m �1��3U�t��M�
��z&�c��@��Z��3�����p8����-Z���]��s�����v���Z�J%�T�I����-[;���h��7��N�a��r$92���1����$����_ܹ����xP������ra�Bz����x��D�8�y1D����O>�؆GFF�e���$` ���bG������l۞bW��]N�9��b%����:L6�N���U\���	CE��A���yb:u�OE�TAu�����9����9��Ȇ��WX�lY8E��#�,Z���;�Z�r��w���Ω����d����"	�ͬ�d�}a��ό ����������ٹg�ޕ˗>�������,�?=��dM��G@��"�T*32<q��WYugɒ����;���l�2P�V�VE���x~z���]�����`hk(��^�@�R#W,O���u�V�*RL
6t7	uЂ�r�{�����h߸�Pʏ���;n���&]�:W"{$���OQ\�y.�6�I+�,���۞x������΋k�_��uY��z+l�2���/��C�?��!x��oP!����	ɋ��}���|��g����@N	yx���%y��TǭXq�����w�ߡ��+V�Qy��ޱ9��J����BX�r����'����Y����:4�(�ڤ~G���\S�VE�*��fA��S�s�͟:�?Y�A;s��A5:�IS�}���腍9T�&�+�F��������fxk��<⁳�X�l^�^*��������я}L\]0R]=`�
\�9՚IT^؏��l�, ��v�0FFFZZZ::;�GDA3�PqҠ�v�RB�O�w�MOO�,W�Z5�X#���u<�)£M���m!�s�g\I|���Z�,�:DQP�!�nϭ��g�[")��)������xR�f���sZ����]��k�a��C���G[ ��SɃx��`�<O)F��J�,Kk[�����&�j��c�h䳟�l{g��~�3����w���;����TzӦg�?�������O;����|,]�z��,�������x13�����<6����.Z��o>�w[�m��~�yK_xa۞={B�����r��	�^0�R��b�]�ʲ�b~'�k��mr�e��	d[�����C:֒��t��({��+�fϴmY��.)��h�ݩTRUU]��o�hLLOuuv�SI�SxY��Ū���ɶT;<��tX���Å�zF1	��<����Q`��xϻ��p߁�o<���+�����<��Q�$��G��7�{�)'�ܴy����x<�{f�Pc����/>#d�'����&h��.PeJ���3���o$�|���a¯]���_����1���\�ʫ׮��B���E=�ɀo�۵��.[��K����?o^2�/pu��_g�1��EF�>���3fD�<!s����9�p�X��g��??(|�X>A.���t>y���0+���
$���d���VC$�u8����W�.x��kO=S�ٱ��o��|� �"�K����	�2�|i��駷6�������ز���c�<`6O&��Q��`Sʒ439E��B6�Mg��[Ǵ�1E�?7�t��@�"B��1ޢ�G�af��{�Dd!��/�/�
���T�֛��\���>���dhO&�)��UrH�$����
��H8j8n��*��N]���7�x#���}�B!���4t`ȶ��/��w���g���o~s�Ν��^�nuE�+EP���4F�[T�8���I�/�������(�8��-��Px����t��LeZ%	� ���z�Q$�s� �\���"s��
%�s���ؐO&Ꭺ՚,�x��(:C�5��(�����<��������S��|;hψ\��0��c�QkD��7C���Z���Y�-���K�D�EPaR������s�ZD <C�EϷa Um\UX\% :��@��ܤU��F����g�k��S���. ���~���kO[(H�a��qe߉i�9g�ʱ��ii# U��;眐-I[`y`�4�Q�4!����z�#%���\�Ԉ�)V�P�Qsc#j~'�f=�h�T2rKbO�����n�:��g��h4:4Y���{o��AM���i����7�t�pذ�P��.���"y�PU�#GP���RE�_�Ȝ��),����E�/���1E��G��A2��p&\<Z�+0[�a�,(��I<���%��]�
+��o��9��ǊP��f4L<�*j�*,�g���5�g���$ѹ�%�8]<?MMM�R-�]r�=�����GOy���w܆�����쇳�k�޷�����χ���e�i��q�	*��h�(ayς�rt��������1F�����7	i	$������t���w��"���ra�?/ �y���M;VX�R�xGk�����?��s��y�:��TI�L˗�~���눡���^����H�.�K�#cՑ��F�1��Y��wI�mӮ�2�&�!�<��<�#�ѳ0 'Q��+�Zq���W$^ޟ[i�`Q��L��3��QHKM�"I.�r��O��EpV�����Ԣ��QF41(��!�����-���G�W~2�~7E���BE�b#�J{�y��W��+Οo�eq}�BM�^��'�#�*h�x��H��0	@ v�7�1�lg���t�L0\��P*��>���<I3j6W7V��fҭ�m�D�����P8�T��]�i3nz+��|�AڠRb�u��)�B�2��<�j�����1�)����٠tUՉZ���9�aQ�ؠp�J�"��'���1�cLzT0F �D&���*H
���d��a��}�ݢB�Ft�I6V�֪�jͬ�S�aã,]v��ߺu�-_r����;︣\,\|�Ņ\��[o�$��s�=�����j���p��_F��F3S�#W�0��5%>�m��n`тt	J�V�h�0�=��6؛(6<Z2��n�]x�#:���&xv*���j���{��:�EI��+㱠±1�����	5^����/�GS�\%+X5�BU���ƈ�ҥ���\�U9���:U�|Fڈ��g�v��JLw�4��@#�;>P�k���x�f�	�?� o���@/�r���5#�F��}����f��z>��H̎�@���� �X���+Ki�2�����(���,�.������d�:���}$j��W׾!�7Mw��]�<w*���C�э;h.x�c�)�1~m]_�<��5��k-`��K�:�̠N�-�5Xu��Zu���?�5R(�ۛo?e��5�{}�f�lb�̠Tl�&S� H8R�Y7@L�T��@L9�,1�81(+Ҵa݈f����h��.�QR�e�c��FS�4����fu���Z�
�O<����,g�5T��Z�(��("(B��e�r\���/_�>����,E�dڶ
_΃�����a���� �gP-�^L���y��-�#qTQw��G�3�a>ĉh;N�D�������_>��㣓S�^v�oo>����k�w����U+��pÿLON�x��k��V�xl�����n��md��%<�9�&�ہ�-	2/���wv�� �>�RųD�Rŀŕ�8���k��@�����!8P�Z>J^��7}�Ƿ���߻�p5}ź���{��Q�k�g��l�VuK�,Y�c�wz���K	���i�!H��J%�l��i6�E�k������yϙ]��!&���w��?yY�ffg�9o{��YX�D.���3	:	�5s��/~�S=�쎷w��w]v�����)M!�C^&͠B��'��Kx��,[��r`d�M�$z�<�9�M����
"?H�t&G5��+� <��>�C�CI{g4I�Ң����J�L�Jd�v�P`�`0��6��݂CR���0�Bo��&���Esk�`���Ex�����@�G8,I�fHhsL�] U4xf0qai����$<������/;��+��<�F7���K���L&�c�����s����{%���3k׮�6m����ַ�����ѽ����O<i�X���-�\p�����իW�b�L.�9�~��b�)���/���SN��q��[~��'�r����x+ ��Yꉧ������^/��\�20�B3&}(�
y�j��i�ݱ}��?�ïe�1sU�X�YHg3�TR�g������֡��r��=j�А�wS3(e�u��5�pQݮ��)8� D|��U��EH����ZV%p���8j���l�-mp�Î΋-���zt=�+d�N�0���:Hŀ�.���͑�t:M_�h��w�9�?�W�ܸ�+���� �iԡ�1����{�dY��!�rJ ;d)�t�6@u�lX�=U���ͳ\̦�'����}�x"�PX�<���-Y�~���]g2)����[~��M�/8���r��G�S��թ<��,MLq��F4"L���#΀��Z��%�Hy�̄�JF-�2 Tn�.�����^v�pM��Nqƴș��26n߻��ѿn��Ć�p��_��3N���f,^8]�Կ?�����7wBA�������cER8���� D/-���7��� �P�e" 7���l��A���J�P��,7����I��f���!�v/*礍L.]v�1�h24s[��'�%���A�d�lI��Úv記W$N�6`���W��@G��ʛ��bْd�5nK��=��o�0����lx��sΝ��O�p�+�9�dQDo����cO�8�K��|�zJU�q�1�/�����^m�w���mn:���W���\Uۜ�г�_��5_[0k�/y϶W;���K)8"�V'��e�y��b/��:�#�HB`�Y��A�KǞ��˖.~��7<����cK�vP��V���q�����ǲ5��а_C.��}?�� k���ǰ��/����뮶L^b�nizQ yS���!L���QC�/��@���$����--S��r}ݽ�|6G�}J0�}y<eu��ю$������(���-� q�q0f!��&�w���:���@4ˉ�� ���^�.��Qm���p������p��̤{���Ñ%�,��"�w�B���.�J/Z����%9'� ���M�$3v@BOY���w�"�������U � 
$�؉OvD�H�d����2��h��:>4�s�
*��Te1��1ڱ�f8=���H�N4����$��/���c�º7t�t'Ǉ�FWK-�����C��9��7�'.��c׽X�MH�R��A��%��<�C��� D$ �HLMY^�ҭ��B)��d����s�%����e	E6Aɖ�$y@�c��$dH��Qsth��i���M����d�%b�$}K�:S2�#��w�TI}�>��)�g�Q��KW��*IH'��ҀBn���fZ[˪U��/\4��{{ֹ'�֡��;��7��B;w�3kV��W���nGYM�Hǃ��񡁖��[���??�&�<[u�M_)��؀�{���.Ls��m�P�E�|ni������P�j�R�kw�耫�_�/Pcmt颅m�:::Z] Pc���}���EJ��q��522����BG:h��nټ�VT��1���&�K��{�����6���\��1+�U5}0�-�ݒ`C��)�ê(G�MB$X6Ev����
�R�����)��	��=R��b��шP�tAMSQ
,!�&}[���4����%��B�n�JUEe�P��ڔ�C�x�V�R颮iD:�ȥ3�n���p<K�PhA���`�.��	��*���N��N�
�iVrK�)PڞlN�]>t��_}�(FA�Ԃ��N[V�bqu׾�f,޻w���f�q��X�`L��"��U�a��Р�)� �G�X�c�w}�T���R�Vh;+�4�d/I+���e�Ƒ�<&խ(}e��>�+Ҿ?�k'H֚DD ]�၂��s�'�ۊ���׶��G�w)a�r!aW��Y�#��Ԣ�W�8���CC�mM�����=�Xb�'"����g�ߚ�d�y�WO^���ϕV�@E�����ZF��vl?���YM��@�(�&���sf1�AS��k���};�;:�c�M7��+�X��������蒤/
N���.'��}L�PTVy59T���-�����v���kD�O�lhh�T9���X7��9�iȒ���S~.8 %)$����##�@�O8���8L]rD<�t����e(�%��7�G����^^��ASs��Q�X,�4%�ڶ����3IU�����L(w�[gD���#"G x1�+#�O<a�2�r(�L��`4�D�/hy�b��
�Xj�0���b�W�kA��w^�G�ﳢ�`(�)����D���6�ג�f A� P�Sל��6�%�J��Ib8�[e<-�C%?�ѧ_��xY��~�2X��&pu��\�X��&��x��a���R�9A	��@8�,	��)���ϝ�t4ן��� BL��#��DH����l(=��ڱ���#
q{�h�1�&1X��� 7�! ��I"�Z %�	 5x*h����S%tՌ-`K��݉��;�ۦi7�����ЎRZ���S���)J�
E&m�M!M<��6��i�e�`̤xJ[}��2�WEkըT�O��i����-�*�-�59@dm��.cjӔe�,����
G��{�?����v2r��1�q���=��M71�G9��/^{����ʍ�ض{ʔ����{���m�/��͚r`_�)��jE��[	:��Q��l�D�-��p�/���s��՗]�C��*��`���uhh/|9l�n�5E�;���v�!c�L��t`����ډ��u��e a�bɽ�9��N����F;wx\^�P�E(�N��T���C����"�`�*�P$fI�*I��S�b2�2MrJ~�whx(g��	b�i���N��]]�Á��������`� $����P*as�B*��
�FFG����}]]��R)^�4��NsBw�0��=.�����C3 �P���M� �.
a'���הG��@*�}?U-��Th������n��3 ��-�����P*�c���EQ��(�v��|�2�q-Bh��Bl߃9Ķ[�٣|�)Y9�0q �YƐ-_p�Q���Y�>�P�)`Pg	2���L]��)�� �*hh*��b!�Į�Z��sJ.���xVV��,�a'���*�$I��{�����W�QA��(R�-�2x����:%�Kr�62�d�æ���1����v@z�f���bP���S�>��"RJ%��l;��B�c{�ߩ�I�Uj$�'ER�|3�q�_�.�EuJ��������5s.�b�����޹m<|��wn�قŋ6�������f����3w���W�����_��G�6���fM{�~9mR�^x����}��͘6�����QԹ���#��E}�;_�9~����n�:w�"l�u�Ɏ��y$7$G�Bǰ�<ADU����ST�}��=p��=0T�^�h�c7N��� �F<i4��T/:fAOWgy��[�k���5������#����;L�1�8 k���H44k�USR	�s_2�vuu��M\�R{��������!<�Q��xV��!r��`��Q���lSS3v����Eehႎ3�۰3��+[FFF�~|h�@i9���B{d�V��ٰ�E�BD$L���k��"p�iCӵ2VEg�M�D�WI�pG���Ȇ�[6M��J]S���l��<��KB S�	'Ŋڻ\��L���R������7z��(��B:�K�g)��h���A%�9�6���1>O�0��"�K�,�p�H��F�����d�����E��(\ �?��"T&"�Wh��7�BG�Hs	�����x�F�%y8N���Ō�,�!"�!/bKUDT��e���*bb<�x��V0rF8�yN�tV���t��uDR0܉i��) ;���L:�d(%�S�,�zQ��$�,%;ǖ�K`�R�M��+-���&�͕+��\贳OŖ#5�^rΙ5URբYA�ș����O��o�;��mk9�5�Z2w�q�E�7o�~���g�ܽ��%s;�T�⎙7�,��Ԅ��{޼y�búW�9]Ys�qA�TȚ���t.���sRo���Zd<�\m!������DjV�~n^ak��Z�zx?y��x\��p��$���r�� �'�ؓ��ө���7z{z��P�(��|��F>�:��������M7��C�����lm�o�DU���W���QC���[i�ٞ�̈́��f*�x�����V4�?�y�%������SO�#օ)7d�;����l����/~���[�ʨ��vv*�,$��j��@8"W�F�Y�2-Dq�j�C�	D6E�Y�$��$��F-�/�܉&Sr�I+^r��#��)�4�����(�ّM�\ �~ $�`�)��o��a��y:�+d���o,�B!RL�n.�e�fD����l0� � ���~�I�!i�9�!3K�C�� �"�#Fw0fR��<�L����5��z@pU.�ѻm�Vҫ��2�I�� m^5D���g`x`?�SN=QE�|��)j�x����i��5�J*G�BT�y	1I儦�pB��,Mf<�ۿ�+��/]�$�@����E`FЉ7�Yoi,~$�F`�i��	��Ӟ�E`<U��l9n+��&y͢�嫰�v{��O[�l��F��e	{�!BW\vnb�=c�`�D���B!w�X�;s6�Z<u�J�*�-�'�u>�����N8u�	�B�������� .�f4�9����VW����'V���m����X�7�/^si� �W�b1����t��u����ѱQ|e�'p �M�.��4h6!�\f"�pU����ܞ���Y4.�*�x���Ŧ�p9��d�0ڣ��.�d����㈿�������,-1v��1��=��|�Tj`�oxd��rF���E���Չ�.hhf?�,�t5�G4����5	q�=%�I��'�R�w����#�����b!�cǶ���AXF�3��h5��"��j�-H�2�7M@f�|�!z8�Ze���l��g�����,����P��0�� �j�TW;�D"]SS����HN	_����J�Sx���}���{��d8��TU�1�q��ar����98��.�1��0����8�R99���`uW�P]S�ZL���:�h�O)d�F��fZ�[N����G��������P-�U�9��Eh����?80���y<�mo�~�_���GS@\��|���d��ȱ@�=�wp��v� ZQ.�N��5ٴZ%�%��UF�kp��
�@�m�E����?�픳�|�g㯅;�JG�AɁ}��'�x��o�	�޼��oo��;VS��쪫�ʦ|�o׿���d���+=ݟ��'{ף�lx͔�>/?kv���}��K��Dk]����B6��+ަ����(�T�sf��` ,����*�Ě���w=�{��5k�a@G9��������B.S�u��3��t�e]��?��X8§�S�PV����"t�_�����U�*�a��6�I��C�ŏ2�J
���y��4IÜ�IR"j8y��ڥ��Ԝ��^*�&^�I v0R�t�����:FQq�씚��Q�|�e�B������FMu�^��Z��CӰ;��9���y��)�@�����.���i	�Y�y�k���
���ˊ,-��aA�.PrE B��p0]��"���!k34u����Q|/���+G��h���i�Ν�t�����g��o╈�"��	����X�U���Jׁ����iimN�o��E%T��q���˛0���6�
��0'bUEݿg�K.W6��Fè���<e[����"+��[<�ao��(�V���+��I�';5k��.�G��S�ppp�����gx4�r�S*�8Q��C)�H�:u��z<.$0�b��u;���V�$WQK�ͳ�����g*�Ǔ������15�W�/��u�{���W�!��#��=q�?���~/v���H��`Ss2!'Ҭ%�E����٬�i�fQr�5�O��h�TѺ�|��Ǉ�OZ{�sۧ0�BxÄ�|,YdL_|��}�@B��8��ue<��z�k�4ɒW�ּ����d�����ǎ��xV8v��=#h<>�)Ś��L���=��+�ߙj�o���M$��w�����$�K����[;洟��K/nyc���׶�ii�w���w��|��w��
����X�p_}mzٲe��oڼ{Z�Za����6�cVJ6�������jۦ��R��&g����;�؁����D�d�<{L&F
��Ҏc�k�g��tL��,MT
Kr��oKJKƔB2�֪"�0%�@�S
�Y"�{w���#"4���H���������T�����h~Ŗ�t��w�`�����K5Q�� ��*�*Q`'U�ڗ�G�����pc,����`�z�����E,�u�V_�HL�.�	3���x�m�͛7c+�M�$P��MJ\���~||��'��-����f��b!��U] ��/�(G����IU���2�R��=�Ȳ*���\�º'��k���@�R��͆$��(��CT�Lܾ��/_�%�"
��<4��,�]M��@@iG�e'D6���ۿ�z3����Ţ�c���3��w:|���.�����cD^-���~j��j��õ�������v�|Q���*:�23�j�K���#"6:*��mz��?���_���i_�����?�ڭ\��R��ۧ~��߼�����w�W�4�����O�s������=��#zhɂ%W^v�_�I����߸�P�uT|f����i��g�tcS[�]]i'_��[�>�D�#�LQ�</n�s��O�N=���S�,;vγ/����5�4ǚSN9���'���ē�-E֑�������u��/�HÔ�=b�Fw�?����w��,G88eŊ�^���J$��7O�^���?=�q,P(�S�N����i����}�>w��X�RnӜ>k��_��/��4�%�}U3!p�e����DoU��ZQ|�p�S����o౗����?�¦�7��b�%�~�k��|�!m(������o����V��3f�\r�ٻ���w�2�Q7�����ܧ>���Z��1�v�|<���
B�W��=�HTg��!E�r,GpT��c�$+X�A�����,�_B�0����:��fϬ�LOr�42�d���^���i��p�Q�7}Q�Չ�G�3E�tɛ
�f���J�u�@2��j�2����Y6�9��L&��bKr��n���<������{��Me��MՑH�ܐ=*�ϗ�d%/:�*@���lf۶m�B�.Ss"�dq��^x���AH��X_jG%�v�,S�B(Z%�27I��E�,JN(,Y@���q'Q����B��T��2|IgmK�@���B�$�JxM�f�$l6�`����1�{)v���(����x<�,�����t�?��ϧs�7��j�����_�dɹ瞋�л��3Ϻ����?��fL�
�`�u�	�V/��s�2�qfz������g��s�͌���}���hWW���!X8ص+�z6�y0�U^y�/>��y�����w߱�s��7��tq_�������SN]�Uՠד���㽱|����,������de���#���e�,Aı��j�>��S�?y��wߟ.R����ַ�q�~��g6�^7}�3ZÆ�O��t���ێXQ9y�ڧ�T�\��	��8��7�l-0�kh�qڼU+OٸqssGG�M�9+�]}�U�d*X�8�cF}m�-[b��u����}��]{/a�h�2e׮������֩A��9mm� {��7�5Ξ�²�h�f���Wx慿�@ro<�\UMuS#��Jd��1e�{UN��_���sc9�qG�paTA|�9O�������?=�����x��~��o��W(嶻^�����Z��w �(ON0&� ��J�&����ɓ��`A'-{�UT�kth�Q���+���R���rA�J�-T�_�g�ᆮ�.�K-��%1Xpd9�m�.�9"�v!�����M���[�p5��ul�O�1�3Q��6w�i��EY�4�Θ��pD���׀g�܏l.+dQ�-*�T�j�$��j���L%qt;::��eIH�J�4jI£����;K�@h}39�=��XÞ�Nɉ�,cۥ�:p�2D"�"̌�`�m�������80;a��k��HDD�t�U�.[���LP��y���2K�p�3N�L�%�`�������s,��?�Y��R0�N$�d�����`||�����q'o����m��_��������k��7nī����#����3o�a��ߔ8�, �&��7˚;;w�UBY������/��r@�?0��_<ZT\~_`ێ�L�_�Y~r��=��s�+ �����D60"7c�l�K�x-T+�re��Ԧ�v0|�ē��#�c�Ү�MKW.|8l(��aӋ#���֞u�Is�p�Ȣ7�v�u�ig�tn�Us���g��D�4��5}�)x�|`Ǚ��[������VY�9�5�L֋|�����?�������Ԏ��sXFK��� ��}�evp�	g���?��ކֆE+]����x!�"��S�[z����-/o:�Ӄ��{�yy�Ks�L��S�&b�[rg�28��L�HΙ?WVyE9�����v��m|<�K?�6:�t3�+�� Y�[w�/���NO�o012�iyg�l�	�����ݽ;��=�Ȱ
��Aj	B�$P���[�쮝��h0�r� ��M	��:QD!*d��&������)r�h���߱`�*�J�\.���n9ګ����u�JJ��EU�D!�������
装�$����q��1�3�����
.�3�L��~|�����?uÄ�>�
V��{�|�|!/rH��T�v*|G��CB^�������k��bn_H�r�P��;b�U� I!��lH+�H������r���ۇ�ĻJ&�7Շ�H��P� %��c��h6���W��g?��f��T@4T(d���MrJʈ��8j�mæׯH��V	@O� 4�C���
��-�� ��2u��lx����H�a���GS6*�٪�$�I>�C$��seCH�"C7��\ā��8��*�������J��l�`����O$z8�qU�7���܁���W���>��_�ZmM4��@6XE�f6��b2v�9���!�BN�C.ϲy�����¶��@�y`���7{Z�ϋnMz�}�w��_�̋�1�E��Ұk���Y�`Φ��]��
G��F	o!cc�S�{l�IY�Ц<q����͜���2uogl��H!��mN�y�{�zFW;���{�c9�(�@��axh��e
��3$'i��/$�!!����?�٩��q�ڕ--h�Y+G������zu�q�:|�l�ǭ��._�a����$xL>o��7�{��yK�=�4�w�� C@��\A޲�ֽ�sV�\�K&:���� c��0+y#�\"S,8��T�J-��Rٌ��v�\�?@mO��ߟzqɒS���uy;�x�	ë�����k�?6���<���w�Cr|�9TŨ��-�X.���'��V	Y�j��h�H�)R�Ĩ'��e���᯦������&
��xV�N�_��8��b3�,~B�*���ظ�p`�� 6�5�u�B!��i����H���� >L!��TGGFG��Ew��������|EM�55զ�����S���p����4]�� %��Uf"l0_�肉}ay�&�H>I��2r�P�
��0L8\}��-/��T��e%���J,�W:Oh��a*CwB�nb�<�盢�(�}��۷ۢ>��G��&a� �!<��y�4���lpA�d�.!���!�l ��$8AjSJ�����Q&X~�΄�A�+�	d��������h���A譡 ���8f������ҖW�B�:*���?�����~�Ou�Y�?�j��`d<�̺�6��r$����.܈��6n�L�8z�D���YI����N;vރw߃r�s�[���{�::Z��@�uLߵsߌ��S��y�unQ<�ؙ~d^x�1���$r��ιf����X����=^��^ߺy����u�Jݚs/j�h;9h��H$�/f�ӼK���-���+z$��[��ݻm�VM�|�/l��x��LUܾm�!�W��v�+���@�`{�A�QP��;�ք��#�x���1ڦM������� �fe�d���g��Û�er�����):ܢӓ�ˮP�/O?��������9��f���-��\*Q��wd�{��_�<��+U�1�!.�rE�M�o�~c�'���~#X嫛*�]��ֶ7~|��^��h(�����I���������C8�it:���+��u�o������Ť�p�e�hp�-��C�F�D���$8d�@�U�;6�6M�|dŰS����l�����nD}�,kLl<�}=�����	�}��u�L6%9�T:G@@�b_����9�0#�eA`���\Q�ա���@U.�F]×�{��hu�5Ѓd�xu���jk���t&��ׯz$\�&:�SI^t���{�w�~���"�s����p�,ˡpucC���n���ylln+�^�e5M:���Ȗ� �D7�8'�b4��V���ѿ�����5崊�����9X*�BNa���*���=X��0������� �Œ@�a��y��G���G^��i
��tȳ�����D�%X��KP��2����c#�_V
N�,�P��@FԘ쏁B��I}?���{'�&�j`��'SR��`�|�_���4��sx3�DT]9��Stۭ�*6�&(�g�}���y���Y�����Ͼ�l�2��Fo��͛7�\=M�\�����D�HO�a�I��o�"��M�6�Xu�����YS�"�<�Z�Q����Ӗ�q�kV�g����& �,�Ӓ�'O�_1�5���o�,���Օ[�rnQIYZ^S��h��7~��w>���?��^pڢ��j���ܾm/9�:VU49�!]�e>����������k�蓗\�\�۵�͈C��k�1���kEyod���@a-lm@顎FO؉���v3g�Ne��/Ν�r�Y�q2:��e/h���Q�q�Z<o�)��������%���b��)5ŕ�օB�yuF���|vmbd��9��uְ��T4�$�ڴ���� k�󉱦״F��6Ϣ���==3�k�V�|�e|���fM�~y�+g�x¼�3����Mj,^�E���=�m�������Eu�ղ������.񣧞[_S��9�	���"�r��jN�+AH�X�j�G;@\B�R�����oM$Rg��K.���2-}��������O--M���`(��c�.����G�я~d�<�d�d�������Z�����6�ط����K�Wt�`���O|�c�̷w�ݰ~�;jkk/���Y�f1���'߰a>�U�֬9iO����>�_߿~�������̃~���v߾}S[�.���H(���5���_���)�5%ah���}x�ғ�C��X"��G��A-b�	lx�-0L��&�X�
!m��R2�q2�	���q$�SSU��ei3��9L6�8��!��	�X2]�r�9�������q�CEӦ0���>,JLG�k�� ��4V�yL�6�2$�t�eW����)2���xg�!����-�-�������P��&ω�W�!�����ؒ�tM#�.<�*���@�!v�0{%<��׌��A���%|�#Fd��
�2 @���x�s�y�L�#V����[�����H��aeu�3��~JcX7sϽ���%����������q9=^�_%���X��!X�����ԲH�[f{!91�N6�,E6E��7\E�ě[N:�Z���q��._Z���ج�L����4���İ�@ �?���H.{��/D̹J�Ͻp���"����7�4������UA��۾J(T�[~}#�LO�D�7^}��.&�U@
N��t�N�7�d��������ɣ���E9���_i�6�&J�LV��Y�3\6{ ��+��?�qNY?sɛ��̓��מD�!_3�e��i_��,x^$����x�������\{!M.��?���
�/\tìbm�
;S��5��`�	�Jwڬ_:��c�l䜓��ɭ��,C��SV�?i�1d�<�,֥�8�a<�(�]ɷ�Y����D�H`E �ݾd2A�!��$���Au�4X���E���Ƚ+�q�7~�EW2";0<�_�z�g�ܹ�E'<����^�Gk�Ȭ��[��_�p&��"����]~����o�9p���ߡ��7�\�i��4r���A�����7hݸ�o��z�y�|���׭��m��|�ͻ��y}��g��}|U��u[���80:"#����vOh>傏�R�/�t띏��'7�݇~r���[�F�.w�p�G����/;¬?������r�ˉp�*���P����-S;$nf*�@�=��[Tem�/�M��Ok��attǝT��$�{�s^����*���#{r:"�M��{�"j�&%�H���9Bt�)����£��};Wi#��ƀ%�~\ �6}�Ȱ��w_6��y�BD�{n�C#HF�rJ�
8��{$3YtnHc,0ǳ�[�Ӱۃ�)hWi�9eRã �)L �m3X< R�^d��c��2q�%:@nA�g��|��3�A����cr�������u>r�oמ}��?v�-LC�;k����Y��u9�<���� Ɓ��gǣ�R�+�����V��)%� Y�r	�!�ԪD%�w���`I&V��Pyp�v�����!��ř�(Ǥ���5�(9�A�U��&Yw��I�� (J ��,��i��#o�6mc��p��S�SH)ĝ*vlJ?������ C�B>�ó��t�4�>��dJ����Ų�  �Q53�.�ǁmzm[��׶D�6�w��~cw���'n{{,��F2��X���T��ʶ3/� �6v��馤r\w�X�Թ��i�����+�RRE�mڡ0������-?}����rީ�������X����3��⫯��
#�q1�+����;C��y.��SfB*2Rwŗ���3������x��tA�(x⺣5����E�ڷ��s��!�jX�<nlVLMWU� ̸�q����0D�bk�|�6��󆪫ձXfh(�Iy$[���}�(2`c� t1��2�/6�G_�i�hޜH8����7L�B��>�N6�	��I}(�QC�/��XaP�GZ�fȲ��4%�ur&˛�Pb�7L����ɑ�sJrMT�A~��/���KT]�B�=� �!�EΆ��U��8����
~�<��*��f��9a�1�9^7v��=�h4�9:6��|k�4$ggM���W?
����?y�)M6=��钾�ɋ��lsSӱ��4M�\�p �M���VR��_��$q�=`� xT��`��R&�r�����(ϨE�h�X�Ϫ��l��F�#2�6�)����'e�?�3�ܢA$,����zH��f�{_���:[���LfBʑ��BZ2ꬃ�].(}i����\^Q(�j�rtc��N�t�2���Z6x���N�~��Gsjnp���q.=�nv[�Pw�W�~�ӟM��������W~����A��n05�{w�����y��ݻtm�50}�2��Uu�p���.�'���`c��$�n�P E����Nɵ���-���~���b�ԦO�B�X=��y��=���TYq��8'�Q8�8�y��X>w�1����߫CBȍ\��{Ł�]Q�k�P�&r��w@�,��\��o�d�d,�eCǷ�%8j2�)���I�@ug��z��<�����3�q-ٗL�ƒ�����z���p�b'���o(�i{Ք|�P����7�#̅*b)q�N��Á]a|����؊��8j?Ș$0P,9V�y�X�#5E�|sS�@姱AX��]r�jA�l���!���"�8 JR𗥑��Wd+�aJF�֑������\�IO�.�!�,Q/
�I]����Q�χnll�)��CH��B�P:���s�p�ᎩNNϨٺ� �Q��x�B���||h������e��KB	���%^�_����"�ict��L��Ye�Rd1t�0'G�Ծ�S�L��?c+.Q��:���}w�\y���&����w��EBm�s���|,�Ǔx�\�ac(�����UnS�23ɥ�T�&�n��C�)���k���>wm�*T�,���fn!�f�O۸�Y9���6�~Ӌ/���g�:�1���LY�|Ǜo�ڳ�O\��������8���Y�y�G.~�/���[{�e/o|������n�)@
��7��Ҳ�U����45�ٵ=��_^{�w��&��*�E۷o?��e�G��<����Vlm�ǖ!W0x���fl��&T]�W� �5�ʐR
0mp�Z��qa�V�t�[�p���� ��&G��N�$�Y�䬙���b����qX>81ϧR)���X�	�stt![�%A��p�w �`[(:�n�ED �2`6M��G���$�W)�G���\A5��+;7��/�������|~\X��h�Þk���0uE0k<�"y��,YbM�N�=�jˑ�D{�HpC�`�aG�x�ą����h�!�˸<~�Ǉ]�\6k1<���B���ߔ$)Ox���S��e���Eay�`�5!�������N�^05 ��OZ�F�j��*/;Z|����e���)=/*��PEd�R��wF�%]��t%���S����G����?dcR��N5�AT�.=�̻E�N@nX".O[z�A�oCC�E$K�h�7��|W�୷�Q�;y͚�{����?���	0SC��r�ȃh=3"� [ȉ�Y���:��;��<e�bW�u�Y�Dh���/<�D��JV_�h�_�t��'�8�Qr���O\���_����iN� �j��P�E3����bn|Z=�ߵgl���ۼ^��Sy䑖��Λ'���;W,^�m����o�Ⴖ&��;SI�Y)5��.[%�+����&-]����Zo��Y�A�ur>�s��f./���B��ӌ����5�㝦��b
<Ch^@P�ဥ`�z)�
�j�3M4�X�~q�+UV�h4�����Ϯ���&�*P�����r���$�]��p8^n��bQ�	�>EM}u6�Û��'�f�����������ՅbN)�+v�Ȓ��#ʎ��G�k�n�����\Z�~��}[����5�X�:Z���ﯪ8P�-��ƃׁ �� �.T ��)�`�����+2���B��	��`I����7cG��~��Cx��ˍ6�/p�� �/U#��5���_p V_�ȱ���vL7+P}>��tbk'9��d"��Tr�ز��u�~|ӏj"�L*�sK��Tm��P�59�����D"r�U/9�EM���!:�l�+�&�B���T���������h�՝x��I&Kb&t�LC���_�ZY(z��V�x⩧���?�{ŕk_{m�3O?�F xp���Z���R%��09�|�,��qǀܵ��G�N�/N����>4���V��Ul�5V�^Gd��֠���	xX�h6�x:�F}<j���|s�����T�~��1�M8ls�k��ĥK��-O?p�]?�^ݙǯX�$�`�	��������jj�O\x.��Q���K���q��b,�4~�r�ܬ3���UW#SA>�h)2���dq��ҔLB˥%��բS�U5DG�^��$-�[6f�h���W� J�x��pX)dYQ���nR�#��i�$i�%?��O��cw�}����x|���?�R�r|<^W[{��g����x{���}��\��[��VKn>����
��V�QCxD�r���w^���vv���6��W\�j��BA���362�]6<A�!$�c7Y��ۑy��?
���ϰ�t �@� ��@=h� �s9��iJ�{�E��x;"�����:���2�*�8<4�6Y!���3�G��מ���i��q@�:�� &Bg�x) mt����C�&ǣ��Sth����ު?��Ч��
�b>���x�s�ݬߍ1��hr�=b�U��S�;Y�p-	<!�f�����G4��KW^Y�$B�J�!�_��`��ญ��������,���8ht�Ŏ��~��_5�5~�;_޹���w���+.���r^I�X�Gb�|>Q�w474�cÐ�(�$�$n���#q��_�􇾐[͏KnW�%�S�����6��e��K���;_�>"�N9q��u�!��~���NK�~s�W�^T�b~��m����H���8<�3��O��L��ԥ'.�j``�}z�i����3�~��tZ�_�_�e���g.�DBcc#�b1��q��uG� �Ҋr>?�OW9�G?�N^p4}����n���ij��[�8y���*r�|e���=̰&��u���.���9{!��_��n��pdsY���b���8����x���\�� ��S_�#���&`�*������X44��k��|.}��QC�o8B³��7_����}x�F"l0DQL�R�u;%���t,6)I����y����F���r&�R�^�$�i���G ��p<=�e��C�|��#��B9�E%��6a�	!qy�P�1��m�m�m�V%��p��o�b�D*-:$���]>��\�.9D�s�п�u��d4Y�:X%>x��%��p�@g��nE�P��j� ƊC�{�g�|��n��7b?i��}E<��(@�5�B�(k�X�m�Z����p%�b�?<�t���"�����:Hя~/�~�
���$�^�q[�h�b,>f�~��~@��Xr����mm�/���3oljݳo/c(�gOu;Y�A]�Z+�Z�*�`��d��"6�F>�25�G��SS��CX��\.ihp�d�ڈ�33�V�44Mw��/��rMP*dQu>'s��vp���
v����@V��C��N�B~�e�t�K.��2n�.���B[s5�>gOoV�||<���fR.��0���C�b*5��j��!��#'�p)Y�+��G]D�eY�Y�I�gA`	ʩ4�M
R�Jy��V[̡W�\>�4rx'yP��Ǘ����z�Uwuwc��s����U~��={TM�|R�4>�ٍ5�M$�#�#�LFM%554�h
H�
"��}���u������QCxDc�NZf4gy�����Y�L�X�8�@u688���m��fQ5A-ے�d�y"����7�5kV醶w��4��tGB;��&?|:b���F.��-+'�� U�=6�p��Gr��*kr��ŀ[ʖ�tK86[x���	�"c���y��F�N�]�`�z_�p}m�C�t]�M������EC���w�\1W�̈_`�(dϥ26��\!�U�A�[&[ɹS��xgtE6
dL0��ƀJX�֑!Κ�����T����n����?Ies�R�F#�]v�$��S��5��֍���'JS�t2~ݗ>7�.:q��*n�K,��(z���wޥJgߴ��VIh���}�SB=�^��J�:����Ą���@`�TT� �0�"�ܵw��}�\���n���C}����ή�Ѵ�	$�r��3��[��eѤ��Ph3����:x�>Z�k��8��D}���XZ���g�x�p�`:�3�ᰦ*�=?Sc����kO˪Cpʪ�1���*�3g�SK�gN*�����qHb��� ���,gUp\�a"+���)y$|~lr!�(2�^`�.b�3&p�aK��i@�E���2��B�_1uG��˹�; �ʲ��A�u��aiGe@�)^@�oS$2�,�c���`�c;��C����[n��6���.]��[o B,N%��R8�/�吶���׷��;�ő�R4�bC:���������h�2k�)Ӟ�!G���nL%H/���F5�ž���?�H&��n��U�]x�0u�]e������w^^.
A{���,���zQW\���آ��x{�+/�q��k��n݊����E-��L��
hG���l*�N�qD�Nc��|���򏭾� �k/�؃}v钅g��-9������/��>\�<���_��'�~�؎���O������-�x�:��e�=~��6�u�}����?����裏><��|r���O�LQrY�_�t�����X�ᕩ�������J4������ _�	�N1�r�"����������pOg��={W��Z��`��6Z}�E��s��~�K��ꕼ�V,^�h��QJm=�s�K������K�,�� �J~�ߖ)�f�u�X�+!vp8�bg�!�%�Kи�iĢ�%��	-f+#]T�š�܉�^z	]�:[���BE���?���?�o�'�h� 0�A�.���E�94����^�aZv��erf����
{���6��QF�����^��.7�7ش˟�����+
7����Q���w���C��*��prm��QCxD���.{�Yީ�dWw�$�uo߈ �P�ր;�@ɫQ�2,dR�p����D΢tJ�I��P�4�K��_��6���-ӑ������ݢC2��6G�
�Q-jQ`���-��0�?���L6���'�9���n��o���ٱm��9���֛K���ǖ{��'�����:p��'؜��}IC�a/���Y�U��S�y���wЮ��/`2)>����'U��(�{�-��J�
�m��N�������}�O���Ι��m��Ϥ�m~eg2�=���?��@~~`s~�����hc.���d��%`�JzF<iu `񤴌�D����hޘA3�E�YW[�
�8~r8��HK��΃��f�y�T3u�ݷ�O�bq+�ׅ�L�'�.��4?���脵�aH/#)qۭ2�k�v�a�aL� �tD� hk��|R�cS���b�wK����˟�@!:V�X�F�p�LS�X����S6%��	��Q��UU�; CmvyΓ9)��e��w�e�ω�ˆ
����r4����,�y��'�
�� 
����Cp9eȐ@7�C��A�❠�8j?� (A�*
�Z
xL���рG���� �DHa8�vS1��^�y��������ba4�� �4q��
C��-`)�#L<�.��xr�����=�#���?��OUY��޿�ͭ��6^-�=�6!�'�|���^����9A�Pl|��3�����mkkmjoo���߲��z{��<�����K�M���{���KV�<^�pH,���4'���p3m�F��-�-����﷫,���QY+�u"�EjjjU]w{$���b�֭�3w��;����u����^�펻�9��Ys;P!OC(��o�Ў�:X�佯,�G?[�>�t(�n�;�I�#�����"d*�ZD��C�d�gxƎ���(Hה��3O�?��s�(�B���T��#�AS[떭\%:8�ӵbɴ��1����	�k�"�<��E������Ͱ�=L٘ΖEd���K�� ��^.�� #��"i�V PʲS3<'�N��W��Y׉9�6M@l�M55�<���C�w�C!�ëO7()��Q�P��(Ҙ�W�4M�󙆮�� Y� ��otr�.=���?��[�l�s,i�o�+�%HM G��ɩ<�)���P�\�i�r�zd�h5K���ٜ��l&��xYX�I�r���	��	�o�D�L�U�a��A�vۓ�#N:�)�[����>߰�7^��<�!�����50~,#@����dXhw�(b��D�R�F�������~}ޛ^4�j˲-�J�1�`Z�@
�I 	�����l�H�,-��N�6܍���-��e�������H��,�/���>|�O�G3��w�9�������V����'��Pu$��}|��E�A��W7��!UVg��u8r�'�DB�=;��5����5�ܓj�s'�H�0m����	M("op������36�Fbq)��Gh�["Ɗk�*��$��,��IL`��$���Hh�;��s~��s��?x������Y�vm�N�׷s��;��[߽`��,��T��3-)ʊ�q��Rb���e�Sre	��I8��4Ԕ��̠N��S���q/O��tM�lXEkX�@�TY`؃����V��8��6���׾��LC�8�Ah%��n���ot��u����������iij����=̛�ms>�)��/�~�/fy��� ƙ��g�Ag�g�0��>���Ҩ8���\�������ǐ+Bt$�I�l�2�R(��Kœ�P�vt4�
98]�P�UE�$8n�X��|�]�)��i���tI��8�Nl"A�|!�͆*�.�1��3�����Su��F�������ь�Jն��Ir],i�-�2��F�5M#��|�t���Ia8 b)�D��XvBU��C�E��U�"�h\�æ����}��kj���UM��x3�1�6���@��eY��8Ɖ�ٴ���&���qZ�W��ei2	�T���ё���
R��06.LkMa�(H)����1	�DȲH������sҋP'�����ښ�n��O~t��������������z�%8hU�>��h�p�0�e�b�����F�f���oM���;w΂EK�{��]۷̙޸hN�c�^���;{�t*6��*p���#sf�����Rf.��%c#O�����{����x'�S)T��:51���b�8wvǉ��/}�K��D*­gN����oh��w�{�ǯzq�ˢ$ڿ��W����\5y6o�bN%v�'�� f�x��+iQK�vt��zy0o��pD�5��bB�P�Ak�kX��5�>2���}��O���]�6>����|�J���Djˬo=|���c۷�0P�k����+���}J����>��O����i��[����|���i"wJ��n��*����)��A�<�����M�� �]Hɺ�Ld+��.jt�l�U���쉡q����DI�o��#�����4����O����5E`���|��mF�h��T1�Y:�-u�#0�V�=.!X7^���
%����c�J�A��7����mq��g�S�eO�zv�r�h�E�FRK�Ԉ�>�oL���&�z�"ASQTA`mS�����J�P�e�L.]��T����� uZ��1%�,Sl%G�q)J�a���Z�穑�˔�B� <�v�7s���J��F������h0Sr)�8��������ё���}������đ��v�,�!�@t�N[���'���	W��CK������l1���>6���2�v-���sb�ٳ��#>6����<w��-�M��R�<�,�t4`��7 ir�ɒ�j���S��x�H�L�VB�7}�֞��B�rV�5�����^r�őH��/��PU�c��T&�	Ȑ�a�&��;f̸���s;��N�2����ʢ�&�!z�p�<��� ���ħ'YHAɋbOm�u�z�����RÊ�9��E��X<�cϡ����������x@���j2�y�}yf��uw�T�k.��A����֮Y�y�E3����������<�m����e��%*6�{�y��8yMw���H��F���l{m�>*�n��Ց�����-���k.X�e��=���M7�4kN�����7�����>�ʔ���޲��5X-y�~���/u����8�S__ѥ_x�G��z��g{�z�ኋ.����Gd�wx,=����p��K�`���ל�bfP��D��~�+9o���_9��K��Zx�y���S`�Ҫ;o�j":�*�6��z�t��Q9�T?9c%m�?t��|1Q[��  _��H����M+������0T15�Nr���V�:���L&�s<Ó@�U�L��5J�c�iE�_eߗ��1t�]��~��}��Ї���ʃJ�t]�u-�Nk�!k�l��ڤp���KY�״f��*�h�����`Q.=�ܳ�"���;��Zs}}�#4)�51�nN�9��	�f�VО����E�|��?����v.�ױd~G�U�yg/��mh��yg�!p\Oo��sW��L�g�>'��1g)����� ��np��Za����:��+�HN1���}�Ʉ�m{�J����aϘ7c���K�?���.��jkG��yY=t�;��%�)��5
e���N��NV��j���x4gXA1F%wnY�}wX�%,˫�ű�,��No��!�l����ڊʑ��!�����ܺ���"���|�a�,P� ��t|����IʔG�r���k;E�I��Ѵ2�3n��E~�S���BJ�I���R��U�z8#S.�h:�LuV|�57D�}����?��v�:�����J��v4Ϊ{q�N��F�\{v���+[��v���p���
]d����O���7��|���]��]��;v�s��y�m���6̜_WGmڹ�[o���ЍW��ٶe�3/m|a�����nߴ�#��HS{��+���~�_����@K9�Ke���Xt�X(H<kuȳ4�[$�G�5Ʀ�"��ǒ0!�0��:�Q(���	����I�V�zl|��ՔvWSÚo\9&�ـe�H��4���l2uI))��xu"8�.�r���2d������IƑ�Jgʖ���9P4�S
UԞ����ǏgS�|>/J,'2,'�<`�
E�b-�R����M���>>���X,���
	�G0 ��X��3�r�������㒪t���} ��|���J6������`��1�v�a�7͘vk �~���\n=WEc�����	��!HkҺ�O�.[�R�,��t���;k��RL��4W�D�����yS�����&T�1 LL�I!�&�Hx���Y�s1��&g��yo�<�������u�ł,čY�����������m�����Ő>��+$�55�����sʂ`��6�@ld��%�p~�%��y� S%-�u�A���9�=~o6�����bʕjRVD�G7�)�s���BZL��ʱ(�AJ�K�(<{N3(�u��9oΌ�����:�=��~�+j�\���
fӔ�?�9�8k�ο<�'���ѱo�Eu����jUU�����]z��3>�\z����{�ְe��ɜ�)���	\hG,��5�L.W���B�h���#�������f�\�qcA����<���m����^{�����T<�~��_��ׇM��7�c��93_ݶ�iz��"���������t:���;w�,��Z
��x�|��YUYq�Y��H�����;����Xs����	��SE�wddᒳ�wx>t�Ͼ�aڴi%S�kFt,7!J�Ӂ�ڰك~�-�؉�b�k�8U�0eɲah�r:��4����iu<9�w�^��M�2�x,>��I�'e���I`͚��A�IQ�N͚9�}��]��$�f$�8�0���4��H6ü�w��iE��7sL+��}`n�o�ڵ����h��B!��$U+�y��L����VR�����z�HO�	2X�D��b>�]1%U	���P�G?�ٶ$�T��߹}gSC���9k��GF�*�*:��)��`0�PҘ'� v,�_��:*R�������^�O��A�:�����4���U�B���6�a78���$��'G\<dn˙B�� ��)8��jrZ(�4ͬNeCa�cv�s&_�ɡ�*�j��+�+�g��SZ�1h:�H��׌b����W���������~���_m��~�0�ӟ���v��~����457��=�����r_Y�[ٕe��?>?��F	����葞'���l
�@h�]'}��mo��T2��<W4�iij�ԧ?�y|P�����u�Ʀ���C���7�H��������ͯ�{��
��d�s��WLa�$$yUQ��H�h4��{x<�H�2s̝6�cR��éb>wŻ�;z�Ȏ�L*�lqKtx䒋.޺u��PO?��ykV���:�I<����.�du��L/&��9+�)R7}�C�<��/ݟ�e�̙�|野9TW�	n�d���8��z(]-�����W_mb�\�0�xB��=q�{�r�(YA�2�*9="X���H�$IN��W����x\��,!�{j`�jHO��9,�5�S���飫����D��b���R����<G����T]e�C���EL�>%ܳ4���c)�}�������CpR4g
�d��!M�c��iE�v�TB��0!Y.��S��2 5�!����W(��}E��4*�p�kW
Ӥw��!MM/7݅5�z��vt��t bV�;]�����V�����������
���ͻ�.��O:8�u�/b�'����\!V�5����I�G8���Ɛ���e�7�+)���p��$�g�1�t6��ԢI���zDZL���dKV�3L�U&y)���*�a`I��'��8�ocL������uRL�C��I�� �(�#�#�l���������;$������:ޥQf8���,_�iL\00۠'�#ý��ǎ�/�`���Ƿl�r�%�6nz��G^�ꪫJ��g�imn�ӱ���{��WH0YԒ!O���r
메�K��÷m��V"K`"�%8|���?2o��	S�z@����k��艮�x���`�m*�w�uk��Q]�c�w����AO/"{�}:M*�l/�<��1-�������4��4i�������s΂E�	z[[=��Z뫷nX7�����jk�]��S��77VSA�#Ͻ�5�>�e�����/^��j�Rr��zoz�v�p�Fu�ʝ�;���^۱��[/7n:�����~��M/����37�p�@����\"���1UIF�[�ۚ�\�ws-��]����](�>�9�=٨����a�\�Pa�!3VW�!N4楈:dH�5��N"�9fL��B�;v"T�e�NtH(�R,f�z��Sǃ0���Lp'qW�v�~�k����R>�N(pa�b��d���yZ�\&ď�_� ���8��i�~���u9�8qtx��z�t.���zB�M�c��H;��A��E$|�X@�AI����,pX�#C�W^�up߉3�X��_}I�S�av��?��0�e��NWU���F1D���,����$5#%c���TR�ő�i��&Չws^,-6���2�@[���a��]vS�w�.
�)��T5���'.YF�e��U��a��}_�#�l�������Q�/0��=�9�1��-=a+�)eV�/a��	D(���TC�'��&kU�H�*<kV�UW� ��_��^=��s�k��#��
[���-x�~��!q�Sk�uݢz@���2�Q���>��cu�������R�ۦ-��*�p������W���MP��J*��ƣɘ��3gϩ���N���}ss�P���}b�ڵn�WǘÔ�lK�.�����)��`4fϦR)��%��*��}>J.Q^/�|᜻��뮻�}�9����g����X��9ެ;�����휡��tb4�R�8�Y���˃�-]�����?��w?���z���g��g�����K��*e�M��t&�KD�NK���wF��.��W�ij�A99����y+���sO�����h�U(�Ot��r
8�|��ty]"&� /@п�v�Ò�41�pJ�ٌ���u�&u���l*�q��"�h]]>�F�P��TSJF��#;%* +mʤ�=45:%/�&��ā��D:��E�-1��i��Ф��0'���*��ӊ�m��!)�!y��x�m4�K(i�={�oݲ���J"UUVU���ɥ��ṗ�v�k"��c(��Ŭ�-j�H��1�
��Z0(��3�<r�8	�3C�QA�J�ҏ������x��ߺ?�̢�Ɂ`E:=��*l@U�&��`C��h &t����<��mҪ�L����)W��H��F
�0�+��ۗɪ����<���Ԁ���7���$�=%�EHs�v����~V$��nl<����r�`(����[z�4XX�8Ͳ�,bc���c���-���M&N$2 يɪ��Z0n�t��
��q`�|��P� ���=׊g�s{z{�=>7|���I.����A-�<ϪZ�|�剳?��h�-���L��t�� �l��6�L��X(�.�oǻ� �/�l�܅K~�˟�IJ3�q�� �@���c,c�h���C�Z�TE���m٭�����Woݲq�����9�ϻ���U��@�j��4&*/�ީO��R4�y�1{��e%�����S�L	U�P ��y3������ҹg.�J�G`Ƙ=�;��n��a�4����ޝK���t�:(}�#z�G�?�dKs�7��9x皫.��u��Ɨ`���*@��Ԃ�J�%��Z2��?�����͘p���L��m��WE�j��Ͽ���5�\���y��]Mӛa/^�h��~tvr����X2e)?R��W q?�uɲ�Ͳ`N�bmM����;�T��^��M������_z�E/�����`�Db�2��CN�	��g]�|-�&�5�N��ݿ�����?:�c�b)�x%������tb�D��iE��6������T,�^y�c�ի�lh��%�e����~��K&ľ�o�C3�|*3cz����ft�*��TЅ �hΤ�D2��Â�sZK�?�U�V�X1:��X����d�u&&dc)����I���R�.A�孖�� ��LcY!�pX�N��Mc"��˃1����;5�t��mm���9��ب ���&�������ݗ�� ��"ݷ]�'����1�Ӫ���`	h��pH\p��UaE&�`�"�z���圼�e�c N���oSS.B6@S����3��/P��)��}���vm��#ՕL&Ԕt"128R�7����.�~���g��[6�U��d��t�O����M{OU����p�$I ��+�J�Mb��f�SL�b��ˣ��+k�>gUkk�}����^�Z_�2��&�$���pC7�b�M���D��p��c�uOus:���[u��e��fu�ٳg��ﯯ�X�L��C�e'ܤ'�U�G,:-�P8���/(*��j`LP�X䚪�����Hs��o�de�s|\�������/�v��d��>s�M� �I�qU�<���~��x �Z����4�������T��J�TW�EmF�p���Љ�>�6��U��s��E�W�9�O�f4Դ��q�c���fj�+��,�SA�����Z�D�0�0�kX+PG�mZ��2	S�r�0�p����0]��a8VD��̥S�`.Q���O�6-K�m��'��X���ɥ3�bv���7���x&^()��L��{��^������r1�Z6��F�C��RͷN[��o�V�okL�+o֏w]m������l�= �͜�|�>U]]s�m��[�>�J����;�S�Ds{8ڂ��Ӄ`�]{�S�7���h��
�|>��^�P�z.�:��穮���{��wvuo�����U�6��m�<�䐞DԂQ��.Y�9�|�P�����t��Sۍ��[T���{b���\�X{�E��޺���,bM�� 7�ig�[76�f�'���́L�w�x�@����iPR�R6S�kE��J|��n]c=.1��s�
x����eNO�Mh��U�m�i2 �U/X���g�=���<�����.L�筎D]��������>m��+V��W�<�~���eNq�ڿ�	>�7)�xaΜ9<� ����u8��P ��9
�*9��}C���{���5矿��v��5��xH a'z}��S*�l�0֛(�%�)�[=>:j(�C��R ��r6��K/}��7l��կ��l"M�-2���Y��N�V�+�eCI�*N��NX\+��$�L�utcu8��b��pEKvM3ڟ���*+H�%�z� xUE@-ɑ �(���0�}����Yʹx��Av���!�z"�R�Z^ȱ@s0�|^l��ϥͨOf�l.�%l�%��c�w��"G�`����xJ�l���d����.Q+k��и����Ay<�/LCx����j��r:c�ؾ�{ל���6�'I�|��C׆��MF�0��~uu��'�'R�pW>�>����v�`���RU$��y�������ӊ�5�-
r4:αB $��t���C��J���b*�7�FMMM��6=|���j��d2����S�R2j���.����͞�h�Y���?��.�M&�^�;O�.��JaN�A�,z��*
ա���;;B
+m�&E��ЉU`
��u8v�w~���o������[�0����d���1i�v�Y8��������ֳI�@W)\�(������9w%����E5sǎ- t��2��$9@�0�I{����3L�Z�נ��r!����yײe�
y�}z{I�J�@M�j����z_&��[2����z������jj��l���ҧ �@�mvMk�Jֱ�l9���
�����q;@���`�744�o��Xd%	@U�w	;��={չ� ��Ҭ�g?�?�Е�*d�׃�&�z��-Sz6K���L�� ْ��u�����PMs�k[75�׍?�\k��3���g��9���n����Rj���'t�v�(�@c�<<d���O�.e�vrH<������i��)]�$�"��F�%��!�w�GF뚪\�odl���2%����� m��H���++-�u�X@S��Zf:EX	��i��A��(���.��|.�*:2����V�<G��ǫ���E�w����T1�LSM]�+!�)Cv+L[	�<K����Ћ��¶I��5�b�0����x�G��#]��O>�ToXlz,��u�a���0�m(Yv������ϯKd㋗.d	�,ZP�`�5���q2����ޑ�"|[�x���@;��$�q�;��?��˛��������%k���[v��={>�A|J���c���T���Ʌas��GG�`Y�D�%Ɠ�<�HCC�y��
���D�;o����wv'a��`�1I�9���8���"(o�a��L3u5u�|Dج��u�9��(5i��0��$d`�c��I�E�e�9��d&���c	O���߂�(y$*��Ci`R ���
��-�hEð?ض�I�w��L�7����\�@�\�yR������Izn��bj#�����p�8�߯�D��T}$�͙��s���hM]���R��i��Lr߾} ��G7`"เp�#�Ͷ�L�dr���k�A���̝?Wr:�FK.0ۍ�{v�i��2m,v"_t�R##Cc����x	dq*1F�s��u�n>s��M�7��4��Sq�	,�U�kk�e9�w��+V��eXɾq������I�-Y4����3OϞ�q��k
����L�T�tY���z��Ug/�ԉ/�6o�\�xy"�`��5H������?��_���%m��2!� �_��_��.�>�m|�:R�2:K�Ǉ�4M�)�����$$���5��uyi��H��+��S9C�iMUL@:&	�J�"I8f]�L~��#Uz!2+=sb��]]<"��g>�DG��1�,&-�x�("}���?�pl,,]���@))�+1B ��d-� �`���6�*��A���h,� ��D��1eT�uE#����5P�J�P]�Ȑl���]��I�\'�U���+�-��d%_�Ț��Ms`` oI��z������FH?B'Z�v�7̱'�[k��F��y���f�D��l�a#ZN���&�P�75���;o�V���x+���1�Uz�(Ej��<�����P%�?-]�f=��} X�𱧞z
���1V�J�O99���\�����tw�|���)��y��C�q�u��ei��`�,�Tݞ1zO p�W����x<��+���?w�ң}#kV�j
n3��{��7`T�&y��cr`��áDj�b4�df%P]��n$tq#�\Q�Ɔ�N�UD*��hC}u<6�d�������N��6f�``O�@0�`�K<2�����L�����24m�˯̙7�������'���{Õv�H2����r�, �����hTU�ٳg��jkk㸦����ڰ�%z�����Ά�����|.+U�E�f��J���R!�v
�L����p	�*Ċ�U�כQ,<x$c�TB�W�i�Ho�|>o�,]��M�����V���W��X}]#����>��������/|�C�aNUJ�b��.�d�E���d�~��yӪ��Y��uy|�Q�(ǐԞ�5$$A&W(�����+�>]�`���Z��\*'��s�n���ȤӠK�吩�w���p1�J��INֲ��&j���Gҗ����h;j���"����o]��T���d&��İi
�REnТ�`1'�G�C$�*ǀ�G� v��;
9b�YM��2TY��8�s��´d�j����$��pg�T�TB,3��&���aN��hl�y\��jP%��eL�����-����D���j˟&D��;~�V�ok�ڏ�ԕ3e,�>\��T�%:[ںNt� y��fE%��[��ƃ��J���$��\ �	A��ܜzʩP���3���hS�����I1nZ�2x�v�W� lUJ��
jD%�E�a[�������zK��U1���]�奔`%���G��8�K�[��S"2*++GF�o��F��Q��O}
N���_��J��h�FV~����J.��f=.�%2A�#R�#�Or(a6�\*�Aٺ����� �ht4�H�cY�"Xw��胚;o�ě�5�����B����rbKsktx���ՑHO���i��P��7V��b�	XB��C��n��v���LeEĽ��r�T8L�E<��СC�P$GE���y�@$RuʭYkR�u�{�z�D,X�g�P���=К�������ʈ�ι����sƊ�m�֟/�$�� �����l�b*yc`l�L���$]���Í���N7�5�RT�J	ra��ɘ���Jq�x46�c�(R�A#pa?(�d��ͧU�p��P@�
Vr��3��>�>Y_X~��/)��-ɚ�,6�a�gN,��ˠ��jBN��)��䐬Ӽ�[��t�;��I�M��P�$�� m3�����(Y�@�L��R����y-�˱�6�k�Y��O�B>Ϸ�W�I��j��22o��s��XVh&�Il=�Y��NfsN	01��`�6v3'��wf��:��/��UR�!ن��\:S�'3�ρ��4l�,��L�60�BQQu�Ӣ���1Φ� i֤�#,V��NS ���yݺu�_��P�V{2�ٶm�������s��+ 	8]C�j�"U�SE�^�Q5UK�S��
�#sD�U���i�s�ƍy�{3������H�v��Y�x���K���淀F�ƪj���<�
�^�H&)?4 ������w�������E��J����'eB���E�(���ν�)2����\�}z[kk+�;��݀���BW��T6��sjkk`�J�<|��k�gOol{����뚦p�i�$y�8,�e2�����9��cc�.W�(	5�j��	����D��4}D _:Cu��i��
57�$�WV��'����\Uup��끳(���ѡi؊KC�e�z��P�U֬(�$I�6m������(i�Sz�������=w���-��w=��v���3�k�ϝSSI�R�HM�|)+��D���A���c��\^Ir����ЕA�����`��>X�d�R���f��G���/Y����k���-*+��=���}W��~��;q������I�`���(kw�?s`�W4V�c��r��?�xh������s�'h<I�lU����u�ׇ *�D�F�eZb���$"4L��bB+[����T.�ڤ=3_*�%ҙ�şJ�`]�N�N��.���Tؼ&�ɇ�����X�
"WM7X�%��G(w{;�5zz�<�ԽȔi�&�"XV�n�tq8�3��ɚ��iR"ow���F���'�x��v�p�b���ܝj��$0B�呺�fE'u�����0p"J���ɤ@� %���x���8�P�	��cX�����ł�i���H&/���d,y��β��<�׮�A�cv����;�g�7m�L��<caC�~�w~���d�ص{�?���v�{졟�fн:�hX�H/[6�?���p��B��{��k�fěC[-y̓�վհ��`��M�MM�Pȉmk�|bʓ�4L�C5������[��&RO����V������W^)H"@y�g@��St�\UUp��@���������m�X�N��'����D,*I�R1���;w�7��R���Ps��������Gxg�����p�P��%8H���#���R��dt�U����x,_���$vh��Z9X�iIR����d<nw۴��H�С��d��t(��{���pS�_��/�b�K{N�� ,�(���,���łv�WVW�z]}=)����:44��5=�����$�*������ �%'��
���J6z�NU�u/;��]?{�P��3[|r����M�z�.�I�ǿ=����K̥��t\�*\%�؜l�K�{�Z5�x�X����deM��Q`��p�ox$�����0�|�
_׉x��d"*���\���/��T2UU]��fkk����<��
>p��K�!�%�O�S����\��H2Os����*�(t���T��Ӳe7�G	����ak�����M��YD�&��"� 2� ��t8���	,����YԄ�)�ɤ���9d�gt���&�eT*�M��2�s����Õ!������_8N+�|�E]3GH"��O�G*"&�L�˃� ��I��L����y!,XĐ
���M�Pp�n�U�L֑~���>���[^;��':�U�V�z��?��a�H�-�<V�b���fsF`C�8��s����/?�T�>��G�nٸr�����Ǟx@������FS�4�(�����F�����s�c/�{e��u�)4��s$`Evs��׺��B�����o9�:cɂ�\���.!+�An�7��=�Iʜ
��2���rR�$��Ř��E��{�8\��s���YմD2x�K"�x�e�����qrp��J״t*����# �\.��t���p䈙�d@YnIY)�X��\���E���6.W����HwP�*
��ȥ|��(%����C����Ғ�.�L�8��I�8�Jn�E�Y10�M�~tR��h���Y����� �;:2τ����B�'��O�峡��ђEx��
����M^=�dS��G��ƺzG\�����j�\.�D�Z����
H�x{i��;k��BIQ��ﺲ�A|򅡡x��}�L9N��Do���h�����钳�Ԛ�Oaޚ`�L��ղ���0�m��Y�U��a��9�N�
��rJ�Y��+/-]��W��*_x�Ū���:��3��4������]����E�u�z����`_��\_����Ö9|�p,WZxfu�4׺�̺@��|!�e��v��Ոv�Rrl*��y7�Ɖ��dj[���X`�Ám�qc�(E� �y��PO3=OY(� �#ioC*���1��0,�,	�`��̙�9΁6˟\de5�1�Q��"|�cR2[w�!ԴVe��8�uJR�����A�A[çT�t:�,� ��*S�l���(�|��2�|N�Y����5����J_�&���!���l&�E��Ԃ�L��E��5+JL��'�J��&�ܲ=U����"�V5h��K��؋G�w��\n'e*�����<I� B W(�
�l�x����<���T��/����xop�_�<gޜ��f����8k�B���KO�h�Io�7N�]�l��ȃ�_(d� ܠ���<�����5UM���l�������}��l�\:58<t���˖.ܳ�0��D*�q�Ђ��=�x!\A,6��<������9�y�g[�b.OZ1��wtU /J�y'�.q����,�gd@��B��+��rQ��lL�bdl�, ^3yѡ#}$��!~j\������b�!O	��TEVK�@�555�����x�P䜾B6Ϊ�C;^���Fӵ�VqT ���,��Yl5�bӋ�H�yOE<>Ȋ������?92r}c���:5��R��R"���b�=�u�!�"���ڣ����������� �~��o?��3�^��>���,'v$=��`�=O��o|:��ՀiϊI�����'�Zg�s����sW�`*�����~���]�=��y�9�tww?��дiʫ��꬟=��6�POn��-?/�4o����o�u�+V���s���_z��_�w�~`d�}����x���54�8�O&�IƳ�d��SG\�E�|eb���9Q�i5i����d����z(d�@ O�R�CYnx�*	t�P��g���e���r�ie�>�D���u欹�M���U�DM|J��^���M�"�/�	�KJ��C��h�ht���ϮX �u��sB�bX݆�J_$��β��
��>�u��zU�dA�d��
�?��a`3��\<��qD�vB�tR��fهKi�W�ZMy�;&��1]���:�������E���B��A]�mdVSsc��(�(Ӥ���r��n���u������a�ϓ�屧I�7�����]_}~�ˋ�,�3��	W����-;��A�����*9yM+$0I�dLй�4����
 �t:������1�x���v
��t��ڵk�w��_QQ�A�5q^E�w:݀���������ڬ��`؂hV�
̪����`�$�^*)���Ψ`2K���?����ŸH���dx'�I�)�7�Ij�.�"n���CL�(ְ�ma�0',D�������O�8�	Er�x>��9������ٽG��W#tt�N
jF0X'�� 7gvU]�А��^���o`�U"�qMm�J&s�{ޛ�g�	F ���l���}�^q��%'uۭ������K�Ǔ���A�[
UΙ1s�\�Ys�"̆n?5c���0��� �9�L�BQ����>y��P�8��ۿ��/���Nf�g^�V�4�X_�\��<:�>�LX�#)�闶M��Mm�w4��{���]tӬ�9C�>�͟�P6E�ɻ�����Ysi_4y��6���;v�I�&�*:���2�v"��!:����t��i�ͧA�lG�U�`唞��MR��W�P̕��>'cM$�
;
��0ʯ���&��-�D��w3�=�%��$��DM[��AV�����,1<W�Yޑ�"|[�<��x�@W�aW�Y����AYZ�buK���=�Τ��c�8�s``S���P>�ͪ��f�%��k5��9���e��f�,��L����Π��yV���E7��2@EjJ�u�d�n4�5�  ��h�<�%,��s��bɢ9{;�_y���Ib���]�h��I��NB6S����r����[?;2�������zA-�X�&����p�Mm�~r׿}��������>�;k�}GI�{j2w����*)�^���g�iU��6+��Y��h8��;пk箪�����뭉��,�ꫯ|⦏��8|�HuUՉޞں:@��l
.��o��t�w�Z�Kzm�N��g5mx��sV�+J�+��^����П���#�\n��� & 8;z|��3�Nu��U��x<�?��y�����袋[[���͘�P_���%˖54ֽ�i��U� "�����s�_�ӻ~�>�c�����`ނE3g�>t�����P�Ú*:pX �`%������{�.\�.Ct��G����b��v��sϯ���۱�m}�-�M�u ˊB&PP)wIgM������Oe�����t���j<:�.0�|a7�/U{DNp
��bE�'�X�pA���M7~��y+.�h^6O�}�ߞfΜ�h��?>�կ~�����B��-bb�5:�LNۢ++B��7����`����<���ݒ��j�����)9�_�����G?2T�����c��t��Xt����(u�����S��,��_߷b�9�t��Ci
�w;�.�p��H����#���C�H���Js�d�0!���b�$8EIU�R�Du�N��zo��Tl�L���޴ßVؘ��wF��ݛ�ϕr���%��k�i.$�|������`C�l#��e,~F�"98Ȕ�ı́���Ϋol:r|0��641��0`��$]�2m��P)3��;�;zZ��à�<L�V?����h��#G�v���;��qzL���K2dh����߈���N�����(T�xJ�L�8%�sv��|��kB3XX͐�"�hD��U�O\!ER*�;�UAEc��X�K�@��Pv��<hCs�bM���E���H�B�A�r��_rI��%��x�V/kT8T+3C8�~��7�8
�.t�z맺�-����&��O�^�aT��\��ߠQ@u��n��W_���A)�2�` ��ڊ	�6$� �@��[�$�;��`�� �|>��p���1C�� �fΚj>��O��0,�6��|����������Sid��$���s:�46΋�p8���8���:_,J.�����r v+��K�
�5XQ�N�܍�>xO�wH���%�����E���#,@*�����(�O8���
�� :�5���͗��0�ǘhK�JV5&Q��Y����K"m�bt�Gˏ�M:ܾ�YD�(��3� ә(ӊHe��Y^ok�D}��k�"u_��	�h��T�	������Y,R������>'���擤c��6ӂ�ٶ�������8�Q�y�����	�7��E���3s֑����]��������m��^�����m�m���%�]�o���vX~�5���+�Q�)"��u�*g/Y�����pWТ����gL'KX�9��t��g,�P����PUm2�t23Ӵ��O�)��Y�������I'z�as%�qK�)*�?��o��n��Y�@�:;/��������� ��Jf�MBܫ:���;(���"|{c�*� ���i��:6'�l?E,6�ɤ�;�v *b�%E�?�V֦a)�2�2�z�+C(�@�h���&W_[�Ғ������.jDE�c�*\#v$�h��J�4"YD���ߑ�74�w���0V����̂\b�=Vjö��z���7ɮ��{�����BM�;.Y�쌳��Wy�hw?F�)�ڕ���#{~��M �?q�'7oXh��U�Hk�����=tj���;�*�%�4����8@/�M�M8V���T�U��7W,�V #vu���7��P6 b�B@.vv�X� ��I���	�	~���uvv�ƪGG�۷�6�cfww����y__��-[����w��}```ǎ�@�����+��Mz����f�:r�ئM[��#G�>����w\�>Xqۧ�����������U5u���*���&����7���������~(D�t��U~�?�J�^}^mmC4E�L�N8<�l���9s%��
�1��$ΪA�sY���%SjI��n�m���g�yB%nX5�|f (H}XXS���BQ�5\S�-'�=Q[M���{�	��u$��
������s�>����/~e���6����'o�Ȭi���fW�ӓy�U~��D��`M����R�
��[_����]�<%g����_z�)�Ȇ�Ԓ�3׭_��X�P���7�.��sۦBv��-�����!�k*��޼^ȈU磺��ၮ��Z��]?�^ɠ��_Lo��Ec��PE^A'������!�����8���3c�'�x2Y�Iy�LM��˲�����Î�]�E�r��/؀B�.'�u��YNWؿ�>U�͘hĭjr������k.������}�!;G'&��|�Sw�N��?<0��x/����u��gy�c���{c�QQ<�P���8�v�JX��j!L�4A�q$1����<��Q���g�3�a���
C�.d�@Xl�$I7l��h��I
�.j���Q0�\�j>t��#�$�Hv�nE�x02�J�[Z��\|�Ň�'�#Y�հ�����ā�7p��{�)f�H��g�{���Þ���k�2�����{�@�׿��[�}��^0��k_�
Z'�6ӊ{��Q���E�ŃJ��i�"��
��.+D�������e�V����,���u���/���Dbpp�������ﻯ��._(�"L�R�a�a�>D�����Gj�"==��l�(����-[6<xpp`����p؇~����;��/�����W]�+��/Z��Z[Z�EO_�SO=544�m<6~`���~P���7�4}z�-��'UU���o`pPf:��E�|�I�ߗJg#����f�y]G�ut�	���\�3�MTtlxtt���w̙��y�����H>D�,��s�R[4a9&+�ȿj� ��z'��s���-/h�D>:T*f`�s�C�y�[y����WP�W����l:r��2!�뻟:p�����g�T��D�����3g~���Z}n}����C���?߳}��'��;�R�f, ��um׹��E~X�>�빸G�
�PԪ�8�,�������Oܒ�ښk6�ʪ3$�U�n���Z��}�[y�J0i-��u��*�����(�������������qq����|��Zh���1]�q?R�#���ۑ��M���I*a��U;i�z'�|�X����v��ڏ�.�(8���v�(�����pz��ёQ��FFGC�)2�J����y9��AC�c���B�Z�O�3}����j,i�β��gA��*�ʹ2e��нJ_U�Ky�*�4W�2���CCVr5���u�<!SƮu�X���
�-�"����`0���]nU5�Ne-*_��o����"r�� &F5s8Aba?:��	<�%ڷDd%ܗ��@�r�!	2Yԅ��bH�Q��`��m�4���'PʳfN�ܔ�PX]�6o�G܄�5��4Yi����R�mm_��g85����N��1�1'��d�����]T�VMC�����䓣@Q�\�h��,I��e�}�܉x�	h��+Wf�)��p Kʸ8�Pᓟ���w߽s�6t~o`tE���`�GGF����:��lo��-�K��-�����fx�	�������4�3��#�hG��d����f�������<`)x�N�-Z6L.W���`�Lx��v���ܘ/��Ɯn��9�`�� �CQ��"�x��ښښ�0h �z�~EQW���4��E����KT��{����7�����fy������v��7�ֵg�Сׯ���[G�����յ��=Ϟ�r��U��C�D��P���~���s0>]�p>���&O������O>���uuu��֮Z���u�D������0.i%T�Kx����8U/Z���*be��௹���j*��|"GMG���틟�����Q�Y-�p����Qj��vLd�%����$�褍�]�>�����5A'U9���UgJNG(����K�z��k���������*E��x�v�]�3���e�1�����!�O� =���WNO��`�B7u����ں���`�h�P��rp�A����x���~����/�b��ۿ��#����R0�B�HX�֮��3�[*}���F�Ͽ�����X�MLY��NSvꪅ(�w�z<������ٛGD�a�J%0��q���L�B�p�]?մ�,�e
*P���.�
��ǗU�{�)���}��w�$^T{=�$%�1�0��H%�=j"FhZ5��B�t'	M�<v�MО@;3_��M�?�}w�dU��͕suu�ݓs"�	bD�tELȮa�	�]]W]3AX�+A�3�03=ӓ;wuwUw�9|�{έ�V��c�3������u���}вЮ�,tW���𽠆�A`i���G�s����x`l��;;;6mܴy��.n�9j��E�&rss"/:��
|�'�
	�)V[��v\ �&�Σ�:Z�jSHEN E��E�-�n0�u���֞b��*�?���]~�	2K�Z�%�*X!�dtٲe��H��/�B�9u�M7�x��*'Ip/MĐ�` �[�w�*v_�k����ٵ�Zj��NK���i�~�����5��b|���a��rN\�ёq���B���#�)�jeR�̰�ȕ+E��ΎN�VT�Vݵ���,/9��J�z��_<�X����O����c^�)g�'�a��f�שxY/�Y=痌h�O6v�TK7��:;:`={<L*���M�|����:�����18�R�(o"�4��[PE�(^]"�7Ò��NUJ�G HCW����N���΢1N�n����rm��T
\[�ׂ��Ҕ�[�T�sO?	V;�f��^i���+ �9�  ��IDAT-[&�.:c)�~y����6X��	�
�-XW��M�����֗A��v�lK�_�\.gբ�p���ů�����*�\>�NË�PAl�!�.8��m��iiiy����<|I_W�P��L�����$!e٤J�Z7z\���pu8�A^�w����c#i��O��Ɇ��'n8x�@��S��$T@H�`{;�j�cky1Z��ʄ�`̓��Y����23S>o���e��Z�������4�,�Y�X"��v����B���px�u1���:��e`x���P�q*Uu���%�;���0">���BHr1��^�;35u��]gE�o�������P���o%�ޣd�{!�P�����"{<�4d2�"qz{s�Tѫ�M8���Ȕ�˘�`Ћ�5p�	�~�B��AL;���t�=w�0�GbJ�
�=A:V���%7p-��*�y\��=Wֽ�Z����!ƅ���87�����H[�*E�5�3��	�@�e�T�����$5�Kc�5�M�����59��[E�hDK�	�����ꕷ�u/8=!�iK�w�*�Z�Q��dPb��T$�T��j:�������:BG{��~�������q������jko?s�馉�K�������c�S�DLQ���Jc�Uԋ��G���Z�$o��27�sY31C�ߝ,�q_����IMj<�1ʑ�8&��0]�޼���jܷ��+�|>�����r�/!���U	��1�t�Ѧq1�0o�ڋ]�(B���^#��4��83$ȏ�����
��Xx	X�HƔ5���`AV*U
0+,�[��z��@��JetlL�2lu��H��`!��"���;����z���<����_����|��imm��F��{���ˑ�KGp��Ķ/����83��w�0��Ww�h?"����4x���lf��Ȧ]��g�*d��#[���"����Әa��Zw︁GR�������s��I/�a����⿹�W�}���������%W��m�����7�MT��&xjr���߰,�,�.? A
sѽi����0���n���xQ�3���L���ڗ�ǆV-_q�'?~�������y���?�7��o��M��r���Ǳ�σ��ED:�W��)���`�#B�`X�����ԝ~!-��h��`aעa�r= ���^�\�jDl �x�|f�n��U��rJ�P��Z�V��!�8e.�p��iQ## 6��M����"<���6��9�sx��;hk���{z�������/�Z�uO0\�t�󪜦s�\U��N����c;w��|"����>aCx�p����hC��?��&>��OC�M7]��3~���?}��D<��?`��G:L�֏��Z�j-5�&��! N@������T4!�q�%U����POwOa�,xн.ˈ��R*ۦZ�AI��#��%�6?��t��_�T�=����Bժ����C�@�2�FJP���d�6"�SLf1gȵ ��7OO�C��"j_QT��$WԐ5C�W8�\\�W^���566[6�Es$h__c���������?۬���ޓ+T��Yb��̳Ϋ㬾�qE���꤃v�RP��ni��g��ǁ��{�ǯ�+է��.�k�FY7����o�G�ڿ~����8��\D�P�#f����ڦN�k��L	��K����ZM.��As.T~�],���y}!O��w=�ࣩ斾�>��o��}���?~|�unlj���o��7���������j�i�w}�_��}�m���Jks��C33�N�i�b��Bw�{����//(�x��1�k	p{w��+vC׊�Ev��U���H,
�l��1-T���J���i��努[��o������wO>��I��{V��kn��{�O�w�������Я��K.y;�h�rF���-#k(��H$��,x~��������I�U"�o�t��&۴k�u%h��m�x�ɦ����O˥�cmR��I�u%�`ۖ��_+���GSTˤa4��9���+�VA�-�dˈ�# Oc�hzj*�҄(ܶ�Td�vx�<Gj�x�x�6Iy��pa��կ�kKs"�=��s�2��c�X:W��A��ص���+U���}���)��Ƈ2��#���}����_�vt$m0��1�*�w��K����ٹT[Ks3+��+��7�L�⋷�
��/��������M�b���g�`����l\�܏2�Ih�؁0ۑP���g�1���f��Lt���u�r������t0�A�~������z$�b".�M�)B�渀ڠ`� B�=�H�wԅK�-��` L�7�D- ׼��g��L0�
ef�����v(�����&&�� �jp��U�����2�ڀ���Md�:����q}�����[�p&2��#�!�Y��ҕ�����|=�e�G�������%^45��m/N����S�ę�Z�@Bat`L��E�ȆB(Q���=�r�!���Q�]ƱZ��C%����v�3�(yM���T�#�����g>yçW�\~��w������r9����߿��o[�b���k�=]=�>��O=�����w��~x�g������TJ�b���b����ָ�h�^��LL����U�����[�:�W�>>�/�|���L�_�e��X��ބd�8D�IP�X��}�C�b���=g��a�������״u��X��������=t�����	+��3m �EUVf�A	f��r����^�/�L2�A�Fzߘ�Z�|��T
5�Y��z�bH����};� RV��88Ϣz����J%����/��/~+���X��mv�Æi�����P|�.��A7���"T�c��h����?�E�"ê���2�}�����@C_s�
2�P��,�s-ݝL�z��dD)
744�65'���l�f!ˀu���;w�ģ���{Ͻi�|����g��k��ލp-����۞�q�Y�G#���UG"1K��uM��^I_��݉��|uH95K�u������WG��I\�٥}b\�a\%�V(;$��C&�[�k�#��N�#$��`����5��������{��ҩ�~��+�Cl5w%��c΀}T�迹�Hc{�úlX�?�'�.$mycBoW��i,{,	pX4�h�KF4���f��̀5�qݺ�v��� t�e�~4VF�hS�a(�>���{%n=�r��u�G�S���vxR�R+��g�@���풀(	lb�Fgt�'m������ٱc��g��~��JU�-��|��p��n����yv��]=}>DV5�\�z|awo�E���{�-��w��gي]{���AI�J��{�F{��R�X(�
���wa5L��iI�_��f�^2�nF�k�C��(x"
L4�/�f�g����. �4�wՏ���w��zN����f2�����.q`(o�iN���R*��`1�[[הu��\|�O?��7M�:��7!Q����뱿�F(/]D��|�٪\1u$�Tʭm͑H(��>��lp|1���>�R�g�Ա���b>���*E��#1��'3[\�|���q�Ù�ɡbz8�53#�´�=.���9�|Q��	�C� 8���ؚy�i��c|__�y����u��ki��}WNOfv�?�W��Lɚ,�1��c*�0gy�V#�@"���.0��J#c��/b-���v��k�f]v�Z��a�˕iA�{l�bi�]$���˹�?��D�u5�8~�	�l�� ɑS,P�&K,px-�r2tuղP��y��_�i����Uׂ4�A�2ΏA�h�����|��J�����q\�����W������O���G�i�#�:(3�}\�2){8��c�ʅR$�"H+���xH׬%0�+8	�0� &fxꠜ&�B�hE�N�B�tt81�&(f�8�<�㐖&r�<��ˊ��d(GЈ?��ORM�ݽ6n����/��n�����pXp%��z�G'�B����d�x^�$b���7w�����Q-�Nٸ���na֑%�5�\��|���aqUk���Vl��-��ݓ���ȹ�]�R]F7"����D�Wo{Y673�~;_f�����穆���>q�;~|�O���n�k������ّ�	�o_�_�*G:C�fD�!��Ҟ��tz�����M�^&j]`�z���c��]���Ǳԫ;�$D�ڄf�_P:XK`��\,F��B!���pιg�|��mc���Ʀ�ޞh8v�?�#�����"p�mEW<�P�U���a8��Met B"�6&I�m%���A�\]-e
��.���3x���R%A��R��@�"�}{�~�_:2>�����W��;�w ���^Og���M���9g�3��y=h���ٙ��კ�1Ө�s��o��=��JME��Z͡��,Q�Q�GEM,�T���+Sk�n�;B��[?�C���,�Wgm�cP)r����n;�v���u��ČiםK���5AP��bZM�:�'6!Z"'Pۅ#��/Q�� ؎A]]�>(b�����%�C��x&��vx�\f�1]ɼB&��2�+��4�n�v�L�oɮ�O`�M⤆�X��B^B�����
���H�i��U�Hc! �9���n�I���(�p�:���V�A�(�F@l�&h�T��
�b���7�[����8,q�%ےz3˲�l��ڞ���\����l��Yr�]���y�Ļ:z׬^��w��?��(B����3�~���92����,Y���*���o�.]��+��G����}��w���@F=�Q0��~�?�=�����dc<�*���z�����P` ���s�̰S�4�%ՈP��%$�h\�"!$0 ��)��:{�n��'���֝�?3lZ�贱kϤ��^}�k�Z����5�Z&'5�
��9��&�\��\)�J�eS���F�n�����D]q��_&>h��<W���Jv>����,�HZ���ia�����d�O<q���%������Q�ǣ�������ka������0aQdK������~�;d��7�n}�Z.�w�E}q�-k�5�M�wln�E�U�O?4����H��\q.����/衍k7��T&3:;�#���{�X��5;e�t�|禯��?~�s��<�K����\|���_�ǭO���oz������V�l���ׂ"�2X:!��.1�� ��bi����9��C˒���M�����A����Ylh��������#h��\�,k�Z�6�u�'�b0�7|d|J��4��B�����?�lr��C":�E#E���q����s�j�Tpx��
`��f�f#�ظ�r�cя�	�ld���԰�p7��d0LHU �[�(�
��E���1%�`]���}c(���6|�G����6<��ÉXL�uX�XUcZ�u�c�!�4����Ĵ����D^&��݈�e!��A(	U�6��\�C1J��B��~�H��8�x���r�B` �i���F����y���/~�Kg�s�����f撍)��3<4�<+W��|�i{��D">���'�4M���Ç���K�<��S�\{mKs��ǶoX���w���������6���ζ֭_��O�z�	�bf���]}��
�8Jb˩����H���������a3�):��1����y���}��MO�YC/϶w���M&�ə��x��Y�_s�F}Fkn��
�J�p��t:}ƙg�ܹ���Y���E��^��GyԲm��<B�/t^�Z؝I��/�$�a.�:h�=<!�I6�l@�z]�LOs�x�%Hi�@����I�$����g�Z�����/1���Y�!���׿�̀��g��3��֕�'"�p�h�Ceٲ�+��ͧm80dJ�\z���FW4���Z�hk��i��k�㾻o���J%��+�������g>37W ��k�ӛO]/+L$���?�s�!�?4����xTs�c������fhD�r�`?���h�ЩWS��#zɵU�Ѡ�M�"\DS��2M�=�<���>��5��{D�Ե+��%���?���J���t�[�|�_$ɉ�|Y�����lU��G��=�����֫��ZR��b�����6��U���N�jL4��))��j��e	�#���b���^�l
�@Mx_>?
F��ULk��U>��D+���7�8�_���H&>
�n�&�`i���tuw�I6��ժ��r�{7y��Db<��R��RsTG"*o�:�'��mm�`���2X��"�r��L���u����i��뛧0�npc,�PH���`�������?m�
V��%�����S���j��.z�y>oZww�a�^����i��^xzz�����4i�DK�4M�֞ݻ���E˒�]}ӣ���Yʹ�`��q����W�ka���4W����P����g��4�休���'-�EN�fgXV�50��͋��i������t��� F1\�tz2��kJEŧ�|�G7��,�B H_,g�L�����I�w���<����!�n~����D藾���D\�ˬȝt�I��T��4MMØؒVKd,��+�/�zl�7��/{��U۶��j0�/y�?�zl��0�7��o�ҘQ���^�b%)��	�^G����z{GƳs��j3M�ɓO]g(J��\���z�o{�%�����|�ѫ?tE{gÊ�sss'��h��&Nd.yז�yx��˼��^��7�9��j&#^�C��<�w�}�6�s������2�WH.�
��dg����5'm��u��#O<�������w�ھ�ݗ����?��;��-&+y�q���B�X^c^��9VSU�X 
��Y�e���;;;@UU�ޝ�T%�{�*�?�0C��`��3S�X$	��B��[�IN��c7PPp�W�P�?4�+¿h�u̒��b�� �6{�[F��g���b����K�kSh̒cn�f���uX�6�#�ʐ�C��A�@��k<TU�����k�N��x�WUu�E�E{�e)�* Dܰ��	�Y^ ej�f����N���͠p�P4�M�xϥ�T*�����sF��Z���w��٘m
g��|V15�����~w�	',�[T�����3��B2��5��`Kk���؝������=�,�I��^GL�c¶Uo�_0�n�g�FhV�4�[��0�Ҷ4f�*E��5�>t�?�spQw�}��;v&�\ybφ�O)��Y���.�Z�P��U�Z�f��k�R�Gc�������4��䬎/�.x���/�.f�<�~�4!�����u1n3"K�#i�����+��C>r��/�~
����u�~��ބH��� ���*m��x$�����_�1�cz�w�{֋��FAŒC�X^�q�0��G@Uē&Dkjfΰ͆�Tw��Ds��H�ji�/_���+�z49{�����[�Z�l��'9�#�m�o��t�)���Ѵٳ�#��~���f'���泃>&ch��w��c���E��	I�=ߴ�o��as��	��$pC�+�:��M,,�ԈG���5��)V�@t����l�>�{�D��퉧����D� 2�%A�B�)���D"��,��F���U�R��QҚ��̡R�n4�8�/��>�q�ڈ������ZtA���zA������X��sုP*��^������kG���sH�@��H� :[�X*U@��Z����#�bn��Kz�ۂ�G��l�fт@}AV0�8� �,a�.bza���C�ϋ�v�����#�e�<Պba�;2����JB�H�(I/V���k �E����f���U�>��H�Wr�*���j�g��K{f&����5C�lN�"*�b1��9��}�郃�o��'���߿jŒ뮽:=9�>"�X�D�*�������\�=#��Ͻ`���}�֊��`�
ıĆ�U!4��<8�j���%����;�	�����ʅ��������s7��>��# �T���T���[����,B V�nL5"��(�Y�愍'��>�ȣ4��,�M���%��z�t�棋������#�/���)`�P��"P�e��I�.�)Y�lX��X.df��s�@0@�6,;"3LXS�@
M�����
�����r"�%f8�|�_�w���Y��a������%R�����};3��F2�j��K�2�<a0��ɬ��s�:��y��#0�����OL���u�|���;W8�Z�{�ߴ��'�}d�i�\|��g�9w�m�Le
?����SN���-���m�_r
��E,_DR����e��f
�����t>��r�Z����;�>��R.���y��E�owK�譤�#�X�J�-�bݒJ�1��|���~7x�nl��"O4�AMc��T��k�u{�~� ��)ǽPȃ�O���1nC=3,k�A�Ѷ	���uHt��~�3��(�Y�--�=^�+R,�ll;^D	�� m#Ǔ�`W)#�}>d�YWS�4��4UUo�aN%	��_0mzj�=�m�B~�r���q�֎+��=��M�c>!�_��\N<^�/����'Pъu�R����kɦ^v��]݃r�2&n�b�����z��8������� ��E0�a_��
j�_$T�n�ϛ���*���i��%�ұk��8�ǘ�NI��A9D� ���%㵤 ���l���%}�X�ٸf]wWo<9x���Ь�qƄ�:2|�)[�l�Ygl���H�];w抅�ɴ��$[�,����n��3����Α��p��,J񄧂�H����Z72�����Vw�ʽ{��J���~o��0gJ�c�&6)c��/Y��v��[\K��h��|���+���Đz}�&x�B�O�����8���R�M�-D�GQ�X#C�
�vá|r�H�Ik	�3�oT-�����oy9���]O���=�_�ff̒��ʧ��e�������ݼ����n���%ь��@\�ƽB�1�Z���TC�C�]&�x�4u ��i�QYƄۍ�ϋ>_�WIw5�#~��p����}�ȑQ/�Y����g��;�46D�j�:n��X�XZ7}�o}�ߴv��LL����}�럻�{/�;g'&�㮖k���}��]���@��;d�3��$,\�t�S\<���b~f*�y�z�����|�;��8ޅ����[G��Fc����LԼ"�"�'��+�#���e2�zô^_{{3�eC#C�ǁ9]{��T{����r�0�x�~�t�n����l���+dwΞ�I��ϧj���d�3�8Z��"|M�%���Ǹ@ 4��NO�r5���z����DgqKOf*]?�l�$�IX���&��n/���$�@b��d"�5'���gYN$���">'U~<;ϽR����+R;���)�3M��i�(:�z��*lJؽK`�q��*�D�;���j��z6��#aa�(��ݻr�¦M'~�hki5�*�J�b�Y�3�������$��p&�p�ZU�K1k�a�r<Qb	��_��W_|qgGǑ#G�ႤP�)*�/�D��6%{BަÇ���N=��h41=53;c�J �P@D�,ۍ��55�A���|zbb��/�,ko������?	�0������㨼L��h�8_kJ򥤫ͱ/��"p ���g�$���+	�Hg� E�F�^�M�����O~�pk`V�{��m�;ﹿ�1��;y�=[ۚ{:��j�����}4;[f� ��Hw�-H�?��b0�ѿ}S��?O�@@K"���J�ԑ��m����
��#rjЮL/mooI&���bXg�}�m��q�e�*�o|�_�2�j�`iqzlK8t`RQ�7�3�q��o�ٷ�������-��\���x<b���r�ѓv�piLH�Ţ�K�V%[}�]�����'��uv4�������[�,�����.�4U�6x��	O&��H@����3T������'��E�V�sP�)�����`�<��tv�] Xx�#�P�'`�^�B-��+PӖsɘj!�b�JYLD�[�g&�rU}��S�|.�"�Yx����q
�+��=�c��<o�*���ݥ�y�Q@%U��q��]ob}@5p^�V�L�<:z�W"7v/�lGDE;�嚛[Y���fM���)N]L�!�Fp4���h۬��Hx�i>΋���H���.�|�ņ�-ɟ^Q�44GJ��x���?��G��;�-�]����⬹~�Z>x`|d��@���r�U�������ю�Z��m9����K��0��H�6�REQ���0�u�SSR�C<a�ɪ��=˗�/�
=�=�-����,'d]�0`b/]��0솆F��U�W���>��SL��7ݭ<|!����d�m��u,���j�,�T-z���pE�2�%�^Q���%C��0�g�9����n�l[L(��d�7��Z@�=�����ӟ�8�\P���|Uv)�k�aǑlp�9}��OHF��@Xw�y۝z�U�G��H4��
��4�Y�-�M�1�4Ɩ�U�Zn�k@׊�O:%՚1tX��UW]5�sG��D������sB[k��/r,�3��^+�`�����������˟��v��1���#�ͽ0���9�6��'O=�P4Y�����/(L�o������;~��uNݸ�ٷ��8Fbm/L�$�����=\ ��t��]ltT��!�nh�!�Q������)�\,e�YQ	�������������я~x���'�xr`�n�	�	ł}K-7�l�>)������D(R�ȷ�~��\��g�]��>��������kN����j�����e�r8�����{�[�,_�lv&����T+�b��,� 3Q#��jBtŲ�W^y����.�а��qc]�Mh����������|8��&����B6 ��&�	�'���A`��+��}�i鶩�|�va��7�nW�x'x���K�|�����hhh W�"+k׮���l���m��8c��"�@wgg*���˗*e���KB{kcGG��=��B�Z��t�wI�i�-C�`�[�j:V<���%?�/�eP����οfffIF�����ggs���{K�%��ćt�L�`/�
^�?��NJo�X��L64�śx��M+�3�c�6Q�����U�kR�$�Y{+ū��Ɲ r�`�WJ�v&ғ���/���R��Ru�����q���e�{�̼��&\�[�pia�?6���Ǧ|^�R�5����LCc��O|,��޶=�L8�iV�L��g���Kޖd9����OZ[V��Z�X.��e�Ek׮=��-�ɨr5�N�S�ɨ4��?gzy�B$��p`��D~������1K�yϭ���ؓϬ^������]۷��m{�;gq$���áx:]�g�J��`e�����t������{���/�}����15�6(BX؄�b�̓!�X��"b�Z"��S7�:e��o@՚r*�4U7~��k<�^�[�E���1��B��Z6g�
L�$b؅wx���c� gܡ�f�����5� FH/��iWJ�m۞U
9��ȏ�}X��,�|���p���������P(�QY��y����d,��t���޿�K�'��?��/�Ţ%fh̶X(�±?�,˼�qE�:k��_��CT������޴�o����~U�Z��6�hX��_E��m�L��<�ЃgMt�E���o� &��ؼ�h�� ��9Q_��HD���n��w_����m,MUep�xdY��'j�a�%�E���1�]lF�&�.��$B�+
�Ղ�NO�◿L&�v����S���G��<&���;_�@�W���/�+�47776�·�h(+�O�!�e�Yu}C�Ć�:g$�g������?�` H��q�"���>T���t�d��^A���LӠ͝�Y �B`z��J4^�j�c�=a�A^�[���j��ѭ��Q�7=2t\m�$t��l�r\Ξ}{f��ֶ��T���)�JQ<M���7HΝ�1AZ�yǊFS����>�ɏ����W�4G��dLQH%R��<F'�T��\.��\���兰��XMVO]�$_Ɂ9G�^�~ooo��Laǎ�?81���<<4�����.x"�X�X��u r�s����ݏ��W�q��s٥��<ѶV&=�����q��'(VkK�o.{�ǯ�j �:<�5���~�[��mY�����ߚ������3T4��y�\��<-�p#���>�oh�d�X�"�6Ml8E$'����c3"�
����\��InC7IO����X��W��-� 9(�r�
�q*���p�dQfb[W5s mfGKfL�K�P(MOϴ��"��(ʊBJI�|6k������:���H55���+.�	������"��F:��
�
�BA��#�G��l����*�uc�V�.ꚰF.S.�w��=;;
E�������$xB ��Z�-�V��i�b4D��kQD�V
?����ݕp4BCV�ઊ��
ు��@#����-3. ��0e���)�_Իc��s��kV����� %�ޜZ�����y���jkݹs/�b���Ѳ5E��ah �AU�1x�M�9<��FO�NuDun0����r!�x|���q?��A0�)ym�W�<��7D�,y-'|I�h�5���(���>nnj�'kW��B�?������V��f����#�cՂ1_���)(P������U+W�D��3�٥K����3C�j�����&A��������ΉZ~��λzbͩg�M��d��m���ML����	��7pZ|�j�BV�t�~f�ǘ���E�o;�Hȅ���a_�[-�cve���[~bl�ھ�ζZR��T,�*�w)��&t���\~�������>�{$8{0�4`E�)�%�tbgKץ�\)��5W�3�ٯ~��1_�`���s3�x<���K�AU��Zv���*�_�rܝ���	���e�0[>��Dç~��g��}Q�5��eQڎf�a�F�����������7=��3@�Ui[G!$�G̍s�B��U6-����g�}v||�R-U�����1��PJ��c���j�R~�?�U�ݽ�o�F����F��_q�:8����Cb*e��m;���т���	{�n^�b�X��\sM�RY�d��j��˒�o|!8��f���d���m�q
.(h5�g�p���>�(Gpg蔃����������(�A7��	loP�����m<�g�������񙙲,+�]���lC4|߭�><8 �@G[����p021
f��r	N�Me����p�'�|BsKSkk��~�S�a��4M-j�B�`:"����)W�K¸�W�ha�ʦXe���'&&2�\�t:���n������_�/tI�ޞ�b)?99=<4��o~�=<t���æMK��T"���1N�X�Gb-��	}G�VG�3cKvh�����#S�eg�fw/�(�����wo�:��c�����6x�iM�X$�>���7߶x�df.�.^�$���\��QyQd�|YW�;�ݫV�r�r���r�x橛l����Ё1,�+46�s��me��C'o� ���������J!gU��\6��+J���+V�|����Η���U#����1	�#	ΔyF�Dk�Ν����
��N�V������l7��켾M��m��fXf��_���{������e!���Y�B����ޱb�R8�\�657cq,���1�K0�~�a�����w������_<������L׵�̃��q�qE�� ���Q�$l8�P�޿�����;��R�pVh��	���G sdC�2��(�j��rT`~��>
C�����W�!�|N�ч�u1Pb��ĢaY�L\��&��I��1'B�=g��|d��C=]�##��"��~�s[�>�����?�e�CC�Ї��?~tӿ|}d|ܾ��5$�-�Mss�b)w������7	ɕ�o~�k��!ilh��=61y����ʕjwo�bX�d1R����%KW�*Uʻ�mZ��i�DӘ��d�"yJ�VgT�ZYЙ��VUVܹu��4���j(�O��$�庘���:�,�O�JC����������Km>���˗���.��t�l����k���XV/K4����>�e$_���.�m�R�Ik`"��/��6�G#`��l�s�"�[�l���(`,�jQDRjEG��8�䕼�bn*��blڴq��!^0C����gR�����p�O��J��)�J��jO6[Uz/�M N��;��5�r��g$����m6�M������Ke��}֖�Ru���N8�TO�o��s�<���n�2w�[o�Uazn��>AJ$D��MʹY����P�s�S�������;�	����T*��[�r���*�j>�ߵk`Ŋ5��p5D��w�fr-��%�Nj%�$�`#\�mJ�(pU�,�;tp/�b�/�L�)V�VtE�T�����#���ߖ-[N>e3�#Mx�v��!X���t�t�% <��B�BZ-Wdp�!��J�eh� bD��!X��B>��90����9?ܞ��I�W]��`��+¿�%��M�v�T�S��82��$���P�!��e/2%�Q� �m_zM�����0��W\`C�H��8��V�}���/���7o�V*�֭����O�e�TT����믿[�@�h���˖-���[>�J%A�c����u�����V��I+W=>knv��5�ZC*�r�#�<�`��Ν;�@`ͺ��iz�`�n 7��y���j)1��۬��hm�#{��ٸ~��mۖ/_��޾bŊ���_�^�6�����6�Q��<���ׇ�����7���T�8�hh��`X���Su�Ej�`�X�붑�a�U��-z�O $=�9<<���7G�$;=5�朰n��cC���
�����/�+Wm�V��l�t!((H�|a�27k+�@@<eE_��,�EAQ�qn��Б^���Ҍ<�F��믻ڡ]C�0vxD+��``&=�&%�W�������_����W�G`�i;)dj����6%oH�l���&`f���$2�y,�+ߩ�P�̌,l���m>u���P�R�xD��9ðM��|>/Ft�Wk��^=��Jӈ����p3�۱#��n��!��E�cE6j���|'Rmy[ւEB��mT��.�
I�X�=���/t��C�BX�����&q�@�՚4�ɠ��r?��#z먰�K�N���!2�M��4S�Q��뭗�,4�x�(�#��9����7�?x��Sߤ*ZOO�����\��������p,�/V}�'�|rMnr/�عb��%K�/^�̳O���D�#��e�P�	H����(�r (ţ��~�#�d��~����n�4`rD^���@U��Fϐ�ZP�C:Q\�M��Ջ.�X`�r�=�H>_�ToD��0X hM;�!�m�����B��>���?���`��d��Z���}�R�h���]_���;�A���ɉ����TS��!v��$&����S�H3"<i��k
K��p����.k������h"��d���;םt+�x�?�*��0�R�4�ك=���p~�=93]����b{����m���v����bI���8�������󖭏n��1/U�j��n������5�(�V�]�w�{��U�*��W���;��7-��Ue��	�+�Y�.�/���4��~L�u��L��oE߮��,����l��#A����8|�p��L����)E�e��)���Z������߸acSsS�T�D"`���"�;D�.�𴂀���x���e<N�b�1H5O�1�e瞧<���I��"2o�� s\��îQy�<��u�؀�-p�4���xHs-�8՚m��P%Q��f��Ȧm�!��Oa�����+H*�H�Ю%9ҪO)o�I8�rj�$�HNئ-I$u'���,��'��R�rZO8���m������zzz@��\�tæO�T7q_Ec�b��Ć��R�Z���U��U�5�kfzRWTI`�H�盛���kjmnK7��F���X��2R ��=�ukGw���{`vM¯|�D�m� X:�8��d�hIGd�̶ `�4� ��~6��!����N�t��K���3 ��z��3�����}�q����k�����	'��&��:::��u��%85�$z-�������`t��}�HCX�m�h{��!�aAp����٘$6�4�t)���BsKz9�V�$
`:U�1ֻ�²���X0#4$��Ɇ4X%�2z�0�
��V�nok����MOOk�%H�F͡##���B����+
�c����u�2L<�\n���1��;�Lf<���X��xKI�ݞ7��g��5�~�-ǅ� tiLKKS�R���J�LLL�
%U����p-���u?eb�pdtPm&�����`e	$�Ch3�WG�y�B���tU�lմ��XD�F:�	���j��w��*�
i"��K�f��r���7�+��4�y�%\4=C��\0_���������
�@W���Z���ɚ���C!�w�q�`P�H�aV2���@�L1cQU{�4�*��8^R��w��r����Y���ۦ	O0�*rs�6��������IوiX�NKss�Ï>�x՚�ŋo��ί~�����
��kץ�37|�y����h<�ld��zzkwW\�LzF�%]U`�ތGb��2ӳ�76,:a�r5;:;�q%R;@[p���&(JG(D������J�~|=/K�p�tO��QA��lÿ[X�J�ߣE�p�t��H�`������Ըt��d2	�Цtuϛ�����^}�Ӭ;n+ m��_�8S���doo�\��w�^0d[��8v;���z��c;�C��d����hِ�dc쬓�p2{�OJ�LY�|f�g�p]w_+8��Y*��l>}�PIgs�b����.��^�������C��'�3���d�``jf*k1G��/�f�V�0�ɧ��%�������]r���dS?9����84�k`OOw�#G���o�Aq��R�&U��.�����s��dl���� �U�t�j!W-B�ĺ[��~�U���b�X�R�-��9�g �/�PH`�u��� �sdttxt|�[Pʦ}��lذ�^�Ő$.r�k���i���4{f��H(��bU�=^�a<��y�:6O�K��l�<0c<Į�1�́7Y�7]p�ũT3��'�S��=cn����q\��QC�gh\��T�17���g�q�oo� MSD�o�DTS�t���@��,��D׌h3��&�.Id�e�&z�U�K���$p��6���,B��aR���!� i��'/0�����r�ѰE�	��:B�8��r��~�����g�u�#�<�g`����ù��w�kxxh��g%ITU�������V˕���?}��|�X���5��BSSTY�E>������SC�B���;`M#K66;�'ש���Hg�f��Fqd�`�q�K��N՟�i� .���H|X�<BP����#��L�s�=�C���.p
��#��+�_dz��>�~�:�0���������"����sy��=������� C@���AUU,G��¼��/[�����i�&�j9��
Y��e����$*��I�[�b6[$2�643��,^�֜iZ�]]V�7;��N��OM�]�mY֍���wzy������V���mJ<#�!�;LF�������:��d����=���ܺ�����%���{��'a�ɪ~Λ��D>_ʷ����,/����Ffnn�r�,�$4�q���f]��Ƙ�����[�P�*��djpnΫjV������&t�� b��e8<�zy�阰������W�Vur"��XD�ܘ:qc���� ��<�#���Ϲ�e1.��{W��i�Ҋ����b�H�P��N�����U�J"-e� �M�=&�%���8p���GP�����lXM�^'�+��6�0(�����*�"b���A�`	�~�9�0n�[T/h�u�6/
�iĢ1�d�f���Z�����oq��O�IS�-g�q٥���䓑` �����9�L�e�]�rE&��{��W��r�Rش�/;:���#���'��c1^��23�_33c�
����' ��d�B,"�7�8L�ӆ˲�쇳���`�0��5��?��,�s6��
��GGǢ���+�g���<(�1W�_[�,�k�B��[/�����СCc��/��3����s�+	�TQ��?����<>�h�l_�����û�z�+˃�-g�GpL�w���s�'}|k<���)������N��T+�PP��*���ʊ=V(*�?��:���H���U�K�GÑD$�EB�+*-�	��hV���48E,#���V�\���ln.��k���,2���/U�
��g�=�z�����tKG���XCc����Weك�w��� �kvpd���H4���`zzvS4��u��د�,I2M�sn��,(6K;u�f�)�Ժ����}��V�\���s���b����R�gkD�A�e���	����#�H$b攚i��U��������WǄ���Z0 �����tztt2m3`P�oӡ%���k�����;$x�!+���$(����9�byKQ4���9G7�1�R7C�[mP��^D�K����(���+����9I�xC׽^�{Y��IU^q�駑����l(��������#�3��|bOg����|q<�t.�����b��
� � ������+�!�r"�_���bART� �M�2��"Xà�1�k�2Ȳ�:����@w����繵�e��� G��/���/�]�6����vv�l�ܻw�#�<¸�6��1��c�Ѿ&=Y�	2�����
;;;S��UY�����Y�\:EV�6I%��a�OU1Y�������G*�>9�nim�r��^�%�-�Bx�3�xIa��y��ƇG�A
�=�➇�{W��xJO__Ood��Tu����ڜ?N6�7�>fV��IK-%�:Z�w�tZ���Es�,�@��Ta��$˦ɰ.�jU�4Œ��T:�ˏo۾#a?t�p���"˻v�ilj,���=�;_�k��_�r2Ѱc�.Y��m���:���	C��w�����?����s��q8U�%�?�k�g?����;4�GD��h���3��ջ}H �5���V��5,G�� s���I˖u+Jz||�t,y��\.��#��m�2C�'4B(G)D1�|�q	[p-�����l에ڿ1�qE����[mg��Ϣ+�[fU-{$���$��a$�Ǩ�԰��w�SseHՇ%�\$�
\+� 闧�pG�e����\�r;�A���AĴGo�`OJ��l�(c]�A�֖�(*��bd����3����<p I�s��Q��r�j�Y��Y�L�g��0k���0xq�`옆�	͍͠�<�PcR6;GB4��s�����9XU4���&���`^~�!�R�a0�s�<kbW�H��X���0U�L4��մ	V�tf<_�F���r���(��>#3��,�s��D�R���Ly�����m�ߦ*��Stt��bT�l�U`���GQw��R��܋�1��ǆ��%I��O�lٲJ�:11�J��ɤ��khh0��;,��zx[�%��j�r5��l�^�������|KV�n��O����o9eŢ�'��R�9/��w�w]r�hz���]�����]e�?~����:�O�I�$�Bh��4wUDWv��]��.�������
vE@��@(�'������N���{�9��y�sg&4��o�5��a����s�������g��\|9+ŏ�z�]+W,�|���˻�P�����d,W��d[gC>W�moimimK�]�E��m554�= FÑX8B?#���g2L$���F'�R���:G�x!���o��'���e4gI�$���H"LHpy��
��
~�d�M�шq)�=������6qu	)�0��J����'j,A^],͔��H��pG>q"�B���5��L�-�Ѡ�@�"��ec��N�'q��ޞA:��8��$V��0�Mc�Z3�'BR/�OMeg��pxj*W�2�d�Lvp��`�C��rͶ�L�6�)=�S��|�,���n0�0�~?>9nZL��FBT^�LA�D[�e9_#��0�C�$C�|��·� ����rUrښ�B)�HAk��v��S�zq7�D���#�ӶPw��3�#��iV*�b�1 �E��h��-x&��ںO�|�/���tT	ϣ��!�s�E�$9 )�c|_H �9�,�r	�C�"����p%�]:�ı"):!h>}��gy��]ӅB",�'=!�1�JU˴t�
���C���3�GHދ��~���DH���}lhh�ZUGFFR�TgG�}����;�-�����b_��Nv;v��h4��ӽm�6��t[�X5c!�F]x�nЄ����� ��sS�0����=�Vkc����tC�d�`jY���ꆩ�^��W^�s3��e�W�Z�N瘳�/0��-A����G�=����c�yl7/*��`��>g�����1�I7��J��%�+�?��7[��w�6|��TfG{o�$:@o����&K7���#�o.+<�M6\���8A`�?"�NPʔҩ�l��a���le�!p���Iû��8��j�b�&��H�!�di�}q&	���@�\��!��44t��L�a���/�p����$\)�t5�X8H% ���L&eCrM|���I!���!W�`r�d'��m�(	�'n��M�#<�uB[�N0��'�!��b�884p���`��I������Fѝ��)�@�/Dk&O�1�0��BC��#����q-�m.���1D2��d)�5�����tM7%I�G�d���i�$��%<U�{�W�KC�g�� �cȎU��mWⅹ�����|�w)��b]��d�B8� �<�#�Udea,� �KD���$�}R4;qc˃�e���Nm�ɒk1���j$�b���ƈ�隮�y�9΁Y�1�#�z!��MȂ��`-�(�3��g��9	�Gioo�[�hժ���=���4=�W���ȏع����=������o�_���doo/8BӲ��ʊ��ÑH.����Z�f�����.aZE�f2K�c�����k���o~
�����}�E���C��O=��xv���d4r�[_�(�P�M�k�m�M#2�O�b�3ʰ*EK��rv���p"qζ����������|绗.]���G�\$,�{��u�=w5uv��9z��&�ͥrN	�c��'�2&G:[:�p��fu�#W6����e�!��$y�N���(�Q��GF��aU�t�	�K��X���E���'�l�8B	Ω��Z����Vy�b�C�%Z;�v)�^�!(/��	qƊJ�q���g��oi@	���+؆Y.�� ��J�@@�r"�Ww�Q��,�����Z�
�g,�u;�l�F����~˶B������;�=�Gxj����R긃Y{�<�cGy��D*����F6;R�9�+z��^do���2u�l;f[�"E�l �"�S�L�(M��BG,�:�q���#����x�s��ʞA�2�i@4Kw�������!��� ��syM7�����B8*���L�÷�Q��$�\*���QN�x�ٕ��m+�Hhr�s��0�����������}�R�IJ����o��_�z�H1�O������a�%P �ė~h�eQ���7���(���D2y��a��ǎ��[�z=����8I�mh��}Jp~���b�~��y�%�4
�f�ڵ�=�����<��e	�c���Ő]i��xْk;���0O<1U5�Wo]vd��{h��"*)����78�s��Z��b$bf2�{�=���>�w�e�8keb��X$l��x<�D2��K.8:�1��z����h[G:�
gR������l�c�_��dE���6�+����mτSd���3�ۡ�az�9��<����% ����v8����%�/ �<�.Û�%"s��[.��vHu^5��\b��!��!�����@��0�ϏA�M8�����A�m;ދ1��v
]T�k�qll$PA��\����E�o�axx��[~4�?R.���l9�Y�,��OY��6�?��k���r�v݇?U��d4ӈ�8�V�������I�2�Y/X��gO�3P����`,��+�����9p���o��c�m͍�cb}��3H�l�W���t���q�/�����1�l���~8��� �<��!0��I�kK���+�k��q�}?ܛ�Xd�vm�U�z�����Jk84�"����bY��0Y��<�c��;���'��ϭ[�V�xͰ��"&F>3��`�L^�gff�H�(":S
D�|(�S��,k���֝�8����p���7�=��˯��m���`s>Rb,�#g ᐞa����,�}N��</�0g!�BY�NOπ�NS��rub,[-�Kp-Ö'xX2�O�5gw��'~�n~��9�u��{y�x.��CSS���^�7��
�B��T�����9�W$�r�	4��I"�yׇ�8U2QIO�]S�g�3����-�illZ�|�����,�UGdHo�/_�/@�i�z�m�D&��)�d&�ɤd����F�[���!�N������������X��������޿?�%��u�Vpx�!������H�9���g�,X�B�\Ƕ��
����b��H$ i�
�hk�fl�TsI-r���&ɻxƛK�ie+�H�*@��ʁ����G .BH��j�زT�Uk5p~�+	��!(��g'&��)��	���X,M⼓My� F(�A��g�D�a�i����,���ᫀ��33�.�JRY�� �?�d9�_tх�)[���A;�y��L���f8�D�a0D#�#� ��t�߰^�h����b!����j�(�/AqJ���zًd5g,�PZ��I{"5���7_�K�u�ٯx�+�?x?$"d]�Q�lN�$���!Ǖe��TʓE���u�O��P�����r�<��LQb	�8N%Հ�6KH�X.U��\	nM�k��S`5"�D��5��:���RwN�A��G�ǂ4��<�ى�tУ�~>�8Q�1-�NW�c�\A�0��Ӆ�JMd���֝L[h��]]���]O_wݵ"��t����	�y�ĭWb}	��Ei��]�{������4������lٲGyī+mq�_t��C~r�k�C� 8�0��s���Tқ�Ѥ�9,��C��2_V�H䊿�����W�7lH%b���_��5�,_ж}��?��{V�\�w|p���^w!��8[������ǿ���/�[4�_�zeC&%p�m�c#�����������tS3+$"���@V�b3������d*��5�Y(t8,{:���m���{l�Z�b]��d�$���:-wu�TTհl��������6UՑ�B/�D��g��z^�ynQ�1��x��C�"����'>���Z�� b���/��қ���>�nl?<�}��;�sU��8ժ���ɒ��޲�x" �P2&$���>��Q0U^:���v]�2eY��RGNG���$�����ȅ��`jj
M�"d:���)\6\�E�F�v<��[Ω��#��o ��z�h�ѶQ���P��:��Sk�v!m ����}::�`�MO�����
�z>��S��k�h����ԣ��6�L@v�3H� q>N�� ��j5d�	��˕	�$m�H=F��2�K�:���@FS@�>|c0?p谨��3���Z�7M�2�f�}�����	���܆,d�s��`Q�~>oQ����&P�������/\��9���D�a�����_��^ww��] ��c��^����!&�H���ı� �>� 
����,Ky�%QJ�"���#�_��N@r�=������s)��dzn&����{>Q��5�ގj�P"��k���+V���P�=B���
8#��;�b��׼t�;���x���V�h	3b�9�/��U���%j��wab��U�Q�eF��T��#�n��w����&0�pW���2V)݀Q�S��3S�$�i5v���Q
�LS��M��H��갌�c��\�]~�%�p������y?�ɢ���3E�F�tB���x������}����ɜv��&1��w��̽�ݥ���L�Z�(>���������l�d��74v���}��'}��|�[�z��������&7>���^��s�e+.a%��2 y~Y�s)2LEg�9�J��F�5hݶ�LQ$@�����N��S��ø�d��\%44���.A���u���������C׻��mڴ���K;24����*CsW��5�S��Ͽp�[~���x��grS�-͎큧���|��������_��ў�����H��@Ω�[�M�\r�֧�Y"����e�7�9a��L�{������Z��7�HV"o{����j媏}�իW=����.�~���n����߻��[n���>�i�N��hI���	���,p��
sF�/��t'������h4�F�3����z�0�͛7�����8f�7|^�}�21>5Կ�o~�"�j�P��"g{�ć���X���~ǥt��>#�H�\�0>>���H&V�^���o^��a������vUU�ݳg|ll��U�H2¡�!��WˑJGD��!�����4=�0�w_�����B�h2w����=��$'''x����36�?o�yB��j���-�Y�t�;�����AϲjzEL�� �b,k�TS��i��+Woxd��c6�4�^��ٵ )�n�ʕ�n�����#d�D:d"�����G@�/�J9�}��="���t饗�!���9��W=����>��O�響DF�98	r4,a��p�N;��G�����$9VN�҃��5��l�r�C=�+�0�n��7��k:ۘrM�l<�k!gj|
�;H儢D4;�h�CI���˘(eO�9�a|��.�FV#|P����h�
�|a��v/�R��������9������<D��G�f��Xv��� �ܩ���zY�ר{A�1��~�s�aa�>r~�k��E|Ī����� �	$^�_ C�K#K��4d%5G��D�gc�œ�<f,37�6[�<�z,�@=����fK�3�D�2xY���6��ǿ��X�F��߹}����w\��{�tu�~��A�������o�lsc��X���d+i<���^`����XD���>G'�x5�c�F�� X�6��2�|n*�̨�=-��<ޘ����z�?[��E�+�;,�3"X�-�"k:�+�~;�j��yV�S��8�<�s`HE�j-ўy~.��G0*p�{��C��s:�Z��oAw��� �D����ZE�	To�R��e(���-'���'^H�]/�����t��J���Ҋ޳��d2s���P��N@�����E��Ē
��:?��/�������p(��G�y���j���{^��������o��nO7'�i����>>2�.M̅���׿�����-�{�9�X�dg���g��3թ���M͙d&uF�LY
ɢd�4Qq
�eDث��pU^�J����c�Wm;o�g>��3s<��b@�TQ5�Mo�;��[����� a�ikW����G��E�d�e\S�x�e������Y�ѩ>�V�u�5ONVM�(�T�P:ɔř\ֱ\����~���y]Tb��Z��e�[�X. sd�Dpԁ��4gQy�v�F�I�-L�Ba��J�,��>���N��M�>gְ�ZM�u��pf<��5P�y� C>���Lo�a�*j5���3	.�\)W!~qL��ɠH]��lW��kBМr����!� }�"�u ��~���=���������L��ZJ��y�_���>�C��5K5�����8x2+	��Z�(�Uw���vu���#ǆ�>��{����5g(���Պ��R<�Gth`��;	n��<�_��lہ(^-;��t�,�p�ҵƦ���ه��.�a�5ݨ��Z��t���k���%g��]����Y�m$0��sʉ�7~��#�1
����8���}���A�r,�������T*p�!���/~��Ո��)Ⱥ�����7o�$�����E��������0�]Z��h��:�=�x�864���=����ೞ}V�®�>r�u�z��Lk�]�n���{x��q�D:�I��T��i��={?��O�cR���O?�f��㣋z�)�<������۽lɲ,o0��z��=0E�Ӳ��zP1
LI_�</r�����ʥ}�[e�%|�A�66�z{;�ێ��O� J��x�0m�3{���C$v��H@�g&�x������''�.|�y�$w���^�D�j�$$���9�G��[GB"G�v8�ʓ�V�M�5E�gNhh-������q��#�	�'���z��<����Of�E�"�x�H���!�oOP3%�P"�B�C�,�2Bdy=��Z'��y��,� 	�M^p�#o�G0GcO�}
��� �?�9�w��}���?&���h؋�C�"!��B%�D��(�!��2�^�b���l_�b�s��pX���|9��5�2N[������xS�T!��")Q���b��$I���;R��-ӌ#�h�s_�RHGw?������2�q��\,i�Z�P*��;�8�y�X�g������g76����c�0��Y�=�X>6�����j�611>=9�մ�q��h8��ܒ��t	��{9�ng�e���u��@��_|1��lv1_b�u�����I���q��|sc$�ĝ�L(�=6l&d�>{��˿��oB���s��g�vsS�Χ�\�vck��/v>�Ě�ް��Cd̩�0�Ҹ���Z�E�G#k�Z�tp�9�z��~����ͼB|ks�	!Gl�rgA�bp.xL����>�/�G����lwWoww�m����kDca��}�%�9ug��4A}*Q�-;`�U& �z����jM}��g�Y�z9�����7nmW�m΅�N&~9�>�ӥ3ɸp���R���L8�x�(����F=����z�[�.�_�''�M�,�j�P��B:��;�q�t�,Kf|Y����+�inj����¶c{8i���)Gxj�iKDEQ���6��%�s4QoD�0w�tIƁ�� �w�{�زD52�kckб�G蠒xTV��uB�X�pZ[Z��G�a�*tH��|8y3�)�&�`׭[w�g�n���Dp�npM6SSkyǭ�S�.<�����W���PG�s�S��M��f�I,��`�M�3�0�P@��hC���d,�C@����[�B1
ڦ�H�J�R������H8��"1l�E��p(\U�p�	����U�8�9y�e�2��Ο,�����XRXH�:��3��?�2a��s]�9J�y�;�j��-ô����]xU��Gĩ5˂Ԑ'��'d�Q����>(䦛�R͍����G˖��ğz�E3)FU�����\tѫ��-�[�o|�3�� �2��S�D��K/���o�����g򹞾���և�q�kG��:�*$��p(�ڮ��"��r@�Vt�A�\3�P��a�P��l��8<�ڦ���B�őA�(���X,�ڵ����X���-%wÆC�(A�R^��8�{|_�r�Z�]U�HT^�vY�4Y(֮[��W�Z��j�[�pѢX[�� �5���G��"(�D®�}GcQO$:�t����~9�Ɲ����Ϥ��CpO�eY9�ư�� �ա�5�9�L�|�I���o�?,y����x2� D�}�m���O�Y/5(��M��A۴i�C=��㉘�VFFF��E�%�m̤`�j��������+K�}9�d>ݡ��̹�+=��F_��g��CY ���K�j-J@�3�\(��Q�"	9�k���;�9��ĥ� .[��oղ�|�[W_}5��l:��ڕڽk����U{��y�?}v|<�-7�A��,�K�Qv��!��޶o_1���'����jet�~>�â^*�'
f'����s�����]�z��	^��)�AСm�P�ʲl�=<�zs�����I9�D�J��>=�EGW��H�Y!��1e�F�F�2M�j{v?3:8Oć��u����h]ԛ34����%����bp����.��׿���+m��f'!okkk��0|�>��9�TO�m6�ZH��q�[�������u�=cӖO~�:�������Mi�b^�����o�yǽ\�-�JA�H$��@Z���N5d6�}�Ę�=��i}S�?�ُ�����Q�&)�P�6�J����=�`�?��%�֡���-����_�y�ԾۛC������x�ŋ��޵��k��\C�#+�b�!vY��w��Ax�SS3��D)��:W(��e�S���b��u�>Nܕ�Q��!��W^:���.Ja8:瞻~ٙZ��?��c�<�6Z�Y	����&0afz� j���G��ib	�-i4���9L)^�C�n5U��Aw�KЩ�KaB�� )�+�2�7�%�qY*J	5�dQ����%�vT��X"�����z�	�^sJ���z�5�1��4M�����}�����H�\GHb4e�x�s�TT2���f��Q�=Ne��s��-!DX��K<� $5}�&y�Q@��<����i�����8V�@J
*����Pd}�S�gb��B���Ȟ���V���W-���\�[��ϰk��z�#��斿{�U��zܣSYXUe	�!
�*"&�n�`	��ԍlv���M�K�#���E�X!��.k������\�������=M$u�)���ϻ��[�4��p�/Ǹ�xA�(J@�1��kB
���
�"�ִ�a��]u	rҲ��Z�T!���V*������em��q�r�/�6��k�o���>�@���Hoo/D!�m$�I�:b9�#�^/2�BI�ω�C�m,�m���X�2P�j�d�S���K�3�����ѱa��c\�ca��|�T�R�izI�^�|��sp�!B1'�b dDˑ�T�F�[��jo��e)I����L�B�	���e�\:xd�X���E��W�M�8�rOw��o�2�jhil�s��<�%�7H+�p	r�!5�y]�b��Da�j�\y�[ܟAĻ��u^�8���T,a6DM��="JX�h���`!�[�^Њ��J�,9�Rsk��hnj"��c:339MU�: �v�3<�����H��б	0ʥ3�Ū����5�.�Cd�L�����S�������yuvv�����"R�Zւ���'���a�[ب��ve�-P�p�9e�M�� ��j��62�3N2����p8
K�6a�wi>Dm��,]�B-W��H�'�.��M��~Ϝ#D�<�e0�$�ĵkה��P4T��8���k�����:24�D�J��Y�w���,k2���H=l�"��p�N�- �>r����/�8
� :2��p6�
�l�E]xᅩ����{ W�,����L҇�y��Bn��Eӯ(��(�(�g'Y��NB�Ğz�@"��*�eQa�PsB�T5��ý/�j�ʀhk퀼!��)"�?�y)���@������mii��i�0��y��+R��T\�Hh�R��D8�JL�EMu�Qn��%w��������nj��O�_��/bM���ad(�N��&�S�V�9\�MMf��3S𠫆!s�rM�,HD`�U�v����Aebrڐ��U��Z�53O%b1Y������ ΀Gz���G�}@7mޔ��ӵW�`	' @�q�{$�#�}������f\
L!�� �=WB�4��O9���Y
c���KJ`�鑆 ��8�AHh���&��{iZ����op������,���Gb�Y����
��L�"]R�9B�*#.7�^�+98z�G��,)����9q{�T	���"k�S���DCA�2��ROO������(a��h��1c����ClG����qcC������G�6��p�Q\	�E��W�N!+�|�x�����,Hkv?����Ba�eD,��2,b?7KL.W7�r�X,��mH	�ҁX8�"{�7Sқ2�4���p�t�g��ܞ_G��e�/@([��۞�U�Q9�I�# c��αzC*޷���N�#,��O� ?W&S����)�ζ	I�&���LLM�;p�_��]��[���Ɩ��z��M6mX����L
z�r��P�R81����_�[�:�)�Ղ?�e�����_���K��X��3���],��T:v=�4L$8�P@	+|M7=�֫IF��J�X�������|�#-�-S��7��M[�قw��_N�ť�Z��kO?��w~������ԅ�N�f�p��~��G����^(��Ԗִ$q��%���������ծlM\�r��[��麭g�XCS"�mY�8��]�S�z/�
pb�mCc#S�}���+G����߾얿y^<���t䵏^d&�vt��I~��`��X���<�m�D:&�8H���tԞ�Jy`;v�@�P�Ӳ�t��/ɠ<5f�<i<�����M����S� ��p�x��4��`!�/f�.C|aU��3�Qg�!��4yD��X��E�1�*Id�����y�?���_�N9Z'�7&�9GU_��x�V-�|l||t``�!���ΙUu�c�P�m�cB��8"p�$8�5�ƹ��X���U�
--���H8理��3'�E�� ��lX��MgD"���C�!%xh� =��Q,�����$�ٳ/�H6��Y���}��ꐫ)�0Q�!IB�h� j5�Vv����xN;:0��m�6�a��������t,�/��޳yb" 4�V��eC�@@	%I�uS�!�2�ᣓFM7�5��C�8� �(NO�!�YJ*�ӉL:�Iγ{��ʶ�w��'v����Ǧ������<sg�f���H�wu�Z� J�-c�T sU,��B!���e0��p��C�3�����:95��Y,1���s���욘G:u^�'� <�Y$G���>�8�q'3k8��8� �>���F,F�����}���0V��q,Z���\��m"� D<����^c�-|�74&�,+�xd��DH:�[��>|p����<t?��Zgzz7o6Fk��?9m��E���온[�V��0Å
\���{ǎ,\� �khp(���޿��
���02�C>����'��r����֞�Y��A֟����̬$}�����Ή�4�Ǉ�-j�����}%�j��j5�]˶�r6�@
4OǢ��FR �g�-{Ԓ�(�lo]�H@p�A�h�4����;Z� �y�����816�|�d�
~�`a�"���J��LS��ޡ�c�Tzz:��,%�8k�pypi����dZ����_V�d�r�/{y��0��#n��v����Oטi�iX�I��
����աeԗUk&l�pHH$cd��u8F󜊬+�D2��H�\���h5����S�2A�T�d�N�Ɩ�X���~��������HBG��$���ڜ�b�f:�D��k���D�I"r��p(G�(�����MM�Y$51`m2؎Q��^����|rl^��j�YR���Y�3-�f�I�Pc�&kX&ǉU���Ő"�z�V����K�����(7K)J�蹻?�`|���R�M��b���ѕ�6���w�k_
�j�P�8>�^E	�\� �8o�y��z{{3�LGGWCCӎG'��� �O���k�^�?y��(A<���/�0�<�����ᮮN�ta����^] �y/N�L��h~�3����!<��!nY��C�]L3p�j����"R�ΥW�m�t¬����(���]%�
*��꺦GP[B@�xn|t�1�<�p��l[[�$�8>8V�K��q$y"��-^��05ʜ��xD�����7�x2��)�a���!�/T���3/=�K�p=w[��) �Y��L�(�u\��l*��\̀XB��%<O.�UX����icS��}0'g"�(�D�� =2'T�V� ��5�(���x����@���B����Cj!�}M�0�GI2f��T"!(|�6$C#�ã3��hU�b@!=܊r���:����ѡ\v�LJGt�v��Q0@��͐EA>��ɳ)�L���q�Ud=2\�&A�W�VSBD������6���BzSK���X,�_�7��C�J�$��a��gv�.�pl,��&�/d��ci��H,����J���N�(j�9�	D\l�f(�`SC�#���z�����9��58���ӓ��H"%Qy�`��q$U�
�R[)���?'3J0e�3�����M���T8�;�v��Qu����ah�X�!�ί�:� K�W����o�{�#C��k?�����{ߌ�S��ۙ}!#�M��|���G�Ǟ���+�r�[n����8>2b>�8��I�Ϻ��x	����g�-����=�L.\طl��\����f@���6q'���6C
��L�b8Y���ti��%
}��X�ۚj�TSe쯣9,8B��`����
$��'�a�a��kZ"�M�,䲂	J`�#5;�*��Iy\�R�������4l���L"�hmh�B��k��s>�G�IG�ka��|7�O�#x%c|"l��$z`a���+w�W$/�u �Ç�S��N�tQ�D6'X�[�j�{2�j.���9�(���r��M�����R��u\x���3���gQͅ�\�ټi����9����r��$�t:ML�E1���
����%��r�t����S��'��bA�>�Ջ,9�º�M6�o^���[/U�%011�{ϳ��ҩ�G?��J�t�ȡ;~u;�^�F��`�6	�_�|�֭[��?��C��ǧX&�+k*S�r���=V���J�AQ{�@kX��K� �����-Z���o|��N$S���iګ q2o{^"�jnk�ҍk�r��]&�����.B�qM��$�(M�΄W@��'T$�	R0 ��C�T�Yط�W��۷�!P �U�D�U�F���d'�PH�e�8¦֞��.y��f xJ�
�貦`�����2�>�ť�`$���I�P(�����T�o}���#�/8kKߒ���X�Qm�����CI&���Qi��:vl���y����#���5�,4��t+�w����BF��u��a:�>p����$d��IT�684
��,�J Bx8Qʒ�@2��c��3��<	l��S�%�S)�B��c�TN�l[�k�&Zn"F�؞(����9�s���K8#C�L��"�g�xu\�c����V�0�j�������xtG߂��V�lkl\�b���7������*�� �˟X
����<|RW�s$�x�u,�"�՟ 3��&�`S��e�7A$�c,ťEYqL��,��ǅ?sL�@8^�����C��O�z�z)2��ţG5QM���c���^� j�u��m�wDۏ�xBY�Z�-��sp{�RR8$ATLN�E"�|�#���`d����O�E D@����fH�}^}�4��8ul�_��ʟk�r�'�����s~��T)[�j���˗/omn:z�(8B��r�(��}��^}|��+�|�ۮ���F��|a"�R3�\O�T+���G<.1��œ]��ղ��mϲ�$o(Y�riv"���mB�d���9δ�.*ù�*�L"��e�Qy۵��' &Nb���'a֩
��b32O8����mh v���Tk��̟�ys��iddɗ�z,\W���	�vu.(+�m��8$�b�8#�J�#|����˫Wo��:�ߐ��:+G ��ɆV۲�J�����#�s�9���{ۛ$�1&#����Y=]�
��K�.]�aî]�LO�V-_�|睿%�e�zͰ�~*s�H���ð/��m�;�<.�t����˳>�9�!��O?=�H��#�;6�X.�ږS*��+555ٮϠl��Aޖ��j�}��:<�u���_��z��2xqAy�j-�p�r�t1�,9��{a�c��;\$ISX	�9�f����SQ���?�����W�,wt�ߓ��[���oߵsWssӑ�G��w<p�����?��c�NΔ�����#����R��*E���=�� �����x$O�O�g����rΊ5A����<�����]����1$�Z�O&±��u=���3�޳#�-[�gy��J�RMTU��EI�%A��p��X��7$7�E�q�Q��������[�
y���y�V�]V�h��Kv6�9t���6��}�_t�e�,S�E�:��	��6m7�]�J)���\���g�b���єN�dY2MB���t(���`J~���$<�_�o�h ��>���-`%��Z�)CP*T�E����$`(�!���x�Z��"]'�):� �]�����2�;4�e���uXJFS�<��tn���9�8���b��\ג5���%2��Q]m8����9�Kx�u���d�͐3'W�58|�#��9��DkB�+�x�=>O��4���щlC*���6�S�O��WM�X�Is�Y|�A���pX!W�1xoG�Ӝ�ֳ��Pg����Ktɒ��h,̳�,�4��B�������������}JvM%����'��������2��3ETL$���o\�ld��㋗,��CI�	�jUSժ����p��F>�~�����݉L,>c���6l1tN`��HDB|E��HŨ�Pܗp�i��;�TA`�j��V$�*qVH�Jv�ZSC���uA��9==�U+V�?m�o~���t�5�����T�5ŀx��>8et.Z3>5m�ի�y��~�����H��O^���W��{$;������<�o�|8fv?]�ڿ���7��-�z�]��}��ܶm�a~n���m{�{_�O|�T�s�ݴ��+^��.+g��pi�VQUU�c[���w��0ã���(�ꏒHu�\�\�(�t.�ZSm���Χ�����766��j��#�eIІ�J%�%<4:R,��+���6�D�"'��s�(v��̩�"�C��@���v,�ĩ�r��s���rybta{�Y��~�G�d*�4;����@.e����tU�m/�Tڿ������N#Qv]<.�"J�V]��a|62��gN��#���\(dy�+D��D"��~�9'(I �	*+��l��sTO)-kCxF����
�3�-!d���h�鹃ÿ��dyb�	Ȅ���"'xN�r�1lwgW�Tz�߼��%�6��Nz��p7O�B�\�q�P�rM���]����5�9������=w���~�R,ʱ ��� ���u��L��NMAFZ�nͺ�����j!���s�0���RV,�GC�:�?R��'�1"d���6�������A��(ɝ�H�y�qA�aZ9N�_,�x&uQ���\g~Ʉ���q%���:uGln�y���_���d�nH	�媖+��j8"R\Ը��|��5�cҩ����p0���Dg[u���Lo߲�{/�bS(���� ���a�e�ƦSmG�Ƣi�dzт�O?:��O=;�eK��g��Mո@,ct�Y�r��\��J%��a���xǙ[�;tl�#�}��1��_���>rȝuIg�~�\�<��qs�ʛ�>���<��ѳ|����SG+Jj�Z�Tw<�(�/ݐr��
}
������:�P�ܷw��6B�]�i�,9.7�-�E�5,�d�?g����N9�|N�B�&8 ��D'y�B���O@:���pm�#�J�@������c�v��-
�Zu�q�T1�0YQ|����6(I�P"�x"�M~�K$��HD�j�,ˎ�y���l��fn�KeMIz� W��,!!&�%�����n��,N�L�
��)�x�2��o����G����Օ�Ok.C�:�w^�������H��$�ӹ�����ڵ����ʩ|�偣���sM�H<,�ZsRKբ̇�H �0~�Y�jՀ�~�ڵ�H�W���#3ԓ�hK�~� 8B��|.�����QB�>=BXFi��X�-\Իbժ��^]3�ux�	�����^֐���c��ϸ����喈&`G�n�2>��q�5�*ȵ�~FB��֚jik�l;��?�oh)�$x8��U�M�*�KhƢIð\�<11500��A��lTedr�����b�P*�Ӊ+W�|z��;�~�{���/�� ��ݗ^��gw�l8c��G�zA��v�Z��b��Ce��`K���H���L8µv�Jx�n�I��kV������QH�,K�lCfy�xQ� ��Q"=߈\�X���"Gn�������̆��6ᔟo1,��򆪁׃Z�e
8��  ��� ��57,2�O&�ڹ��	�䃱���4���01�G�)GxR�8` �z�''�Wp����/��ˑB�g��t�٤R}�W2�{5:�HF�jQ2,j��W
��"
���.����#�X��N��9$2#�Y��0��"�5-VR����P���j�/��!ı�s9��F[� $�P`�T�bI�#F9=�#W£(��!o��*����Y�Ecj�TBى���BM�$'(�����%�x"1<4�n����KR�d�p��D�G	��g::��	+��`�Z�%7���K$( Y']d����`������B�Î=�/��G>��h<y�o���%�~��M�p��7�Z1��<��k���F��P(204��>7*�l� �/�A�,bp#lp���^�?�E���}�?�\�ޫ���e�f��y����K�٩x,����d*�@�$��/^ی��q$��O������	B��Z\Abʺ�_q�T�[]D q�����X:�pP�X*�-_������V*���I�?�-=�@.(R6;��N4jk��c����eyaf�P4�pZ�p:����������
����\�����7�d"�f��m}���=�=Iegr�"�"D����.^ڻt�����gv��]W/_�����F�EK�p��b��_�����,L�cG���p�:�Y]���4ř}F��b>'���o��c0W��-�_t�x��ٖE�f�`�!E�y	���Y?I\�S���N�	�9 3�S�N�1Y�E\)�@��>����SgI��V�����hI���d�Nk*�0o�-����M�L�#p�SSS�V65�"B�\�$��S��$vI�y�����#��W���rB�Mtr�be��(�P�2u�k��@I�P��|�QP|!U"�?�?���K�� �/�#�Z�YK(�d2����܈��j9�M�����?D�?���j���;1������?�����i�BA�\�������;.L�6��~�UWU�j�5�}��<:ZSA�?g��E��j����7�xddlf&�q��g�}�=��ɻﺷ����C�m�D�Z��t�W{|�#;��}�E��r�&�1_�cc��P�xM��\Q�����^����[��Q嚫��o��81˴ |v-�@L\H(��c�8�j5=�il�h^�rlʤL>8�֑����uNƁ�M�1�5o����U4�8vl ޴��3�nlnj���4m�䵢(�D!�e,��HS���ujYN(�mN�#M[:���s�}S5�d�$�^}�r���o��wBJ�n��+�|á��>s��zՕ{{�;�yϱ��L���MH�tA����ݷOd�f�[�t墾��`ICc��3Ί�SE�{�3�Q'&;z{[�Թ�\�o!'LoW�׾�ծ�ni��z���K]t�Za��A%�h��w��˷��-��sWM�>���6`j�B��@��ࡈ"���{��RD�Vc�Z[S�M��"��J(���0S et,l,�[!����໽:I,7���fy�_��O�Ѭ�C�x�u]��Dw�@�F��
!��s�zЇ�a�N��x"	�,�Ġ��0-��)GxRkN�kΆ�֋��Dr�x2On��������{�~�;�E�R{���f����j��0nNq���mo��Pt8pH���bI'�6͙��V����������>�9�)��K��ʠH���3D
��W ����onZ�f�VH~z����+o���+�������k���w���,~���[;��߿���gϻ��t:����;�z"�N�\����7D"����xIX�rE4:60������g��di��?�a:_�r��WN���#��ފ ��h�p�q.���#1A�#�4��B([,�,�o�B@����Y���I����"����|��h4���3���mW
 ʟ!&_�d!�KM@�c�%f�{aJ@f'4���q�u�$k����m�7J���\���7c1n��OŎ�~�YgM���e|�صkdHX���s�=R�d<,�����3O==�����p�e]���L�(�V����Z�f'���Ŀ���Y�f��uk֮*�
p[�6%�Zw<s̵*���<f�Y�����p�9g
�rqwc"�v�2�dZ�q�T7�^���Gz�3ɰ\�+M���g�@`���W\�z�w7l�p٫_3x�<���?��봪��m�66����d@�H�	�1K� ��AۀN��Q:�`�Nt��Ș�;�n��O��9��j�(T�]�F:g?4]���8j4�LX�a�J���2&Q,m0MM-�:S+�u�B��K�j���T�_���^s��W��=S�xɲ�KV<���P]�|��lN��/�ʐrB��(3��*�'���؊�!���������o�!;1�eh<�;��T&�����і���mY����X�5�s�t�ĝ��s�M��7N$2�a��L�0N�y[ϋ%Ej����EC����S���'>�-C��-h�ַ�q��_������O����}�J`iߒ�w<��}�ۺu�.�%y�s{;:��=��qv<�(X��/{�gמ|��;{���E'tMgebhXKg�u��"����[�z���6��X��!U��O��r���K�h���ܜi��4�P &�J%��!���C#�ZE���d����c��t�m�|"�'X� ��hC&��c�b!��I�s�/���&"��JH�����I/����	[D�i�'D�BsS�%]r��-�}�\�P�3^�j�.��:��ǄP��������U�x3�#�-:m�y�T���ѵ��ݿ���+�xb�9F世�Ɗ���}Ȩ����t���2��'o����Gg��і���w�RBa.ܰu�B��eJEF������������û��z�����o.)Vʧ�mZ�wSXb�����{���AqQO���}.�R�,�[Ԑd��e�|�J��eKבCj0(�M�EH
��g�B�R7Aq�YG8���\a����2�w e*�r���s";����$&�p�b��u���u(�S/������yA�V �9�L$C���K:�$K�_�:�Oj�@����a����؀]�z��Tnbl(����39��*��/�َ��@�]*`\�3]Odx]�%�S>��J>0峟��C7��ɡ�/ǅpܐL�qL���P�'���N5�H�jY �$hm�'P{��E??e}FJ�y��;Í�g�$��b�86\�����DT3���~5���-X��c�c����ƍg������dSK/XjUE��������;MMC�(۵L�`�\�vu���A]ל����;0;�����8~B�C}!滎��[�9���O=��+_��\������KN[�ֶϱ$E`>N�G�u>x	�wL@FC�͛��4M�p5�h!@
+σ��D^���m���K`�p3�Y�E�������T4*�˩d�!6+�L�e���`0��s�i�I�N2��^S�D2?)���A�r�L&Y�a�$�_Me��������l�u������wQ�/k�vs�:� �WU�J瑶���%A�b"��wM��G�ԋ�?��X\�&�ܤ��Ö9����w���Wo��N&RG�w�q
�����w>�v�*/��p���K�����ꡐ�nh���9���ܒ����,��ɼS�c��������[Z[���[��\q��W�����bG���'>��'�}�;�O�M��Ǯ�@:,�E#̸������ށqT������E+iU�d[r7�w0`�iI ��B	�7�J7���7�������%�[]����y�ٕd��$�_�Aȫ-�3g�y������_���uf� ������Ux�P�
�:.Pz�54�.����l-78�z`|�Օ>��J������F�Ii��#�d�8�$oSZ�"L�$�@��	�[�b�<SjV!]F,V�X���Yjii	�`�q�B��4v͗��
���F�R.3����� I�a��̢m��R�#�`)xл����"�gG��(6Vdp��9]���YK#u5mǎ�����C�-��9�}{��_��A�12A�<a��f2��?�)���D����Ė�S���'ڤ�<�*r(S3�M��)���ǭ�*�:]n'�e,K(��c�$I="�g�l"'�.C�A�9p4�M�F�='���������3��<䍍��*�`u�BWg4����>�c�d2U�Uj*z%�������DTc*� c��Qv�p�Y8y��Sbw��
�b0\V3Uü���"��C�:eg��`y��7NS�Hl`xxpV���ʫ���X������c�X���`Y���
��M>1��N�|^�A�m	�B'@tHb!f�v&�����������Q�*j+�kkkG#�]�55U�\n��)�����=���� \6B���666����"�5k։��T*�xɒ��V�2X�����W\��7��ko�A&K�"x�P��y���[YY�A���,@�4���]H'yÔo��In�����c�S3��{�.,���lA�fw���4��ޛ�$�N�J{����m`�8�F*��Ƣ����p�DF��h�]V��������[��i�����⽫�ۼ��K���y���G��G���s��*�N�p����ۄ�� �1�+�Y�)�vk�I�=��(|��Z)
͒��"$C)�4X�g-pceQ��v�a$)ҌD������h�C��gO���:�8���t��M�8�f�iO�"K	�z���"9���֍��Ƀ%P����{}^��B�QdX�$��w�8���1�V���-q��]]hZv6S�}UVV��:�ڏ�r����1uR�0�o217>��nV^A7T�t%q��USS��"�6x�D�O91��#��DQ�.�vK�XO��#�[<Od��`�F���;A���_��d��2�����"�eo��mS���Z �z���o�<`�F�_s��^0yrhx�gd���
�ƍ����i����q�r1k�4��𽭭-u5pQ���6�X�C	�b�HA-�EVWWb�g[�=��#![�%2���TttX����J����+��楗^ٴ��CIF�E�p;]��ﯪ�$ˮх��;ܮi3��\�j�ރ�d�َ����և��+����{k�A�;��K��Z��.{a�Kpb7���OȒcڴ�mm-��V�^�k�P��7�onn�ӿ��~���~�{.z��G�����>�7y�9x� x�+W�<z�(܂�������1eJ��#�F�"���^�h��Pܴ��������aHĂ�.�>k��?���^��O�[9�Dώ��"��]�ԏ�����L�S|�T�xkKu�tS7&5L%X^SVQ[V^%�r������Fw���3�୨��40�TS���=������_}}��=�tf���;��d$���s �ۯl{sێ����Ӧ{�Ϗ���y�c׿�����_>��~�0X8����bV�b��'lN�)>5)K˶&���<�S�˽E�-S�jKK��,�:vߦ
�	�y,
G������j ��K���'	n�a:_�~<N��/
��,�}
:�`�����c_�A)�����[/9�%�f��c��Uߵ�"�gi���l L0�L�,X6�)&��W�0�q<b��=�r���(��Ҷ+�`^��$�4-8.rV	��4"�	y#Gs���#��H�����s!����~N���\^��)�ۢѨ�3������:p�Po�Дi��A�����d\�Ew56�c�G@���T\vŕ��E�O�@������c�,+S.ڴ�swܲoO��E��2ݻwסC>w�ݳg-x�g_|�y�q���u��{�%K��E��B3�
�D:3��"��m��nX��g��)֢��pi\ �zO���z�c����5��2k�ȧ�Ƀ-G/�|>���l��*X[��l�������I"/�Q���c�\��K.����Α���M��\x��eK~��{�ϟ�iӦ���ڪ�O�f��3g̸���;;:A�|���~��ׯ_�u�xk���ʪ�/��Fҍ7����g�om���_��K�^�h�-������鍊n�P� ���J8�����~�p��ǏÝ��̓C�]=�y�/���e9�I�
�����A�!_����!OV��U}ꩧ.��
̌
�I��b��U������p���m	�������1���N����C����u��!_�>z��	�u�}�Qp�Ea#�Y�,��L'�CU5�bX����g���o���o~�z�񺙙3g.[�,����s�F��}�������/�sΆ���U��ȁb�#GX1?���I�&�Z$3�3�!p�aO�wiH��M����qp�����5u�/ҿ����j @�)"r�Q��bO9�CtR-H|8��O�4��� �A* "��R���<G@�'z�0�t(��@Bd��C���0 	��w;� ��L.c�O���$K�'U|���v�Q��аO��(�-�,J�qN�8w���r�p,:�d��EJD�n���0�c��ԧ ��dZ7Y�H~�ǂl|3��[�����!�z�gm��
�8�pՒZ��^#�Xؿo�3I
uM�����������\*av��y5�f{���.��9��	���;e�f�E��Q���ۺu�囯]�V��7��[ U�b�R�aኪ뮻�O���=�����'?����狷�q����fj \~��)�;_�7��$b���
�U_���~�:�/ �{�y��,e�(:8�̠M�,3�����������N�F��cǎv��p�i�$R>��4E�3��[��:/��"p�њF7�=���}��v��3uJx�̰�#���.��M�\õׇ+�k��睳���'Ղ	�[__�q㹒��ֆ׭Y���+����F�U���olj��`���ȤI�jjj2�Ȳ�˗�U���j�*�wpʔ)�Xd\�2\^�T���3t�|��^o�(:EXGWU�e�Ѯ�n�FN��$�^��i���L"�\�|9���>��\���p|����N6ki͋S�"��w4��+��,<C ��,i�LEfo��&X�z�)��9���n��P2�a�8x��ٱ�t]�2�z�o��ZX�ɤ�#��A�KN�����<O�۝�d$���r 9Wlf�Dg�kg��{wl{�Ԗl}��[?{}lppڔ�W�}uά�s��
ych8�A�GgiNY��N��\O���򅪪0����He�t����I|��e�6&��Ȝ)*17������qh9	�#�`�9S2H��e�qX<�&q���o��I�-�n�܄B�-��8� �E�/�`'/�F�]>�����r���JB�#��C�_ⷂ����R�<������x,9�Nol�?����W��\͕J��7K�?j�Q��x;��UvE03lSbMKw���+S^�G��%�k���؆������$
�i]�i#�`S����ah�2h8؊"��p�xD0�~쟵��3��D��I��-0k��+M$�dE���t���S[�����9eG���ݩY!{���1�'��,"]	���W�8���h���Ͽ�FZ�0hE�t=3nS}�͜M��m��aOh��n��c�G3f�t���Md���;g=�,0�$X���Oɤ�/y�db�z{�?Wt��!OZ���R�}�*�^�z9!�I.��ЭT<Y���] �s$�8x�`uu5�38�IQ�q���l8?�J�VF�
�\�s݀�4�.GMM���3f6���A?\��T-?��**C�gm]����,��8��A�)���"?𠦦��9� �SQQ��h_WW2\gx��v���p�֯�$:Yp{��ɛV^73����q��_QZؓGݏdX +�-Y��>����b��,���0�E��U��K�`hyYv��4���X�l� ɝ]�tv��%������.ohqbž���='V�:MJ� 9��بe+?��O��mp��u�[��9g��g�Ի�օ��@�.�۸u�3��z\�����iuS?u��T���M_������z���:z!%��$������p�<x�!�o�؄�+*uӖ$����n�rf���E�|h<�>K o�Z�Đh�d�[Ƌ��X:F`�ip��+j�@�r`J�"'����Vy����d0�U���e3�T\۶�k�%���	�v2�����	�a�,�/E��o�mz��T"�kR}ݺ��_߶kxx(T� � ,0p�N˱��g�?4��u($(J��(�)A�dd2����j��r��Z���7��4]��"}ĨC�X�H�g7կX����ϽM�T`��b�#���ry��>�̧i�V�R�v�� �{�i�+�MZ�n��ԓȖP$쾾���(/S\N7'�ݩc�+v��$���R���ũiF����8=�3	�� 1<_(���ká��r��bw��Y���Yg�c��טɦ0���sf�`�J35C���@��}g��8���E�S�H������j��4�J���2T^��Z:�ʂ��x��Ӗ��&`�jk��&�6�룐E� ��{���S����u�S�`4����Be���Ç�a<"8\�L� ?N�k49�֒Φ�z;a.���>���sV6���:��Fc-�m��w��:\Αhd4=��K��v��᎞����{akss3(Ҏ����A��,+�����N��Q=�ZA%%� �'���M��t:�LGGGS�̑��7���"�e�#��	�Z�R{夨�ۼF��p�8��y��+}�'睽 �͑C�#��UK^~����s)U���K���z�ŭ+V�EQ��pT���ͽ7~�FIf~���7��<�u�P�+���\.+�����G����R+�y��֕I1n���?��eF�A����ql^� 杕��
t8�V��]k8��t{A��+�WQI7.�N�v'H
<lX�>�൙#G��
�
*h2��,p��� ����x���"��#	"�E`3��'ƙ������e�$�-����̈~�W^v��6]x�X�����b�p�A7��Cjh�̦|�;�fTW�tuޞΟ�O&�����T���g�;�}�v�ӐGx_#��C}`�͟��oX8^O��~����R�9�:F��.���O��m��}�vG"	5�l{&&�L�Ȍ8<4*����
���ϓ���B�F*��r?�Y�L(�?r̲��|B`��N3[=��%B<?P�,gKX5��Ԡ�/���r6� 
������LoD��Zްm�Ӊ���,�p4,�3J�'lK�#ey$�Y�F����G�y��Pj8D�]8�ENx�YL��&"��~��G>�S-T/�8MM3�r���}ڊ-JX�����k����p��t����e��pu���6F��U�k�dA�fҊӡ�M��� �I/Z�h��Up`���AK��A�� ;���J���CLH���@ \r������
2�U[S>LqC�(������,ӡ(����V�7�]�`���:\Qc1i�A/D7p���EUk�����\V;�֞�dA��L�2�7o�ÂF�	~[�N�-hs�I�pct�o�ш�Up
����o�tz}C#�����ɮvf盇[Z���p!ϴ�Y������G5-E}G*e>����m}�_�)�e~�������w��T�z�tZ�'������U[]��D�L�I��C �fj̣~�Bww��)�̙<���solX�
��=o��k����w�6k֬�AlD����MsG��݃��W�������C�����DMM}}],�5���G�;�y���55)����T-��ZS��
�x�A���ZQ��LЬ�I�K� Sz���ÄA���\� I��5���UU�^y��f`Q����P��6����%SzX���n7x����/]�a��d2#�rY�5�w�$�"���)9��oZ�_����0��a�& �l�l&kj��۔*����R�~%�%�J��l���i
wI�,)#�I� 6�,�uY�9�RLQ�Z3���4_O��H���ɘn�	��m���K����Nmk�T?	�v,��=�[6�j�ʇ+�F8'P��j����E�S"�K�H� �E҃��r��_��C��+!x"�T92�S���0kaJæu��`6�d�Z�o�����pAe<3��5몺Sێ�!TV���k���	HS�r��<u�������2��<��zttt8	� �@�ق'��>|8���
ee
\��={����|��O�3g�%1���>����jƌip�N��r��M�>�V.���4'���nllJ�r
j�pS��l,znΜy�L���2p��Nopz\�|~fS��pT�V����G"���t�3�>kA�&\8� ��h���}��u>����#Qx,�|>�s�oӦMn�7W�lJ�jc�!�)N"*'��x�K�DxR~̌�,�]�������:����]0��S�@WT��u�g?������D:��=���W�]���N�O/�v�t{�U��O���::U�I��ڏ�����O�\/�e>������2�.��;3�� p�&��pә�����]6m���_����?��O�׿y�������?��t3筩������{�_��O�kj������3��������I�y��mp5�ۺ�ڐ�=�o=q�DxZCC���|u钳F2iGֻf�J�٬ ��D
�)0c��Q�ɣ�LнdIo٪c��$�D�U�x��,���b%��K{K����O��|晧A�����Ra���(�~m����E�mm��[[7�wCp�Q���D0�M^��[�]2�(����l���x� ���ܱG-��˝�JPf�@st$�ȟ�������:gt�H�5�P]�W!���䜜$��%=,�S'U�ۡ�u�töL�+��ߍn3A���|���������A�F�eү��*ǉ��0�������"vF�ˊC-X�ޥ0(!���߮�LS/�+�l���*�&��,Q��]*䠿�k��მN���ܢρ�zG���s�v(P\��E���nrw����x��IaL#Y�L���#�,y!����t�{�=�/=w��h�9=TY14:Y�(��=�FPH`0�
?�!Q)9��� ����e��B~��r���c���ښ�jEq$��"�0D�\dl�s�M`d����qT�1�S�l,����Ď�oΟׄT��1p#�h"�Ow۶7n���&�yA,�d�w� ���5<�;��J����P���n����بC�c\[2��ٯ�:�K��޾�G����+�����ԩS{�#���̟/'S���hy�G�ܚ4 	`]b�4Kk���BG���_��I����5�e�v�/�핝��,��0��T�HL��+X竜̺*�Z$ǔ�̳��rW�+e���o�馛���mņs/�xE*�<��s���5kV�_=V�T����{|����u3��6bD�JQ��z�l�7�j}>�
��S������k��K.�L0���TIAb�0���7������� �XɄ�oĢ$�M�~2��'~�_�3������>V��W<�*�Q�̙�/�&P8|`K`�Y�|�g��/~3�I�YؗƑ�N̫�V!�v��GN��?�n� ��f@ej*�� BA@E�L�BA@�0�+��F��EE���ȤRĴ������`I��8GQ-p�Xc5�%��'b+��͇�M���^")������-C��O~�{��vsoú���T2�,-�'�'�&���Mfm7)q����q��h3v%x������{����{���D�C��������T�tZf�C(;#�wO��dJ�^?(b��==�e�I���e�w���kO_{�u���P�V��v�<�\NDUT��*��w�=��p8].���0x�C#x���/�E�D��兏#m��M�9��t��8 '�����"O����3.����§H1p#AD�߿?T^^_?%���92��}}}7�����ʑ�Iq2����|=K�uY�+C�i�&��kG0Ta��k���	Ü0x�W�M�G�/oS9.Ųy��P��"�n���n���^��ķ�m�{�e>�C�Ԭij�H(HX�r���$�ql��k9ۻ�X>�o<gu:�9�I��f-U�w�;���h�'��oR}���1ʼޑt�zr�N3�6u�P����gu�SƸ�eC�m=C#�C-m������]|��C�heu�]"�6���!���e�:�AŌ ��0�B�7�[S��&�w�m��de�"�E{�2�,��\�$�n�^a|�j��"ɯ_s�s�=Md�����LT��3���1�T�m���$I�>��w�_���w��n�^z�P�l+�'���al��XXφ��LjH��b�P�w�+Zj�)V7`��(�[@p�`ǋ�O2�_����)]gyt��E�F����=�����?������h��{>���[n8z����NM�ܗ��\?�K��y;�}�4�cx����i�b��d�;��H�\Ͽ��V�1�pp�L�w;���Z��&賤�p�΋�~���OI����ZCg"�H��`���7{NS(Ta����o.X��U7M�9����h����W�:;OUˢ�$�p��?�%�pe�R�T�n��Λ�5��C�2�ǟϩnHE>^ �fe��E����pI�CT"x��~��_q�$
h���V?L�-�����x�";�<���R١��Mn��'3銓῏�XȆV�\�l|�3[�4͙�vI�hI"��|�g,c��5�#ñ����I`�L���D��\�S�����8�ڲ|բK{$E�f�4tdj�R�SZ!ܴiSLC�&c=�mG�k������|���<������O���VQS�q�FXՆe�w���?�K�!�O����F����ʚZ�`�w��F�ߊ���=>w�2��ks�f����?��+�7>�]k�i��E���R�W ��A��I�+�����vÎҿ Éecz��aO��(}�pÎv:]p\x,�U�cJ;�n��HV�Yf2�����S��f�6(���Z����%<���(��N�i$,y��OX� �n��i����:�h�m{ U�((�sUL)�,D�:O��L��,�
ҋ��1�2/�z,�L��8
NG�>�n8>�{ږ�S(���Р[2��m>6g�Y��x�'���d8��˼� nO �t8��Nv�!.	�$�r�[���v�,|�'��_ګ���-g0cr�e	/^�R���~�v�pE�,�&^i|N��B 7@ȿ.7w�,V�b�����)���r�պa{}.���uw&�1�,�y�d
��(Χ�<Z����s��ɪeAo{g�,�?�,���Թ�!��x��iX�ո��\�(*�h|dd�Z8<�U�r>굋s���
pO2���������/M��x&S��.K�j�|+��:t(I��W�Rc�l�LAVf� �J���̛BMM�G�\
$_o�	����������W����S�����Z�6�����b�N��P�A|�bga)O�M���Hr:�(n睳�s�%�"C)�gE���7�5X0�b`:TT	7��>��c&.��V������Ni�Ċ���!��Ơ�M������ Q`��LDrw ��.Y���gQ�Y�il��e��P�5����C�o��R�b��z�yyN��ԟ���Ƕ���ɕ��l?��y���
��n��#G�7�ܽtيW^><���sg���ښz�G�a+V����P�</91�Ȋ�@��mB c�f$�i���E^�	���uR.�3C �^5Y��0P%�2�D�)�fH���|)cd�0�!/���OD��XQ���eF"�@�
�<�����^, 0I��]RHsF��F:�ܩ(�|�U����eZ�͏/!T�z��],���4b��P�M�Iԋ��f%y;�.�a�0"�Q��!�L`��2QdT]v��bk����q6ϱ�N,�ƶ�����'U#���[/^��'��,#q.OB>y���]�=-S����7��i�x��>ˎ�����C�cH8���m���q�=�<���f�_��r�0���'�{�׾z�C�7�vĢ�Aߗ��'��U���h=���}D���e�M��6��`$�B�^_ ��nT-[g������y�I�b�aI�^r�02�v˗/�>���X4�:��-�j[z�����?�͆���3��,ڵc��ū᰽��K��ɪC�H���t�b��"Zvmm=��X�E��$ӱ***M3 g�J�:�:����M4�ś��T���Q�H`�.*K�!c	d9cǺ�R������1Uf)�Rc#0N��:݌��k`)�a�y�]x��F�Ea8�i��ӴB$��H"�r�r>���aP��KB\�ڰ���"�H�Iu	̚%s^{���Դ���Z������\f$&}聟<��G�Z�?q����~�ٿ|�+��/:o]�����3|؄���ok
,>uix%y;�����P�o��,t��|A+��[�RB���1�ԙ/Y�4Qo�S[�J��b^��A��m��]>�(�w<���ĝ*V{Ж8��2e���S:��i�1��C�L����q��Kh�'�	�7�V�IJ��V/&�-�K]E�X{SDWa������$hK|�N�`O����%�|����Fl��ʩ���cWࣵuSZ[۞��������C������=NA���Je��DL9�Ts�7��<���#h0�]l��(4��N.�[��ǡ��;yB������7�۳k�������Y���7�m�w���7o~}mU��}�]����������v��=>�ןJ�#�����ʂ�K��@��gWT�@��F�n4p����i�n�h!!��ʰ��K��4G��ĳ��f��[�d�� � �S�`���F#+W�cY������P�ښ��|�J&�y5z�)K��N�<�t&�K2�W%���N�e�]]=�D�W_"ϴ�|N=�,f��坍��#<E�r�FC��&4�D�VtM(�PbC��&��#�	C&��p�N�0����c�cx��J�Rc���)eQ���B���`�XHvd�ɹe��[�����,,���C�t�'�����n����:�UMn��f�Z��,��YΤ���7}�YX���UT��N�Zv�q��X��Z��8��R��ȬK�@��d�ޔ9�V3��#�H,��*�!]�MM6%,�'��{1M��UU;pT]��!���Di��7�^2&imee����E=Ni\�t��fz���3���1-��"h����B���c��D2n[cQ��Nu��X���O^�À�6���U���^����6e��K��T8�#��$-G1�"�59:�:�m�H�v5��k��Ť�Y�˂���G+�-߰v���*����ZG�s~�áΞ�u+�0��*�>�Gh3����5��x��DX���w��풜�C�z���X��u��wl慟���Ġnh�jk���`5<��'�{�T���|,�����tOkhŉw��u����6�L��?�'D|�͋"��iE��Yۢ͑H��D���X�]l�{��t��)��@��W�^�������/�y�]�w�ߺu�%�7o�Xĸ�"K�S�@_(�7���|�<�7l�|4=z�e��u�5f���k�����H"�}Z�2�������t~�����#6��;wꬆ:����$�ёz�����ޚ��)Ջ�M�9I��,���6N?g��z���P�Lŕ˖
Ǌ��h�Vzp�p*��eaw���FJ晕gM�ۛJ%�V��l��/kz~J�c������[�`bf�&�דɅ3�T����Sf��Q��}��s�I�-�P�2D�DlLC�,]�$��%�~����h�6�*�'�X�4A�ґzN�.�m�2��J�'���ʫ�N��S�a[���Ȱ�!,o�C�nY<i���*�f��"|ǣ�X�YR�A<���Og��g�U���e�n�CU����M�Qq��� 1��'D�XSl��.�Ŏ[�$�1x �Ƃ�A�FDln��_@�B�'��Hd j�2E�_�	1zJ^���"9>{�g9NbM5���<�7�[�p4p�r�B�(S��R`�f����#.�M&��SWu\n�TAڋK�՞�|	���ԥ��t(N����cǎ�8k���ڻ�������f�|�ؗ��Ŗ�c~�kӦ���ȟ�rݵ���?XVY?��C�ƆxQ����f�;�,:�����U��9u�d�S�G��D� I�5V��hv"�J�
����x�Up;L���3p|��㥂j�X�����Q �����K��;~���'_��k��׿���7��H+h�-����E�DQ�%�p8Ƌ�l��C�Cp
��r2��\�����J)�J*ϲX�4�x�}�[�±Xk���>��%��Z>��I��gCr9�Q�/���?��-��Ƕ�\����n�s3������pfx$���-�#�{��m�?wnF-f��[�����3�N�!�:#�0�.uSGT$ȵ��bP����`ڱ]U�91�9�D|��̳�E�8�X�[�I�^���t��c�Y�ϥg���Sj*��(������%�s�eh���\85�$�DܘzAgJ �e��lإ
Q��-RzV�OX�&
����'�}.	Γ�ұ޼A]H&:���'��E>Q�	!ʿn ���T\,�VU�.��)5`�#w&o�'�cl��4��ۻD�Q��x�JL�	�Y��ĲTSY������<�E�l�p�@�.(����Ŵ����������5�v8X�~��ܲ��'��	�|1���W��Y����RJ2����x�F~0�y,f5yą�����qG��m�$�m���)��)���>�x��c��g�<���ˤ@U�+�>�l*wɫo���믞�l���V����u���W^������pт9/���0��Dű퍽�<��w����۷777;�?��fL��N�׮Y�p�\�ˇ��XzJӞx�T��K�avq�ADs6����J ][7i�^�_�?w��u���l�׭_8x�Ȟ=-�m�$��[��!�	Q"9��$�N��t������;������y����Y�&V˜Ǉ^����3����7ǡ���_o9�<u}k+`�<v������;�E�7wes|.�ag��H$�AQ��b��	b)��;��+���V�&	�`���gD`$H�&���&��zi&&$X�m�܄�j1�FLD,�A��cY4�����+��H�Iԃl�Z��k�)�����R8f0���z.��Ǡ	�%b���jƎ'I�X�-WJ�`��2HP��xz�l�M�\�M!�On	�i�hļk�E��M�� �|&B��O_{<?��Yn�@��Hb��� ����:A�8#��x��h��KJ�LڣO�n4�� �������.�8LBF/���BR�ɓ�hA�4���\h�� A|�#��F�&��	"�Ƅ�bؔ�ƍWa"d|ZN���Sʀ2��	6Vyü�I����Y�f[z�������)�_��<[�~��_���u�Ϟ;o�Ν��p���s�,X�;䜦r�ĩ�iА��r��������=�gϞ���G�Ã��6_r�W����ƈ��[C;�F�ș3�ϊ�����+&+����%�H�`$,3��QF�������/�u��᪩]������'��qp��c��@B�50ю/UՎ�yh2�!�^�"QM�~+9���-�\+V�%f��Hu�۫��$G־E;DYFq:F#/o;�ͅ��J���60ڽ������u�$T�r�,�[b(��É�Nur���/�.k��
��\C�7��'��l)5K�^�q��X�2� `K�K�,;>{T�Q�9:�nK:'��4�ƶT����`!1����/��?6o��[b�1�^(1��z\nЅ�T��r��h�m�c��^2������"/2x�� `�a�?cʢ �x,�3����%܇�rS���D�G�����g�2��ElO�.�kp�?��²�\:ŕ9ݢ"v�Pm�B�A��an���i���鄀��Z�0 A¶i� �IlB�bY���NmR��0�b��4$�`�8xR�M�Q	*!X�v����W�AVs&�y,��جMҖ��T�Fr�c1̄+�ߚӊ� %�{Ҭ��H2�8��y�8�\�����w�|�����9�����G<��Ν3�����jOW��V� �((f�*��UK���o��W�������]�������'4̘Y]U�8]��AA<HH�2ލ��堏�"D-uňЄYFf.<{��0'��}�>v�'��Ǉ���+6��-W�wS*��{6_��T�*H}D�I,��%�D"�Ln�?�K�a��(�1KĊŧy�����QX�
L
4��d5G�lm:�o��	~�i��O.b���v��>�vyDgM2�msn��"���28�4�7�F( ��z"_H�E~2o
٬�t��M��f�,�D"��K�Ģ*�6~Pc�x�S��)�T��K'd�ހ��E�$��IQ�m�LP�p(55f�T�2��� GQm.
��4T0K�����m��2��kbK2q�mF7L��eQr9N�S��)���8�X
�h;�� �����(+���)J�o�rV����
Z:��hvV���w�+�'"�c;�y7��8���`�1am�ra��
�gәx��W_.�2���^�������,Y��{����҅Tu��)���.���_O-`�]0�����adS����%����B���.E�ƪctU�M�4*/�GE�����Z�אf���pX�vND��T��h��r����#,��%��EW�g��R�5��"Y�x4���Z�Ǖ_��������ǳ��{�sEc���ӛͨ�d�W�'RI���9:�yd�~DY��\ ]ȷ5���0i��B$	
>�D�=^BVsۄ���򗙍���x�+σ���/���+�_vq��Y���D'���Dۃ�|�?�H�@`a��3��>�W���X�q��L�y�/O�MkX�~YYe��������K���L*{ۭwP��[�Ƙc�7ΜDJ��΄��Ru�o$�7_(l�r</d��#���WQ&:�L�:r���á���i����Pʓjk��`0���F˔I5<�>"�=�B76�������#��%@h$�,�eɣ�3��d6ϻ'��gUI���K�d<�suC.�aJ�"���zW�]�&�G���V���\�Ԫ�oM=`8O�t�ō�ҙsa�1߮T{9a�14N�^�~���L����NW�/�3<�(��XL���B6��&5�G(��?�4͂$� j��J�s2��M9T!l<�.3�YT�f*X�N�0�j[�Y��0�G�+��$���S�duuS(JoowY(��g赀IO�~|���`y@S�u�l���8ܣ��ѣ��/��ޠ}2K������=�(���}�N%�?�v�-�LUWW*������|42R�ٌ=!`���1�$0#!�X�R�#���@���d�m�c��$~���3cG%MB�*�t;�˩f)>hA�c�M�,Jn�Ҍ�	~(���t�@�a�P�c���V*��.v@��o��Z̄\�Iy�	Wʔ�N�cL��TX���?7FM�v�����岱�㭷��x�{��N���i
#f�Gv��h!cD�2pc+�9�d������l�ʋ�go��w�������5�V��_5�j4,�`X��Pu��s�V���I�1���-=&���X"#v��U�r2�x|�eW\1��ﭛZ�-��7?����~뭡���i�yMc�[b�3��a��Y�N�mZa�Z�;�9Ҽ{߁C�ݑh�%(-�NU��/}�;en��xH�e�ԇ��߾���\��3��sђź����W�4�yr߷��ݯ��y�*[C�:�zJ��ӌ�7�*2�Ь�9~gѡF���㽊d�>��H'��y�/�LÔ�W���e�52�ǈ.^v��{tx�WlAQ���c<�/a
(�.�`�꒮�kY��K�|�!Ͱ���',&�q�ܑH������a0�]q�0��f f�$˰[a½n��r�Ru�	�@8[U�٢�,˼��0G� ���UV�����
�L>��K:)�J���#�O¬6A�����Z�?o�G�����������c��Nk�M	0�,6�?�fm�}��X��+�v5w��	N]ͣ%g�R2ʑ}�N,���g�?=�	�=��������ǋ�,��}W���=���_��!Z�JR�R���Kb�3�]:gNӴD<����}I�`����I�R�m*�K���1�6>�L���)qW�1C��L�FlR��nqL,�1-��~<��9�3XK$#�cAA�J�@X�Aӛ�걧VFl�b�h��o}7�������EB+��V����y�j��X���b��0�I�6��N哑���GDS|�arm��L\>��4�K S2vv�L^v�;�yZ3=>��	��w?�z�{/�̥�_�ӟ�x��]�^RUU�УY�a��KgSy�A����
$g'�~�*H(�#���ߑJ�j��xӧG�J��w�|����y�����gW0?~���{瞳0�c��uX���4�;`���v͚>�#���[���
\_2�E�z,�L��������Ͼg�h^ӱÇa�+�.Y7c��i�ҁ.���(�5��&��:X�p3��gL��㉺�_�H+�ef�W�f�,P*���Jb��+H��wy]��7��7G|���D��sF�W������S�}j�ޱ����s��֧��
��Ioӈ.�V�o*�����Ɵa'av���b]њ�d�H��{������ʪꆆ�N���uI�����3_|���Z<O�LH5'2���k�k�i�)Y�e�w80�2��+��vU�e.�c��I�iu����װi�XQ�r�X��0�|�b��
��d9\Y���<vHAR!���l��ip�N������ۻ<�}<a @l����Hk�b�E����<h��x݉D���[�A�Y��Vb�f|ya>�6�	��/��{����^u�l�t � C8HSO&��;L��A��X�����N=%	�H���ϳ��"�ɤL��Z��i�2m�����*ʽ�{�~Bm'u%I�pB�l���w�I�8-�{���������4o;�xec��cL=�w�\
(�r����V��^(h���y��d.��9�9]7U�(�t�h�h�|�%��2fh��x��������嫖�*C�x~8ɘ�B�6Q��H�����rщꜝ`<�j�s�m�~�k�ۻ�c_u��ܽkg2����=���k�<����r����2C���֎hDIe�֯_�C�ES/���Jtp�Hgke�%�Z����Ǔ�ù��h񚡮n��pr�������ӷm{3Ol۹�x�;���+�kg,�ĭфV��GF��f�"k=��c��`��~�<�k��5�U�׬*�Z�.+��T���2Gjo��V_���TVy'5TT���z,K���Jo���~���]��\���$�.�E2�h�������Xi�����2�~�3�i=��'�Je���.���p�ْ�lim�����_��߳k�cOm]�lM����jg
���S��L��ASg�
F�@oNp�}�����o��6�l.��M�y3/��\�n"�Y�q$��Y����ޞ^P���#�?����ghT�B!�T0����B�\.�t:�ۏmi����4��	+9��Hs#
'����?3�yW�3���p2���7��H��5kV8�Za�"#q�YR2:�pF";#�#H��S�zV-�xM�`�6\�,�CWiA��ӯQä���/�"(a�����
�`�mX_n�9d`��(��>v���W\y(��������ϝ��I&�7,�N�}6�L}�)�U�rŜߩ}i\�)n�	2��['>1�gBP˶(�#Ñ�D"�A q�0fO�6=�e3�hdH�,#��2(����k����Y@������}��˯��o|��ѻu��������o�g�������;�/l۾]������|�{w�}gÌ��#C����]����_��ǙT�Ё��=�H]��{�6���3�̞�k������^q�۶m?޾��˾��g�;;gL���<|x��ԑ#�g7�:r��c�?�g��G�+[}���#G޼��kabd8?�+1<24(W($��vm�$N76�Z�c�iM��8L#�H�1D&��^�5k���׿��������oe��g-|��f����&�s��F/���	���w�TUF���s��{G�}��k�������fz�"��}���8�v`������e�(���gO�@1̙�9o�ŗ�����ѯ�8:sɊ���j�*��U�aU�E�H^m�4���7!�<qy��`�N�ݕ���n7�d�����W�Z
's�=�z�/O_�E3�=��;Tc+n�T�M�Mg�H�2�����a9L�
C��)"�D�-�d�Tn��Z9P���>x��8+���7���q*X�˱�|�)e$���+++9 �`<�暏&�����c�"ThqS�,�E6{GG_��*X�`�ݣ�d"�
N�KS�8f̎�J�,����J���O�"�W�C�E:�A�����[��h*����������=q6����3O��z&�eTg.��l��cu�E�-4�0�$�.Z��XH\��̦ޣMb�6E�g@�c)��F+|�9�-D�������v�YVV}���;������k]���<�r�E�赾�2Oںĕ��O���x��~�,bZ4��y�O�T�2W@��	����aD�Hn �1Gc���W蜷��{�W�Kg��矵f�?���[[�ܞ%�dc2m>��'+���<���\S�0����'䪨
L�`i�z�-V�������dVK��u�4�lz���F��,]x�UW�]"H�-[��X�b���}_zvR}��������|&�����a����A,6ΜY��'�5ᚆ��۷o���>�s{����&2	�S	TS�y�}'�h�p������O:�y!�1Mɱn�y?{�Ϗ?����_x��Dt$I�u��k>��e������<���m���-#!"�����<�z�7v�hN�DCu��0s�r��n�����}}�A�A׸�n$����j�l���y�>������f.\�l�?�|��W>��O��֋�Zr���Sj��n���+��"���J*ψ2 �z�y<�l���׭/Pc�_���`*�sם>yF%�,g`;��K���	Z�h�"v�Xž�{�y����q���`E��B�e׺�˶�������*�Ss�X��Qs�HӦ��h���� �,^EQ&����p.�nX���F��k��?�1��I�TNr��$���ˬ�x�D�&�&�{�E�o4[G�.0�oX�����!p9�l*m�T�ĉwYNge�R_=p�'`;��/,��x�$x�'�n���y,�)l
jL �4+O�XN�9U�`׉�.L���K0֖UtVYR�
�:5�>x�PEy��7����Bƒz�H$9:�̦e�@�� ,�ј�IE
pŜͩ�����ϥ�	����D��~���M�HD�9��_����_�d�+<3�6.�ZW]=g޴������@��E�|�{�Y񑏭8t�MW��S�Ne���$>���/{������ƈ�����J���x�lɩ����;ۻ�����M�}��Ύ��TC_O���ܰaÖ-Og�ڰL��?=���Λ���-�}��p��Z��Y���m{e�o��]�_z�C�%Iihh�R'o}B�e�����u���H��`�a5�S
��U5�f��ib:����p�͞Y;}���ڵ�Ȃuk~��m;vϚ��_7�!�̟��?_��+����+VK�,�L�{�ڕ�$��b[C����H���HG�#?��C�Z$�rt��
��bz����4�3A��7�3�ý��l��t���ןx��L�0��_ny�������O�x���ț9�ѐK��)�������p�U�/h���{ ��rmx��N?gz&S2�$$$!�@ "J�"(x�ED�z�z��U�"6�B�B��FzO�����{��Z{��	�ʕ���O�<��){����y��­8#��h4���U�����w�я|��)y�$��zX3�\.�������O� �����\�A�a"V8D���Д�*�s��[�]|�/���fM5$I���{��R�m���O��@T.���PzU:5sEC�H$�yǜ�Q�k�A�3|?6����E��:^�k�@��C�!�y4G8R/J��f��U�"�`�K`�=�Q��gY�HHādF�G��\^��O,X0�Xð`b�G
-"&1aŃz�B6>�>>|�K�
�F��c]�QƱH��জ��9W�H�� �*f��E�_�o?��O��#^���J��x唩�J���	�����a�K�M`z�I���a��ϻ�?��N�%%�k�a�P�)>UB/�P0��K���%g��������U��?����o���G��54e�|�ݱ_|y�s>~�%��~��}w������O]��{~6��>	~����76�����b�������oh��ɤ�=���w�'M�������?�r�g>y����/��S�V���ka�d.��,�&�Dj��'�j��G~͵���LzP�颞ӆ
��l;ܛ?p�7(Gz��ܼ^��llk�,3�a��N���Lo��W���EY�F����}v  �j�MVB��>K�9]O{A��LJ��؍���,Ytbp�jkYdj�]�M�����f��o�T�d�m�6\�66�C���r�=�5���0�_��/L:x��p���4�y_.V5e�Cj��L�	%H?���)�>� ��^хw����H�ǈ��ne���o��"�j	����oٱ3$s���Ϭ�?����r4�H�c�a��JA�D�epk��=�i�T\N3���ݷ�	ם|���h���n@�%�L]'���Fjc�>��Fod�u�`�"�(����BQ�XN�H�tH3�"�\q+�J"��"|߃`S�ȧ/�	��v�K�ض��l�XwP���ҁ1Ǳ�(!"2(BXO#��XS7T��i�&���2��"O/FEz�F��t����+~1*�Bw����'6&� A��C�u�f0ظq��H�֭k���}�i���h�С�u5Q��c���
&���0�(s7{{��Ԩ�g���w��@�!��T{�{�<����T��>4�w\�>��T��e��5��Ƒ2��+0�00TjhT~t-�D��'o��OtGS��ޮ�B4��C�pӗz��Ug����SO]�У�����ޚ2y�@_׽w�{:�̝֦��͙j�{�}?��0�U��U5�u���ׯ��{��O�{��Xhi�o�Db,��������g��՟;M��_��tU[v���L1ʰt�����9�Ro�-Ggi�OɄm�¾W+ql񼏜�f�����+�@T��A��3ӣo��v��XX�<k��r8�EQZY�����Ŗ����wLF�v�����2�岰)F�Ci�x[u�`_
9:r$�-�9�:g����D`���9�V���q�B���$-����jΙ@�M�=�7^OO_Sd��g��S@m3�X�rv_r�����bh���3�P5zU����_��(3���&Yf�~�����e+�8�J����<R̞��䏭:��"�_���
s&ox�3��צ�'��F'�>�'�q8䚆j)�*�|�GC�mr��v̳V�ɺE����%R��ɩ�~8��h�/�J74��[*���p,���p�jB�q�D���l8��T��eYR�V���a�V9p?�ˤ�.<s+���1�)�v��I��XWW�����0i;�~��qc6�x���.�&����G�C(R4f� Ǒ�)���6�h��8>�P�j��%�������PR�V���*��hBZ��oGG��m��<�c5��>���',^hV�X8|�`4r}��4��O�l�6�3��cӤ=��Q�)��{ܞ�dks�c5�����Y��ϟ3,�m[^�0���>��s�Z�8.A�\}��é�k.9�����M�><���q5f){\3UΙq��Y̦󉏝�z,���JgMU�i�u���p���x����N�W���\_�����[���xߞ�,ť������a����������ۮ��C!PlE�ͺn^v�L����X'x�G�����}�D�:��fMU/#ÁUz=���@�MB���v�f+Pr�l�P,b@�l3���x�r���ҸFE�3�k�������B1?m�lQF�`5�2i������A�����sb��BJ9r��,n3�E4X���`Y�������8O��fq=l�Y�8+V� K�3�0�����׺���/�9	۽z��m,.�2i�AcV� �UZ;H�/�m��΃=�^{5g�i�Uu^Au��m_�U�Y���
��&Љؤ��BY���&�5KT�GwJXnM��."5)��H86����<z�0�.	�V"�^��1���x�E#����+z:�^~�Ljx�1?@jQ�\D�~WYE���h�ǩu���e��ɜ�ɽ�@������L���9B����F�Ы���L��%��Ū��g��q�|{��n{����,[r"ŘS�����*��A/�5���Rc�C���z�~͘>��3ށM�+c	�3��0�*����PS��rK�Ph��C��ڒ�MYu�T�N?y�aX�t��w�#K��˪@�����%����b�ݴ��D�*��Nl#Q�Ģ��IEQ��7#i񜮖�Ml��u�8D�������=�{w�޽L��ez�RB������~򓍍1�I.Y2[W�Im���ۏt=��R���HYy��p�����v}qB��3��22t�ȅ�R�-��r�f�%ܠ�bKf$�<�".�;Tp��R��VtOj��>i\M�����4	�ӆÔ���Y�2��Y=�a��)!��FF]����eut�l^�l������Ѽ�R�Aj��Q,�X�SЊ�D�Q����
�Cx�*��o�����VG�^�^4��2@��Ǧ�ʑ$i޼yF ���Z*a��]O�fO�6�ɅdT ��&�M@}�=ʗ�F��낑�ͦ#���SW�&nݵ۶�ViXcv�`	��"�t�\.J"�~�\��G*���i��S�0ɐX,K<B�wpݩ_�fy�Ĉ໹be	���RX�+Wku�:�#��!��?3ƞ+�X,X#���6�J�$��0��1I��1���B�h�|M�t$�$�Ȟi`m�pL5`c$)�rp��&�-D01~���+��00~�M�X��*�n4�-+��t0d��0a��'&S� �kjj�_��h4�	�(s]|�i�0��VJwF�>��7��1���ώ0�:���� ����3�4��0�UUr�-f��p�t0YJ�\ooG{��+/��sB<�X�b��N��j@8��Ԝ�p
x\Ρ�TI�lj_�t� ɩ�~=��'#�[�V.JH������T�&Q�u�[��7oނ��x��H7\�@�,3�|r��޲����>eR[O?H��I\LK���#�T���$
#a�j��S���U�!�:ܞ,ۦY����A�ȱX�����=F�Yuz�+����yh�w �w�h#�A��}��s}�̓SÃo�ߏׁ�A`�p�K�� 3�'�  ��IDAT���Y�aB��0��LG4���o�lG=�T*Ph8j�̕"|`jc���&E#h�'W(i��>Z�pT������""�D�05�����<�z�`���!�� �N_O�m���oO��cl۰tC���m� �|�bu�{�K��GҦ�?���W�8��}*��L �v��A������]��$��Q]ÿ	�ö�H� �fF:F�_�fE��R����F8\� 1<��PiK7i���	������8����%���7y�+���'��}�b>�(�?�4I�����Cx�c|�$�½�`�l�ٚ�lq����uԵ�p�R��˘<+�/?��)-�"(�*k�X���%e2���/�5�	�!��,X8שQ&xM�f4;��P�]����PI�;F�z�/B#Yw�3�����wV>4���U�_H��׃v*覞E뽈�rG\��׸���QD��H�zs�@��~��I�����E3p�E4f5"dF�e����to @�յ����[�-_Y][�I`���MѥB��,�/ť�Iz1��a*T[V䪪�Zʃ��jgW���Mc�T��B8$65LP�v~�4s�,,D:��P�1 ;I"{�S����XuU˶74�lS����2��Isy\����=������.��X�q�^R�����b���������6Oʛs+ӧ��Ճ��sϼ:4TJg���l:W��x(�[��c����}2�k�!dǦOo�8���?S�=4�5wɴ�	u����Y��:�&��l�{��q��D\9ᄙr�X_h�MX$s�!��#��z�ydw��j������(���{�[�oh ��M#����m	�� sJsqiMsc3ؖ5m�N�]�fM{�4u����sΜ���|ޫ�&m�&���taj�DۮH KY�VFa5�pA�8��Us3�a�T&7�����rװ#}~S�=�%
;���_S��pE����66�ۿw�KJ>l?��#<Qd�Q��=C�+B�j�����s�r,Y��S��q��ű`��v
����4'��\M�@�rGO�lWI3pF	y����`�E�6.#�<� \GA��P��P#�Z���}8��$__M�����~��AV�0d�'�o��v5��oi�2�%
x:{��?3h#��-��óm��L�Ew$K��M[���z�GM8|�GJ����šu����+�o�׵�c���|0��CW�0�h�
��������4��H�%���;r�/�7�5O۲y3��}��$�f3�s,�ځC��2Vĵ��T�ep^� "�b྇��sM|�0jB�e�
�XB�4���?w��;߾��:���u�p��y𑒁vF{w��\���Y3�r�gc	�IH5�����n��~��w�;���eKQ
����`��4Nqa�Q��y�u'�p/1���mD�5��jIE��ؤ����OX������<@A��X&��X��\�&��N��1�GX��w$���tY���~��͓"�H2��(������z�(7�%��Z��8�SA�ӆ��Ԙ�	h:�mZ�F��{�@�J
:U�J�@���p~�����^w?,*����vP�('�
�-;˂���������HL� h�����k�|��q��-;��-T��]��-���� 4@˿6�DI�[25Ь��!�%�es؆u)�ۂr���`����`n�m�'ab�o.�� ������y�o��)\.A4!�#}M��d</��]��
�����92R7;�3�á����\���h��A��9���^7�}�W��D֒9x���}��G���k�"�c)�iZ��"`Ye%bQԞ�^�LF�hɦ��ax#?��r�M�x�P M����֊a�X?w�sY˥l�OqQ�mp�M��R[[?z3��m������yBH	TM�v|z8��L���10���Ц�L�u<]���ְ�`��+z�f�5�|����V֛���g�g�"%�""��P�E_�����;����~��*Q�8����ӹkϾl!5}Aۗo^�s�u�u{zw���mj�nk�c��~R?�熳���E�������7�$�9ʃA ,����I貸��ɋ,	��bo��*�����L��
đbb��_�|{v��>N����F~XV�b)��P� �V����|k`�ߢ=C=���-�e�q� ����7�)�x�A/IG���Zi���/���$&L��x�4\�n���a�}Wـ��N�\t��D]�|i!�>\j��1E��g�����FP	����[��"��DЋ�Ai?�E��'����W8c���L�D����@���$������z��!��l��r�z�T�,��J�ӂ�a�4��q�̑8f�m��&;�vI�ۘ����<��n�ʵW�6��� 	���������*�Q,Ky�)?�B�Nb��m��\�_�%�x�*ֈ�����yb$3T��pOP�(�q.�q�Q�������!���q�8�����B{v�K.�#� 7BB�g2��,�:�>��U2��VJ%�{�<G�J�͘�8ќ�xQB^�r%��þ�t(fDe箃w���ᎎ^��Zۦ:����4(%: ���Nk��[ntl����`�x���P��Ks�jNy�1]a;c��F�tM��,nB5�h��S������a�N����,ʊ������V��;vmz}wG.M�Է,�2�^��Q�a&�5�Ѭ���hN����,���\1� ���h��4SQ'x��|����N\=����(��j��k�;�Z��qi�fL'b��ሼ '�X*�kϒ���	NlC��Q�m�0o޴H��q-===Q	͚�d�g3$�
j�!��؆�'�I���U��[��m�dcb%�z�SK��8��L�;��f��P��U0��v��,�����8����m�c��w�mٻv����^V��q%�I�Jx&���Y�g�\��"/�!>��x�����O�T8�C�"�a�H3�����L]�Ma�%�X*j��긴��Q{<Z���༂����t%�g��x�����8yV'VC�]ul����w�����c�Gr�Ϟ�P��(E�P��d<4nB*J���4~y+0:�F>+������U<B�!�9E��(R�vuwd��r0�%v�1%$˂@���R����h�\*t�ʧג�!��S����ݐ�+�7�� �eU�Y�fŒj󊰧���K.�;�HסB1����k�YG��p�J86�+8t��R�K��$#��Tӑ����S/������o5�N�w��n�5Q]��?�'����o��w�����/7���V.���0�p˄�����+�Bci�*���CA���;��bѴ��vf�:�>�rҟ��J��6U.j`�1%PI�tj��+��7����Iڨe�D���qFih�4��KNˈ�Y�PSH�1��;���f�ĭ������Idr)��t��p�(h�/dr�����6tG7��)�}wI�$�����[����'xL��������Bnr��h(�J�VĐ `�p��Ng_���K]�L��p<[�K2�u��;w�%+3E��������� �&Z���;���/�i9NUU4�nkk�����q�[�$�y�^	�_|JlP�Y���I''L�x���w �J���P$�p�إ�+�<4�H���)�`x�F�̷�m��h���I-K�/��~cog?�zwh����� �[�Ft������{�v۬`��7p�|8d���,�&D1�	��J���M`kp<�0-0�q8���@�ypM��y�07E����1%Ǘ�6� ��#�ฅʋ��<랂� [c��o;���qGr���ܱ��G�;ׂ�=��Z�w�6˩t��x��7�ʌE[�^!��+�u�6��{OI�Z4!ah�a�n����k�fݣ}̶�`�	$�D��s���l!�ݹw��i���MA ��Z�+0,k��C�,]����$�Ѧ�J�(H�Ly����>��7�r�)���7�ܺe�ds�ғ���+j⨷�jN����?6�P`xF˕	�:�LH�9=�(�%K�1�r�]�I���g/�h��y�yS�)l��]J�*A���s���wY���`�EPV�k�6�yQ�9���]*C�f�V��\�9������eЂF��ʲ��b0�3�G������u�"�↓�P(��#�VZ������	�)[/'j�@�Mg��T�kj�"�Z�-�F���j����u���Uv*���]t�,S�F-ip��ڸsߎW_y�c�P�Q0�H'-؟Xb��!�JKK�ʕ��^}x���{��;F&U:kJ�:>�r����N<+˿���������&1�:OH���:S�CI�f>$� :����
��w���pwW���BQiɉ�.���z���nǎ ���T���;�f���N=�o}{sOo^��`p�7�����'�-�V>V�"4��ol��(*UA^��7^��4bPc��(���OH%���ʲ-��rS��(m�!�[�ː.+�Zq1!>$^;�a�o�/�ѭP����֎L`�����
�����~,��u�#��9�`���4&�`4���_F3	��Mh��Z	��&�W8������M�pX.�ьJ�/��'M*x�`��d_A"��p,�S����W�%EZkn�R]�	��Gb�3��p#G::� �3������������ex���p
޼p��N>e1����}�ŧ�(�/�p핺Qxsë����g.YY�0��n�,Ō��QI�*�Tf������{����kK�&�a�٘�B��͗9>�@�Y2Eu�̹�� �58,�aU���ܐ,��J�%b��< E�&)�!�]&{��;γ\(W`7�����_�X��o���?���W7�4����u�l�������k׾28�,�`e\z:M	}�?R�7�t�Ʒ���#�u�����p����+'N�{�/;��ȃM�W�:c|ø={�hܙ�T�\(��9��Į���?!�������{���?y����W_�M��cl���D��(�$ɵ���k�(���b^{���M��a��j,8|�p�"L�/j�ZOY/�u�#��L��%�=E��(���1�)�r�A�MQbA�z�� nZ@r<�l��6�Ƅ&ص'�x��{��Aj� ��qs��@0ڦ�+��$	��9 "-lӬ����Ɉ+׋:���y���)�����.v#M��8����n�LD9�|���*�׮��g�T':�ߗ����^ppx��-��n��R�G3~-�g!�Ht��*Ѥ��6D���؞�M����Ԧ���Y�X�i�`08�Eı�ٍ��_O�Qa�,�H2FR�FWD9@���-�_ΕK��ڪ`$��3�k[*�40�v!�WG㢭	��>��!^_?q�\U_�6i�i�\���?88����y������/����.��'&�Uoڴ��;cVs,���I���ܘ'TezFU��0�����)pT0,X�dF`�4�ᨵs�d�m���8���Y�J�,���p(�2^�Q�^���Q^ �afhZW�sB�FC�'?�iУ����Ĥ�;v�67lݷ_���{{�-���Sϟw��{���{��r��u�h��ͭ�ZƷ�-��;
7��8ҹ��|~��_���W6�h�������F������������TQ��x�1d]��W��� ص"���$��[7/Zt��6������ ���gN3�ǁ�%94l�f2�����WWW�Ғeβ��� 
���8j��d�f]7tU�ʶmJ�Q�)�q�wܚ�0��)�E��!��zx�hl'����4PZ�d4Brp�4qz� �S+F�)sM���׹馛��a��D����̷B�������G�N0�ňJ,8"�bmS����P� !��sh�
���N�ø���b�K�{�S��"?�G6lx��.;ᄉ� \w͵p��P�t�IW\qE}C|`8V����T&��ضˑ\M��K�Cz��5�(y�����;���Upc�N�nY�9C�x�X*Z�)�y�uÄY�8䄔���|�*V����>�)�o��w����ch0-
��-ӆ/��N����7n[ۄrWW>�/���	���E9���UU��)�e�*�"p�E��#G(� �W^u�O�`3��#�;v�
KҊ���>�T�
��iV�i�-{_SM_�ɧ��K:�pG�i���̡�|�80���T���;{�z['�����w�ܱt�I �Z���?t����n�����P85M��T�ml!e��]jL�ͮ��
+���^�&i0�G�F�<�-���-��7/hրK��`��fՊEAJ�?��c������p
�IL�1y�ɋj���ȸ	��$%�z��\ �S���#���ISX������d��3v��>oaz��'�r���}dB�p~��O<�f��}��ퟺh��olL�g̪�l�u硥'�q�྆��Ɖ�:�g���������6���@I��Q��0]�ƌ0��WS>Bt)1���,1�<lk�`8n8��gN�����1a[r�Ք��{����F0��L� (����~�}�s�dWґB96w)�mVǴ���k�z�W�L�&��P���G�xx`�6�NB����ihr�Iz~������>�r�\�چ=;�s����Y`AbY�aּh�G�@J;,��ӟ��5.&��X:
o���|r@7���pl����:�}�S/�t޲iC2�Q�A��T���_��E���"�@���
�G~�M�E������-��n��+wl�K��o�4��]��[Zƅ�M7�[}AH�g���Z�.�j6�G��Gzl����̒Q�Z���
��`��eZe���� #lJ �K����O�mh/���ZV¨�N��#�1u��H4�u{,�ܡ��&_.򅬪�ҹ�� F�J����P�����Cu}�L4KJê�q���p<�(�fC-����#���w���M7\�].��??��֪�QC�!��pٮ8�����H*���z\2-��k�4`�T&��,�QA�ETS�p�'λ��?*�J��M_�ꭻv����~�sۆq��SV..���/�o�r�Gϒ$*�C��QxcqyFz"w�a��hiFkjz$5H�*Q�JU��ͦ��93��ҳ~���,0�h�A��W^�pn�Lg
��k/������ּ؝j_u���N\��.PӸ��=��dH+-V2�uJ����p���_�{`GY^���P4���&�Dl��KO���{׭���D�{.8aѮ�����}�����z:�Tu��_��e۶o���"�m@J :��hXz���7m�bh��t.[_�<�#���uy��0Z�M��՘�d�)��ieR��ޞ���}��ٿ�����P/�ޥ�o'���s饀Cz��!DΠ���&���-A�B��Wè1���E&\��^{C��]�)i�
�GX�!�\+m�� 8����qL~ o@����gAi����}�А,qG���9A8B�{����c#Ђ��DLċL���w���P�׍8���Э|���J��m[���pYQ2�������EQ��*���f�=�&ͅ��뚆%��-�ʪ~�g���w�{���������4��������2��l�T����hpQ4�6\�'�#���?3�q��K��Ff�e\����[Bf!��WF��
l�FJ%�v��j������R�1�VQlӠս�}�h�~��E��l��"�Y����(�X��Y�䎛�d��	R(ܟ�=��K���XtBݦ����v��2u��jz��O?����ӕ�D��=��TAS������N����`���8&@\l����R������K$%���4��#_tm��Q0�,<a��y�a���B��+W,8a���� �d�Y+A�~��	�PP׃]En���xp�q�V
^�Q���2yb#���%��F �i
C��L�C$�T<J/[ڼh����R|��ɑ��U�׎G���;炼�t���"�2����npxTG��&т��r(��lp����ǔq���L�R7uz]����\������b1���Kϯ8i9|VUsS������ʺW3��U���&�:��U� .��,�����@(�Q(��w�I�g�|����߄� ig��-�,\�ʰ�����&|Vy��C�ᮡ��<���듙<'
'.\�r�b��$X��V���(�T\�I�Ƒq�~98�Ǵl��d,IP�d�@XH$NђA9���5� ��\�W��!p�8�?�����1�#����Y�j�YCcI�O,+�٭�P�ǵ�c���9��0J�H��dq�����X���C>�Ş�uv�����@�18���x��^�D��H42���r�D_#�6i�ka�����a��ȭ_���։�t�*[oo�Y����k����;��/L�2����<��/�˻ړ`SB\r��+�Xt�q�+�je�A��n�vߥ���MO��t<N=�{��}��|�Ys柲��9s���8��U���W_]��(��.����j��R��8Aì���g>����Ζ�	�wޛ^�����4gsC`JgYp�M6y����\y�Wg�>^	ƾ�����w�{���׿?Q�Pmc͵7��e�]���?R�ϛ;w�y\��#����_��ּ�3.���x5���j~��]%V��B=ɤ[����<K��=�}�t�t�B��˗���}�p j�j'M�RS��sߓ�X�ssN��Ă�Ϫ��}�p@��X$.�jY�xX��Zd��z.=�Ezr�l��+ͳ��9K71j�{��Ԉ������<7.4P$N�I7%s�
��E�a�vrp^L�)���e)�2���y���Ul(���0͢�/J@�HHM)�8]�q�-PS�k����Qc�|��� �.��V��(�^{y٢� ��V�魵_�Ʒ�rJ�
�_0�����q�ū��@��#�N��d�xw�e��͛7oڴyʔ�B����~ۯ���p��-��ш@#��ޗe4r�|Y�x��)#�}��s�/#�����[��tQ	����VE-���/�Dc��w2��@+<�ӡhԛf��V��HsԈ�9�!���DYvm�E-*����/�4��!r����,�hs�����qL���^|����#	K�V˶�ʲ��E� ��O��8u�1l�Y�b�H
ӟ���P� �0�T w��h=�cT�6u���L~����~�����A���<�A#��ڪ6�ԝ
!A��S�����	
�"�ps������If�w��iº��/=aY����Ov��7�p^����o����(�T�����ۼi�䶉ͭ-���cY��G��jc�{�@zUD�9}̘���N�߮����[A�ڽ��;�,Y����e�5�jh�����+$I���[�lA:�>p��}�er���{����:��ƍol�X}h�s��z��˘���Z�6ʹ����ƴ�Dz���Ɏ���mk;&ϟ��_^\�t���]Z,�ŧ�0(���G>��fN���۝�Z'�]�����66��@�G?�9�E���X@b��CaM������di8SNR��7oE��CCپ��V,�_��s�eom��«����xn�˳fM7���~��?�;wv�h�����O
9# �[ƃ��8:�ɪ�j�8uC�C`��k�0� ��4�-��`r �%E��\�����E[8�ɲ�H��:Y]/(I�2a
F*�\����I����Y�:�~�ܕלE��"�\Yʹ?��i��t��iW�"nh`��;�ҫO��5k��C�t�@�x�c��|~8�e]��E�D�.#�`p�.6b��#��TWɶ�+��Ҳs��S����x`�T���-���;eb�������@�mN�k6V̚��榍���ƹ�/�&!?�Ě��x�L��o~��H�������ww}����۪cs�a�6`p2�F>���L0>eM�p�駆upf0 e��y�cP�%�xn)���:�G�U"`{I=�cKc�k>��3&>�!b���Fep#I�L$�ʙ6��dD%���bq�cxb��S��P
]xL��c��-����۶�ܾC�L��x$m�4�2@Ҽ�A#0�
�pQ��pC��Ȳ�sh|A\i*��f�
����ԯ��eO<�����ܾ{K2��JYQT���X�-a<$�\�7��p�7�.os�Skx���g>;g�mo������o](�5��c�����\}�ym&��dS�=���ÇO?��+��L@�J�Z�c�0�-�����-��}�����'r�R��r�lO�|��6�]���	����o��o|�j�-�A�φbN��MT�6@BEk`��@0<iZ�`W ��d�d=�qAe%�����~|I���&��94a<�F�D<�M[�<��?��s�p�=�<�Q�Ф��?<����_�s��)m�l�O��A�nѴ�@�7[����z{{�J�����e��������Ñu��?��Ú��/��m���;{r����,/��5沥O_x	�Zk��t��\M@�@�8�p �MO�0n8�W��a4p�[P,�ռ.K2\���2qB	��3U�=��4���HkfAt�тΈ.�.�/�����ϲ��[�~��P����g֟q�Bs�I���`'Z�P��i&*���p�x(�

~�%��f�[:�8�X��*�2C���2���*��e`�����͘1������U�;{Ŋ���J�3'妫)� Q�5�_����߃#��\we_&�2�ն����ͽ��)���NkK}c}�6��ji����T]'\/nI��0C�j� �~��q)�vu���`'�!	X�������k�<~��������ڰ�ΰl˫;e�
�
h6�'U >�˲p�\A���i�_���R��mq�8��߇��}V��}�qL~ ��^�8qb}ݸ|�P��J��N�_��|^I�G��e�m��ˑ9�V`Hs��I!p��6L؝�4l�H,�q���CK�Y$l�.��$�

}�#������/��λD1�!M�$�}�P��r�7���*Qb��ݧ�9s'��T���`X֭"�,�17n����XSSs�e�-<���CMU8�+
�X���\ܪ�9��cq�p4C��SV._�x���ۻ�~��ݽ�ŧLkHfߊ$�x����Se5�����k�rm�2���V�̘��ɡ�e���0|h�KC=ŪP�^0d%3�MA-�?kɒyk�nh߷��;���K׿��/=�rL+��twv��6����)�����h"���6U+'j�Է�MMgdMu��Ҁ������3#(���&�r�������^|��L͝������=���"c+���#G����:��/��/��Hl⤉M��%z���ɺ�:�=�P jx��.΍�j�b}���ۻ��i<����ylB�B�M���O�2i(iK�*�@k_����d�����q��՛�53�����w�IM��������$X�WrY�+�5�yc_�@uuM[[��� \[_�g҅H�n�t��[^e&h	����ƫ�D<顑� sؓI&	P!�rA����f������b.�pE7+�2\|�\�G#��UNcC=l ���`\�g9�Z��Kj�.��uU�Ě�(�8�7�c�5�up�'�N�ɦ���ap1��w�b1Q�˜��%]�f�`�j"��U��7p�@�ن��S�q�|
 �po��0D�b��)E��Dd%X e
&-�`�Œ (e�� �H�1E�ό��R�$-0��h��9x(_��&��a:z#߃k!�����q�2�����Xޤ��6AF�,�:E�5��i���~��%G�%#,Z��ki-�� 2�dl/&�V�ft6U�#ƃp �_���K��˻�H$x֪S���@�Íd���jA�}����/��A-X��'���X�:����O\W���I��ݲ��=u꤀��_���/j��:|��~�b��\>�ٮ�v���olx��U+�
(9�'J����6���y��0��
1���L;�M�&�p|�Hk�̰�SW�9�-`�������#bI+=���o�������훃�`<$��|���{�)'-~����Ξ�R��y�O~�l:��K�5k�9`�M�2,�m����c��ýJ0^�Ќ9t����`?(�Djй��_�}��_��fQDj��J�/���;�ޡ�ʁm�� Q��d�8^عk���`����t���kŊ�}���t��79�1y��\6�wJ���o���qۭ�6��v�'�|��g�9�����y�2��A�')#!�������O������+�P�J���׼��'�|�MS��?��˻v��[��ǭ�����KT͝3/��9%�z��?<���G&�N,��n������l;����ɲ��]r�r� ��Kp�����k�	��GN�>�ĝ3(�l6+)�c����������Rу�+�Z*�
y�'�ݏ�@?8�Ƃꀙɀ��Qc0wn��E�,��
1OwT:5BJ貽�ZԘc[��,��]���s)�d^����X��R�f�4<kY:�S���8��7jERG�_ax��qf��apD����pł�h=V�IJ�P2*��<�	��Gxl��q4!�D�h���!Ch�1�J����GY�8��0�6�eb�@`HK#�?�qS�M;��O:g�|!	�R�̄	c*b>��+�43e�F�"����?���46D1p4"Ly1+�.x��p��عB?�B��8V4�����t�mb��.����7����Ԝ�盛�E2+҇� ��5P���+��#������|���˔�eEQ�������wW^�Qs�̞3g�}�����\�2��쏝))T���3w����/v����!f��r,�=���o����D��F_yf�e�K0�m�6���ۑu�	������W�_�a��̫��xZs�5�]��+�Y����M�<qh��O?r���q�X�"D������M�u��ٳ�^�i�H�S����O޳{�����Ib@-��u٢%�f.Gc�:�cw��3f̆�̞5g������xŊS^|q����屇A:�JO�4���4��I�� ���߿��+V�zro� X6�>��O�羏��d*��S�nm��aC�e��k�ݶcg({�W��̋�Z�q��GJ����5i�$\�E3���K�T<�fy���6���?n��_�����x��-M�>s���5݌%�� ��҇��C�<���v�}��_c���W���P���/�������B���o����Kk]G��mW57)���}pY5��N�6�C�VL�H6?�W";���L4�_��5�(�4"��X$�%$Y*�e�?�,�Ҧa���u����a]�� GBfi�����r$I7ܴ]��Z�cy�J� I|5�r����Y=lY����a�%xR$@��y.�x"�F:.J��QX������p�X��:V� �ީ�E�9@A�6}|g�Y��Xc<ޟ�k01-���Ň-LzL~`#�P$�_*������,�ԛ8��8�.Ip�!f��t�;nBB!�}`�24
F$Y��˗���H��}�_�$�V����p��e��i����M�ʍ�!�76!��!lc{�e(�&�I�0|�I��O=�G���� �*�"A�6�.J�Gu��0��WOZqG��(#z���=p͞=��k�p��(�џ���G���k�A\^��K-���\�(�8��b W��&dh! [,�57�E�p�n��c+��ҸV�q�l�;�����j��/\��-�$��Oj��ߒ$%GY�tŒ���A��>�f�s/���ί����{�%�e�g&�=�vwv����RT���Aǲ��l���.���;&�ؾ뜳Ninj���u�<a�_���3'.:n��_�6�n��Ox.���<���ڦΘ5$w��ڸ^;o�	����#�rm}c��ڸ�����S�3g��� (�%KN|���fϞ=mZk�X�V���Jp�ls+:�׀�s���E�5 8:}֪�׬y�_�)��-o�,�
0w�fq�N�@�����*QF���S�U_�M���{;������DGGwOw���O��V�at�������uwA�g~��>'��\��b&�~Cz���!d��!��+�.F��0��M�R�z��<��cN����(���Z�z�#���]p�#�y[$ ���$�hӸۊ�^b$)�	-�����x��8#�O)fw�4j��X&(�� �p1ZYkƶ��{�����H�a8l���N��>:sh�P���'#���8���c!"��</s�������p/[p�GGGѤ����i?���$�S�D���=��FbH�%"4C��q�)����H�G������z�$Nm	��4_,��bA�8������x�>d4��!|g��q�g#h,��X�RÃ�'���nF��j����������i���T_�(uP����$���P#��0�:Pw�mDH�.��Q�,G�;�8#�Gd�v0�u��1c��0��hY/A�Ba$�n��ޞ>�%�LҊ��m��ML�`Ѻ�8A��ҕ����N9�4��1�F�����C�I�̀T�9�j(���/v�q�x=��j���j�`r�1��g��ٗ���sW]}S:��.�?�S����"N�%�0('E�D^p��"J�u!�)��YS-͞ڶ|��V��zV]0�e��M��bY��+��"6��v�&1?&�ë�e��fV�F�Y�.����y�/k�I�n&��H0A{��sϾp�'.�iv��%'<��Gn��W��`�������h��$�Q�T|!J�]t�i�6mڻoGwMu���bl8�l�5��$���Z��޾�ꚺ`���.bx²�_��SO?���9Q�C�Gv&ӽ�*Pwww*��$�-�U�Tʑ�h�o~y�9~$�S`,�����}X;jDb7��qPGU��u��4�5��0����A����gb�{�$t-a�*{�|Pw�O�P����&,6���ؽ`��`ká6i��żj袨a�4�wu��@
	'r,����0��:���~1^�X�>��'T�%F�qL�3�(>B�����#퇻{�id
Z�^<�=`5I�&���_�AK`
 r"�a�&����p����]�����C�oۻw��n�������a�$7Ke�ᜀ[�x�~��ezaIV$��>��s<x����a[h�{�^���{'	l����+V����^,��,���;w䲅PPfǐL��
���x��`uS�}<"J*tNh�bl�6�UX�W�+Tj10�3��d6W*��r*=<u��p$��W�E!�/�JN���>�YS[�u*�C�М �d�=8b��L�J-UT�pɼ�6c!�W�Z�Y5��2�� �3���*	J�-EB�A�Q�a��L��|���P][��4^��D$Ɨ~��.Z����e�����Y�C��W<�^=
(`[�	~"AS/�ϑ˪�̹���{vאָ��E�s�i�԰n�Y���}�U^��x�h�fF�"��<�50�F�lf�7���vz8+�}��Ug}$�D��x<�߼��W���<��@;;.��-L����=��d\ΏbqmI�e��o��ҟ��#��#���ݝ��Z�xr����7�K�X����~�ч��D�:Uh<�����³�����ڲ��ĥ����w�z䑵��<���͝Fc�]G�]	�P~ڂ���(���ݿjZ��HC���ڣ|�>���${�{� ��,/��5p���a�fK�Qoh'�~(�ŸN���S$b����>���0W�lf���0
?I�ıY��e��t�eY���6��V�/EC�HVEh���6EA˜P��'���r!o�M�	#ID;���?$��"�_�w�#�ƃ>�N�#JKSXj�ZL&3�������ݵ+w<9M�L A��^����\EA� � ��bV��"����A$I��L���ܡ�Ү���U�}f�r�Of3�_�>�v�ⷾU(�����gI�+� �b^ӔL&�9�)5���2�4B���C�t�j�`�a�T�B�ؔm��׾6^v��{x�w���HO��@��Ke�S��ɬ����`�7�+� ���*��5��n|I˰9-�J�|tx�u<X������K�>ߐ�~��3��%�q���Z��8[i;��"��	GՑZ<44�Dr�I#��ɺ`j.J�sΉV*�p�mJ��CJ:ޜ�6��WU	X:�ǜ:}6�$b�3��'O+�G�t��2Ka[Vo;p�)�;
�M����p� �	r�b��
9ft�!�\3Ar=�5uQ�RIKg��Si�
�5:��9�V#ќϬ[���u�47��f�K��L�ܲ�kvM��x(V�ɠ((I�.
������g������L�|68X�T:j��S��*6,���F��*e'�M/[>��Ҽa}��9oq�1KW�.^4eʔ��>N�O���l۶:����_��+��kqy��Us�#ⲚP�=�:�s/yXnH�#���v�1s���E��'i��{���,�5s��9�5��.>��G��O�������Y�מ�;ӦZ�����1��O�x��;9�}���O��?�O?~oo��8蜳�Jg8uq�6Ya��'׍'&��b��*�N̿�)>C�JZ��+n�sR�e���<�`����
�Y��6l̦S~%p�G`>�\ve����xX�R�`������U�i��թ�rB��ks*����LS��:U1��q̙�"�7{�QG~�T.����P�44c6RըM
�L[�`h@��g�������t�o_Z�.�J�UL؃Q�n�G��(#�45zgT��V��;֮�5����3�8��l�t�eW.}�%6�/�NV�	'9wΜ�����1öA� ��6�J����\�$ry�!_)��n�qƙ�#�#�S:���-��E���.z��:]�N�a�>�vDNٱ3���:�9������#�u�2������U�V�����e�����#�s��=-�π"ѱP$$�
�
��c�y�C͔�fA;�\K�ۆvto�����H!�ޮT��0&��*k�F��I"?���H�5��-VUղҌX	�+�ǹ&��eYRs���l��
Ks%��[־ܒ=)�K�=�|� T�LРD'�ܘ�BypB����9�v�Lz�+a�I�.��M�l��i���5�͜=w��-s�����?��%�Gi��f(�	|�Tk��@F��d3�τ* 6+�]����ٵc�������!�~}���P���̷��!�f�J۶�A��0������/:���~��_����B]�R	�KO�P��4���{Ϳ��|�OSր�G4{֤�z6�hY��3?�K�~�!C�=<<�Qٻ��={\�k�jz ����I�:���Y���3N�ף������������П�!�����	�J
8&C��U²�֝}A^w�qCM�}�����o��w�RF]���?�G~x���_��۞�ۆ�z/���9��[n��������� }!r�(I���+��Z��N�������D5焁	���q�Hh������7g��:k��b����\��Ҧ"�������(T�͍����[z
�Vh�������T^�Hf��'׿�ح��Q�GHa�XfKN�b��j� 1@οk�_[�i���H��Ig�ښ]�:��h����|c�\��1�,��CÃ���@�62ƧM��h�}T���[<���.x�'�?U;K��F Ě�����{K��=�Zh[��6,X0}ժ�p�M��-+u���׿���~�ۯ,[n�z@�L��bU�<���2�5�Hɏ���/��䒗_Z���/�b�jH�8���"^��e�1Oxi�O(����|��Ķj�㫨AU*�1��<�q@��l&_(�R��LdU?�����5�3`ѕ��8Q�I�Uz�|)����MR�$�X�6�:�|�X��'O}߻��s���8	A�sY�U-w�� �Ew牗Yuב�W�PD���(2��G��+���{�vՙ��n��w��O�'O�{��F%;�q��I�r����d���R��vۃ��|��3V>�e���g�@e�<�dU8��:�x��͛��57�9�)�����)]`l���
�Ȧ���@�����sM��-Vk�X�]�M��5%�6�i�bx�f�l���x!�I����Za,�3Q����-��$�x��H�,1X��������'�|�A��������L�7m�2>>��Ϟ���<���--M���a����V���
Ɣ�یuzP��04¥A�XkA�h{��o�/i:���	�u�v�F���@�ި�R�	�T,��+F��;Rv��!76:�3�մ��Ċ�J��	���kc�"|�CIP�P�Mtx��+���#�#`ϱLGً]��{���Ѐ�=���1|G���+B���_.�Lmx�R��:m`GqӦ���g{̛��q�s�XՂ���\�kX�boz�:*���u ���^|᥿���O���^{q%{�oꩧ�P����g�u�~�46Vxf�S�������[�АU����y��c̄h���"�j����<�����b����T�|Ƽ8YH�/��ķ�)V�J�19�X�,TT�l�[��'|�G)fW=B�⩘�E��T�#T�ƲS�J&����a�nn�5���i�����F��%@Ԯ@�(����4��!�\՚U���oq�)Ϝ9��ԒJ��H�K%X3��
�iB:Ů�u�)H@D!퐈2yMM9�k�u��'��>66�l��\p<-�+��l�-����Z&eД���!�sʥ���g����W}�����1ɍ��;߱m�m[6�r9���dd2�u0�<W[�f���e�ɪ�!��\b=;�eҙ�����3C�'On�귒;0�'����	�FX{+6�+�@��46�F�������/���y)�	׬T�e�yi���١Ϝ=e���/�>}zK[��{<�й�}������ڶy�ꕯ6�5Ϝ9s�5��`��z<�F�ϝЃ��jAp��Jz��#�kR�+Y�d}�Lŀ�͂��L���_x��|h��u,XD��Y�~eO�BB����a����W_}�!��.�_�4F�#�	i�Ջ�PԬ�w�ح�Ɂ�9*�L!���G�,�aw�qتh�:.1#�K��jK�"��_���e�עEK���$�"?��y�8�������b>���7Ϟ1���}��C۲e��3�o�,w�Jr��gR��HS��>�G#�!��H<���֥K_.��+�.����<�ȋ�]~�SO=���~�c�nnh>�$���,]��ƍ�W�Y}���y�'�_�7��i&;�1%���k��~�{���eM"3)dvE��h6=�K%��\O�4J�S��`�f0(,B�3Tف��g��P�Y�]U�
�'u�!E�qTo��Ϲ�k��
Oi���EP��zZ��jd�V�)U� G>q
�r�O��qXbG�"	��O�X�X�z�}���5eE��`�Ӡ�u<1�ULS���!K<���&�D=/k�%�Ih�(.�&��	:�sg=�裙Lzƌ���pq�q`�?v�����i�����z�U�ȓm�_�jY�0S�f5�s�'8��r8)eP�L�*X6��z��6S��0CQ�a"�m����j�̙[�J�S��x��,�U<�֡�>s&sM7aoR�C�i�\U;��}g�xy�����hlA;�x(�XL�O`��*�,���T���^�?�>F�!�*A�:++XD�Keri�Xf�#�`�N�<��Iy�o/�x�M��ZF0Q�S�tj�u��.���8���0�N���\ú��Jw�q�?�1hA��e$���и��>(W��.}	�i*��ԿI��R��YB����G�D؍����꣏=�TC�ŏ�jqHU��&�[P0��n��_�nE��F���(����l``�����ʦJ9FY��_��kK_\)��&��"��鼖�V��Ð �p�����^Y��ϝ�N�K�10Y-~�-�xT���A!����F�TC�*���j�ZP_��?�~g��C�-�߿��۷o���>m6I4���[�`��=�4r���@.���}B��y�����[���~��)�
�ä;�X�b�x�i]�r�d�q��8��$���,�Q�#�%�	�a^�+5(`�i� �����(B�����5��h*��UA�����G��DF*32�-�l!�]},��
y�֯FvZ$"	��G�e2�+����(�!�`���_!��3پ ��F>�����@UV�O�D�H-�srKS��q��=�w�\������ٓg��5]o�ɸ�9Nf���*$�r���a�!���@�6��0��TT)�)�������hY[�5�i*�����
O!�3�� ��Uљ᱇�7H��!.Ίt�}?<RMM�����Ռl4�-�:3˦!�����]+��..#/%�0�k��3Yk�m˖����ԐqJ��? ���KW����^q����3�8�����jD^�Jlg��Y6���"C�.b�G�����I�M iY!�_�_E"0a+~��\0/�J�n+���=�w�ɨ ��I�] ����u�����L��NaPNh�������t��G�=LA��0�����I�Y������C93�!����I��;n��DM��c'21M���茑�y
v���ҥB$΍�(��?���T����,{i�q�^К5����֬]E�w���7o\�x����m۲�7X� ��u�����4K�4����Ē�We:����
lQ�6�m+� T�@�Ѕĸm�VYt�5�	g��"CA����(�����E,{�!#KM�v� {t�S04�X��@�f��0�/jp[�L.t��' _T/}[1��Ѧ|�I%_p �}Vk�V�ޚG�#~.�瑛�����k[ �eLbY���L"5�b���7҃��AR#��"���֪���x�zxF �]�L-P"ǩx�K�
L`�r��{(),��g3�
����3FNUr"��XL�*c+�v{!�R��8�-S�����Ԁ�dϫ�O�)���BCC"�Q�S_��� �I�ZQ�X��Y�����V� V 6N��4�esM^�ơ�q���Ν6�K^���\fq\�xj�"�A��~a����u7,}ṣ�9�[.����Lʴ_~ymWG�纊��J��Yqq5-k�Si+B��äf�~g��F�l!b�6=�h��I2�B���+�c9A"A�ILq�z+ZU��@o��� %6.�O��n�"��8�#Y��
N%l�w�?�[�͑0y�k�����&����7l��`�-�c5�?��GS��}I�g�V(�N�E�Եh�i����j�h^�h�O<���s::S#����T*�2�4u�I�Uy��|�f"U).x�����ի�v�~�N۫V���{�N>��?���]z�%�2#�~��Ʀ�}��9��y~%�F��g#��aZ�GF�{x"�:ՏL9[,r��1�$��?���R��I#/����0��ʊ�8UnsQ�'��H���"�j �T�ߗ[�!u���J�հ��2;x�a:�.�ǹ*T�ji���|��W�qeh���[n�ٷ��������F :��t�	b�b_U��(q/**%�18I�FL�"�Cx���ElD�5�dJбrT�aX)�I�)X�M'�&�FU��\�h�4�OȎ�
.K�J�n+�e�e)�ʤAW�B]��k�f̄	ܴqc�#�
�\,Ξ9����w���>��n+C^
E�C&rC�rN�]�b�ڶ�==����E�z0UI�Bkk+�U�L�"fPC�dM� _
^�"��+P�>zWC#��L� !MO4���yAD�to�t���`��(l�B���*%��g>ю�� FR\�7��&ݰ&O�z�!���o��M�[z䡿�}��)�����gR�W�zB4�@��Xd�64Bl�H�i�5�v]i�)��R�Q���*i�T�֨��,�=��D�lL��,	�1|Y�AhD!H����~4��j�Ob]��k��U�����%�nE��G������	~TO>񔭛7m޴����$D(}�ܞ�Q����2*ӐrCe�U�&��3f�T+�T&�{�=��o�[_��*��|vGYӵ���Z6��<�3e��lPr8E��c/��5K�~�4����[�b�^���?�������g?�����P����;NI��|C�{R$����I}�O^4�7=1��m54����k�����Ï8�S�pf��fqp+XA�|=�+��#J��B:$ g���T+c��t@��q���0��Z7a��c�8d�1��i!�=ay�%�aER������@a�\y�a{MӘ��=��L�o5�F�E(��s@�idb#��d����"fx��v�Am���7�yPj\��*�/)4	Y�]�I��r]�׫J.�#����W9�g�#����R��]6�!��}V������_j�A
F��M���cp�B<�J��X�A�"�����C�\��7��
��O�,y�`���W!CGėP�R��������߻Տ"���C<�ܳ���Ypc#�͍����R���\&=n`�C�i0�T$�VѲa�<ը��fZv��#jq�r(2uBn5��\�=���gZ���L�!��X	:Lq��T���<0S��*�w�a[�A"���e%�cZ)�Ⱥ
7��OT�B�D������y��4v+·5b���+�9s�̝=��{S��pM�U�D��C`�׋���iEJ���}C`��f��C���4S�]�z���:���Uk^޸����}�������(��C:U8�Ix��ږ5488s��r��Ie5ML�޵��gO9����p+|��SN`��FBjUw�(��#��6���fC�����R���������>��?ؚea���y�V�D��j�R%��2��ې�=yE� Ӊ���������1�UE(eƉ��*"��[�.<�t%��Y��1۫P��J��JT� �"��C].NR8��CC�e�du�HI�����:I�м E�<�
��rQõGDZF���7�.6�Y�:� �?�:l�jQ�_��>18�F��J?�ջPq�ɠ���}�1<˒g�)wr�R��!V�ٲ�������(�8W��(h��8﮾���S�QѬ1"᳉�j��T`�
zS�w����6�e���T\>Ҷi�6g�y�b
��K+����s�Z2��t�>���)�$�_�D����Զ�6��uN>�BX��0=A����8��Ue���%T��	����NZI5T��@����wB�ˏ݊�m�A�]{{g�Sv-�k�u##�]��2�mށ�!>u�O�����(FB&�ʚ��
=� ��IS�z���r>e�Z��BW���-ٽ��G�8��_�����JٵؗZU+�{L�m
��gT��Q������JeH�;h��J���u����g�O�!�����l��_�u��M�e`���㹬�Dy�|���3l����`U�cQP�\,c����ಔ�#%�bE���jh%�����ŐZ��U)R L�@S�����F�בS�EIw�X�J���L��s�JrT\��������<Q|I1�!N��r�Q�$�P&��f*V���Hե�
�0�2?�p�0������$�LP�jM4�	5n$�����e���#],����jΨ~>CƝ��cp��1�$,���Oy���7Ns��?�a��U&O�P��g�G�����U��!(B��|�D��
O�g;/䪓�v����4��M)�e9	5Á�����
Q%�F��`oz$qQy���N�6�߳n���������a8�<[�]�Ic��:� 9�TS�-.TP��TC�`�_GʅP��Q���8v+·3$����J��I�ew�n	��R9�a5�C���D#��66w��l!��x�$�$C����C����g���� �,nU��Z��
�l6��_��NM��G���V��D�󚚛�ǋ�������T���"X�`F�@�P$ՐV%ؤ̋ <_J����Vn`�V�w��j�<j��9��W��n�>iR�Y��h�"E���K�Q�S�Q���B����Z{S�Ža�`�p"v��bL�sNM4B��L�UN��d	VD�>�Fu�Q١�%�3�a>Xs�ᴅ�_k���U[A�Fң�����rF+5���2� BA*�.d1DKV���Eu�;�������s����~������O�����S�J�"wV�գP�#�Q�T�&2F"}�$��)�u���R�����f'6d" �`V��hL��󉱅S(�S��;�I۝0	�%�,�#���vCk��j�P$���BF�\�I�(�Ή�����(����u]h�VUŞ�8�ZU�v��dV�jZ���JÚ�تa� Le�H0]? J�����A��c�"�gG�YV3ÝJ�W�@���S}_~1a�E��&z`ΤW�ʞed�GI	���t��!���e�֒��uP`�:�JYᡮ+&A$�u��.Q��`(B�0j@�U�A��PU�����J��\��`�7ޯ���,���?N;�i�X>���>v���U�N���r����Gs��IjN-����ԭ�E���=�*KK�R�U!EHF�P$U�&L�p^.���kp3NHy)����AF�ZJ�����$r�]�"�8rt>�c��SlV��1�y	)����,��.���'=DT�	��E���L��bu+�6`�՘�R��i��N���$�y��8�⟒�W#e���4���?ac�Yo����jO>���ĕ���ɡDR�#-ȱ�-@���?G[���iD2��B���oE�-k��l7�@$��\�{�b�8b��!��$�O%Nt$��d�kA��O��?B�B�:��,C7��We�?�X6"�㢪����a��v��kF[kG-�MIRԳ�,ĂI��H$F~E�)�9`�z��켦zNe͚��v�'��c��l�������@���u{G�ﻇRx�kuA¶������4�x���>"�a�k@�y,~E����[:8|�N�����p���|4J#�C��"�E�)����Uɲ#U�(��w	ypB%���LMI����֗U����&"K3 ��1ɶz/�z�A+) ���v��f�d��Y!��a������h�)z�0ab7HH�O�J!-���7�d�9����ӲT�L�)������m0�iA:K�W���X�r�ӵYu�Ү=U��ѓ��)B�$v+�����Kz��{$'��	T�A25�p�ń:2�e	��b�zZ�Zr.c<�El�P tMI^{�W-��S��Fb�j[Rͽ���`㡢�8���V!��j�M%�EQ|Guw����uğ�����H�.0[P���"QH��\jR�I���u�')]'&I��J$���
?�3$2�J�,մp��mFJR3�Sz�Ņ��.��k���
R��CE�ѣ�9���L,rE��J	f�6l��IH�d��]�\L�k�-�N�RY��{^|q���J�H��b����\�����&�_j�V��숡�����eٜ{�7m��ơ���2��ؖ��$H>���w�U���Н!7�i����y`�ay����`�2���$Ԇ�?0L�\T���U-���ţ�H
($Y���߫��
AzЙ
�"=2��3�=��%���&�l�P@BSS7o�p�wE��(��A�x��Y���R�ʚ��b���������-_Y����9L���L$�1���*�hyO:1ň	V��5�߻���Qp�	Lj+�}l�]w�e��WM;W\QPK%̈�G�t�����RDRJWI�Io��m�_C�	DU�jr^	M��7� Z�mQ���X���#F�LXZa��`S^���U�"�%�f�*��yX!�X����.�����W��U�[�x�Q|X.�^��t`��zCD�M��F�,�&�c����u���	���7����PRD\HK+���U4,vc�%ΐ���#����F��� S´y%�C��o)J9Q	��5��y��^�E�
��z:�4�R�T�̉��W��~y����IT7m�Ȑ&�������`(3S5��M�p����,��*�m����Ċ�w�ح�ΨE�`'�]�'?�Ჿ/7?��3�M��BT���z�
6̌�8��)-�n5�W�5�v7م`d��966���h��K)2ٷ�0M�4Mɕ�[
��Y\�Dr��T���S2�$�:��) 臁i��ᱬH�ԅ��(ȥ�$�0�`�A\��G*�����nMu5D�2CaHz����)�&���T�"�p�˫W��.V�����i�b���Pd$��(4�RX�	k��E̲�;�:r����>+�g^X�����I��*%�hT�)�*�T�����+U�$=W1���S!�}�r��ik�����>��;TG�Ub� y�Q�,�T\��!B�������y�b8F��a�� �����cQ�؇�>VrԽ��ۓ�I�.�0�s���t� �KU?�`��v �5�E�
�nL��е[x}�b�]�zo���?�1�N�Ψ�5�'%;)ٓ�+�(K��1�5*��8�hz�`�RL
��ekH����:]�;��w(��PJ��F"r&�q�a��8��}��S.@}Rt��D�T�dE$+1��}4�iZ��<��j+�hy�sQv[MZ�#���L�Ե�3�e�Y�N/]�ꖾ�hR��un&����9���M��Pr�Z��q�����4��.�؜ٝ;����w���d�q�?�N )��Z`�+gg�sI�>��ϿK?��c�5&[`w����Xn�ڸB��2ID,�݈!	�����&\8lR���x��=(���@A�(C�KK/�x	��i�၆|c>���n�U�)(Uԫ�N*7`j��|�H)�4���Zf.Y{�r��
5	䯭�޴�d��z�n�DǞ���6m�+��tg�f����9�T8!m��R�!e�~0��5El|�̼��p�j1���I��1�Uϔ�ʼc��������F�s��N<���ʓ'�)�:� ��%�7����%Y1B,�dZ3r7�ɂ/~ERf/(˙Ld������J�L&�R������(2�F�Re�iOE�l����N��H��5�q�N��j�������S�\��V=�;�������t�ϋQ�p�N�����=��@��ኳ���s ��P��Y��::Êb����=s&r���ᦔB��=�� ����~���!*��OˈwR;+�tq�k���&��Թ���eU�1E�]M��@���03���7W|��v�E��?�M{�;�3�i�`��OO��c�]��wǌY���S;��5G��\��/�n��;�z�{���g3z��0y�ꑏ�ܿ�'0�w�E���m�M��Lb,�&N��R������ �8n[:W�8��)�wK���%}i���������ʾ�^E�m�6��S.cy�n�x㍠�o���%��ڰ�hhu���HZ?�"T�u�V�ow�,N���ʢ5����s��l��0�}��`0�DD�CQCEE�֒��GNjl��퉗�cq+�&���-};i�R�L�Ā�j�M���R5�/�F���Q�%��Z�T`�V���TRi;�K����������%'�J�G��/�'�Qp<ps*.�ʵ<��ʭC���&�%�"S���y���v5���P�̝�~�I�]���ETQuS�]p�!����0s�`'[��ilh����y�J4�����|�<����n��<nx�A wӹ��jd�|�J��Z�d�l������$�(5Ē�xr�
f���2�f�n%p@ӌ���lnjnj̧R�P(67�b����!p@�(�h�ܑ�����Lӆ3���V*�+��t+�M�)���;�*ef�f�\AxBy�-���]�&�� �ptd�i���5�t��)0������ȇ{���R�\�Ҹ:6Z�4e|�;=�"��=�����B9���S�	�?ҡw���1�@��pޒSybɳSgL��쌽t��k���/_r�m��k���������������Z�y��A���W�����O���{�l��)\3G�
n�"��xT7�;��)E\b��$"*S'�A%.^�ߋ�V1�@)�@W�4���4epxp��Y���S�+��BO�*�J�!eFiE��$/;N�X�Z6o\���X.-�nmi*	-�H�zu�v�Q�3�nE���F�.����w	�b��; �m;;��[[�:��[�@��&QޢU��� �&2`����/}	^W���B�:-N��	1��%�dV$,"f'4"�sKFUpО�"_���IV;.2Z�1_Y�*�}�-�:bt���ÏΙ={�>���}K�
�S+��VG��%O�u|��Rm�y�@-�3�V��T~���橼jE����ѣ��7���zv��f�#Ɋ�@ҫUY$����&Ɨ@HlE��aAN�u��L�>2�>�cӏT��|��JE�ͭ(_"*����ֵё�C�cڔ�R$����QR�$��CT�Y�'�)q�<��>���������M�C#W]qչ�[,�}jɒO}��r�����◾|�7�n�K_~��W�Y�f���䒋g͚������N��h�b��k��^���ض=}����;/������`����?~�q�765Q=LT.UBf�Y�����?|���A��r�	��ԧd���g�<��g�r�WPkڲe/?���}��w�w���	������?��ө����~��B�/;�E�q������g�}FS���J�񫮸���C7u۰}i��')!�P=ҵE�b^�O�ϼ�x� E�Ѩ�����t�����O����=�?{����������~���_w��WV\|�9�&���C>Nem�:�|���2Y��s}߼��O.����?^*#-~Ḧ!r�q���=Q5X<q��B���j��И:T�.A_�;���u��e�F�G�[�G�G�dLk���볘�5F�bQ��5�IS�L�-l��*m���"!`ܝ#�=��P%�<.�$�B݁��wC�=�+Wmxy�kű��т`PP.v���$�JܞAm�4�._�rӺ��6:��R^�S���!��!��*p�&�z8�9��$
%��3y�C�d	���P��H�R���x���^X���mJCcgql|��ɏ?��o~y��_�T��)Q܎�h�V){�Ȉ0���6m23y�2ե��bp݊��m�P�U+�F�~�����ݷ��c��?w�g.��P�ͮEBW��U5��l��b�D'p��� ��K��qG��)U��3�k�F��M�G5c�n��g�lu�/��Ɔ�GO=z��M�)��9G�xאM�F�����?a㦍���Gu�)��
��;��ܹ�Z������_�<udd�����ү^V*������>��_���^�ݯ~��w�qǓO>j옣��7�eI�����_q��{��q��i��~����o�t�Mp��|�3M��|����G	c����0e���o���/�w��G���$c�?��=�ȉ'����z���{���O;��7��ˏ�>����6�����+�{H�uk7��_~��@b���?<��#��u��5�֮Y��}h�ԩ��ݜ�T~�b�>Rv.��B�@�Hw��d��7����v��TݴԊ��v�����>��Ck߼5|���S'���߸y[�e��&Mj��\�f�Y���{�6��P�\LY��m�	�	*���"��<�*J�C�NijT�1J�-*2�߬IT���"�y���iGG�3�<���];ޜ��>3�)���H{0�ŵ��/L�1��{饗̟7���c����#U,�k��~���<���$�
o�Y��w�V�oyhp �Cm�`�$�!<�x�vǟ�S��T�JN�d�"H�DIY�D5�?�ѭ2ࣛ�UR	ʲoI�/B�4�;��T�r*U郜�+��Zq���-��N�ztNi8���rY"�,���(f�κ�?z豓O8���ظaݣ}��k�؈�B]`;V��*E�0{u��m�}t�=�d�����Ks�X+TQ�r#���ޱ_��o\�1��ꪧ����HZU��=�����o��u�wh"�:`H-(Q�Jf�E ����i�����0��JEda�f��u��1���l�j�t�5�~6Կ�wO���Eg�3>�(
{�~Ʈc��"C�$7n�8}���~���;N�� btxV�˥�^z)�J�&��ʫ�:��C_{�5�P��tC�P��d6���G>�����k�t��9���w�>/~��߽����,���hJ��4x�+_���448��/���_O��^xe�
XӦMۼy38���{ﴙ3��\��O8��%O�+_�#wuuQ�������SO-;Α>r�9s�/_w���E�}���>#����Ti/W�d��T�TRO�f�9��u,�]W�tJ�`,�U��Z�;�Z*ee��5`>��#�9r6<�痾p��_]������X�gL�Gҧ��b�� dc##`<��4��c�����$H��ӹ�|P`!Ʃ��ʩ��_<1�
�pZF�Tʆmc�i�2N֛4p1�k*�%K��xe�a�4GI���༲�.�xXu�����J϶��n�vF12p����!�-��I+�_t�V�oy�G(�����q 2,�03���j@�<Z0 ��B?;%C0w/�#���S
(jA�s�9F2�P#����N�V�.�:"2�,���dR� ��`�a�d�ҍ�<��S�������W?����ۦM���O|��?��S���R�K�D	�����<�+Ղ�]��7p$vA���ɰ�.�[z�+[���{?���r�T}����:�B�J_����}��kt#�QTM��h����#]�r�|el�\�k�l�z^٭��ّqgpX[�҆(jb,%�t�BȺ�����GDc�᩻NW�֫�������D��@p��֬}uū,�zPMz/�<��Z�v�y�D3g�x��'f͚%)?@ �y�X����j����l�a��būg�y&��H����A^�|_�+��m��=��|��I�n��-C����9��k�����@��喖������FɫP���9��Cy��?���g�}F*�A8>(9P��;v0�ޛ~�=�p$ s�
�8�C��D�&GI&!��w��K�� ��A˔�3:6��Ɔ˷�vO�;�_��?��o�SN;1
��I셗���Ҭ:����a:::���J�rsKSql��K�R%�k��}�(��~�DK�S������Dƙ$4�/fr��`�CӶT�Ƒ�� ��}��4�N�(�����L3Ʈ��M�`/`Q��t*
��>5@h��glw�p�xSC&�h�V+��)�|��n��>6a�H�c܊"�A��!$ؾZ��������D�������B��U���#x3O�wPY��!i���b��,���<������Ʀ�/��fۦ�%����3��oz�ɧz׾��z{�rbzn*�e�h�r�F�f�V?��#һTk��|ta�\a{r�S����;�Tr�26��B��k�W.>���n���"����dPE<3�nkV��f���o�\C:N�nhds-�ܿlx�pzʤPѩ���ȁ�pmc�uء�o._cت��4���p�QՈ��
<�خ�1�JE��I�&576��v�E=jT���ao_o:���u���=��%�L֞���+��:���~��w����љN���bۖ�L��0LM��������	O�ե+3�xک����ﺫ��ᨣ����/ǲÈBp���6uٲez�޶uh��3fA�y� |� 7�P,�}�]��=���'�z
�`kk�7ި���h�~���iᡇ����I�$�����z�,��Z�o>��S�_~�US���\�ɯ^��-�������<�7�}}.<�ڡ���ѾO괌iM�h���۶iKcS��Xh��e!�HEb�P���~
IES간3O�G��#���@M���;z@�e3)�i��^�+!�D��\�(S��>(�-��*������6��X!F��w�
�c�"|[#)�&آ�Ll�r�bW=VAC���Dݢj�MT��%?���dh�U�eK^�H⺰{K����Q526*��>02C-���8�4�]��B��5�7�������e��;�p�ŝ3ׯ�v�eW���>}�	ܾ}sSK~d�O]%D)(M��U#��^l�<����H�Q���P� _��A�E��=�=�ީ��ϝ�#���##p3:O��ϼ��^ze�z���x�C�u�o�R�=���3~��G���#�f�w����6]D���܁��z���h�k���6�mK(�Y}+��_ꊮ�l
�3��)�.��] ��S���O|��]z)6���O0�h���A��Q)-�OI%{<� O���/|�^{����y>X5�li�b�_������ׯ����:h�Tp�Yk{��{��.Oq��9��|˕W^��Ca��J�lvdd��\x�)'�w��p������a�_3��m�6n�� x~+W�t���p|j�-\�p�ܹ𧶶6��5�]=�d��2q��w�����G���T�e�_�5������?�9�mY�3f�����Ǌ�|��_:��_�伌ّM��٬�Vn��Ӿ�K�Z�Bq�ʼt��'ߐ�JE�L,1��J���✝�T�OQy"5d&��b۶m�<�~�`�aYqRm��A�@<�D�+"�/��'��*I��x����O!Ry˒����R�q~�nE�O^��Ep�!���˯���K���
AG�q! ��Sw��^J&�`��ۻ��X���u�����_����ؾƏ(���#�! �a�R���m������KW���}$F�JrP�qWt�֯]=mڤɝM�Û��oڡG�V��Ozo:�o�]��C;�cW�2��;���X���y�LiK�-D�)į�{�r�� D��ڼs�p��<�y���|��/.^�h� <"�8��.ƙn|��_��?���J?ʈ����L�kQ�{��镶.vҩ�D|��t[f�����ޭ���G,n]DS�
e�8��k�>��oA��@�h1�H]�T�U��%�]��t�ۓ~M][5Gũ�2>L�����;w���?�8h��e5�����X)�K�1�7���888:~m�h��>�O�:lhh?���l&n���9|�� ��%�v��{��]]%��y~�X�4��\��������~�/4n���M--�����t���_���O:�;���m������[��旿�e�S7��<���ϛ:y�M�@�^��K�Y|����{�9'�rJ Ĵ�?��3z��fM����Q䁫B�OuZ���0!�&��f��&ۊ�?���F�8�x����N�����G���(��ᐿ\��\49�oRg��.ث�����f�����K�=/�ZX0�DA�,�҆i'O5S����h�aZ�Fd�\ӑ�F�=B�m�.EWO��	�(DC���FJz��a�	��q�[�N^h�rDǀ�	:������(f��i|�� C��(;����V��{~h�.ר�A�#4�nE�����
�lAŧ��44��H��Y .;���'��y\Wy-.*(*d=J丁�B�d� 1@ο[r� ��-6h�t0�f�f��=)��aI,��X�`���}l�i�P�E���)��<�p�rq���>~��SfsS����xnC.O���I�p�6Dͪ������
����'h,AHD�ЈG���y�R�J��x�w�k�dSuTK�%@�VDY���}���}Ee� �tޘ)_��mE������Ǽ\OU}����~ق���C�Vq"��r��=Z'OΩ���RQ�6|U�Ɋ"����mT����ڤRs�&6C144��3>y˭��������b۾u8R�I�q�u~��E��O�F��{��~��w�q�S�T*�bQ�t�gDJbHB(���ϙ3g���?���𢭽-�o���M���=ݰ:F��L��m���s�����g��̛�����G��o���%ǁ�Κ5���wӦ͠���F�����Dfp�J&������t}�)���|F�`�dv2T��?�TT���W
���Sk�L�������
䐠"(%�1���� ���%�:؁��d3HS�<��Y
�g��e)��
$K�T$X�W��n�������V�V�9��k�Τ���s��F`1�K=Q8hq#I�:�Ǹ�j�� ���������a$��nkU�:3퓷����M�M�ؕ��0v+·<�Ynj�*�.e���ر]3|tt�s�`
مJ�<B�7�iA�=-;F\�J@M���K6X@Z�x��R�T��=��S)�����@.&�v+O�2������A��*�t	s �U]�;>>����y������iinnn�2�KA��auj5��F�T�~�o�r=7��E���" �t��o��Vլ�ߗ�qK��c��e#)��<��\
��W/����	lj���qĘ�<
�y���}G�O��(�gj	�v{m�jH-���[��tm�����MU�j�8�ܫ��}�G;��ϓu�ծ�RS��f(	x�с�:���.K��͍M�tf���/������~�L&���4k��b���_�ꬳ����o����V8��d��q:� D3>�<�wX=Gu�I'���}�G�~��ߝsι�_Ke�5#b��x�{���/���	�s����\�h�}��s�a����_>��s�M�~�G�{z��{�=�C���A��G������8@���C�CY}�/�&�;o��i��:C>L%W+m��:�(�3����u,�򙢃�j�
v_ /I�1؋X�ŤF�z�^�D�9e1]��S���U)uM5Q�jUar�����t�@wal��V��O��UJ���bA��z�N�;MILD%�ˌ�.�Kj{�	�q����zc�"|ˣ�5�	��I!5�M����epAM�_�	c�:��Jh��>/�^Pͯw��U[��!��\��ؖeS��D�$,DR*���W��1!Ia���+\I"�j"�BU�P�j8"��	t��2uK��톓544͜6�������.s��1��9e��+[���jV#C����%>�*��,|T#�v�E�����+[E�Q�y���ώ[ʦ��͆w-����X�Z�%����M��l֬�b���8a��๬X��p��ӳ� ��p��)]*5]��|���;�F��[��ք����F�VGgg��3�ԥ�^
z����ُ�>������<ࡇ������?����c�w��\w�u������g�]�vh?�o\t�G��O9����<��cO<�č�6���~��?�䓚���Edj](�~�����;唓�Q�җ�T(��~@���N�����);�}�:P���η�L����}WޅJ��;��(�0�JF��霷��ԛ[Z�=���.����o^�"L�C�x}!#e.���?��'�qBUń`_�e���$$�#OB�TkP�<���Q1����F(�`����I��<)մ:��$�Z�7�ar]�>^(�H�R$2a�S�����dP�~���9��D��U)�$s�����A���9D>�����J��p=�p��d�l�`mI�sl�"�=�xHR�H�nQ�)d�@e���gׂ�=�u�$
� B�Z����j�l��3��0�$d4X�n���W�1�#�l��uǘk�
��Y�\�� �eCC5*�@b+����7v&�H�'Y�JxFQ�p�\�S�^�q�p;���U���(лH^����;��V�M���\hs��$�ٵ�l�B*Ȣ��Ը�,������?�cX�|��sGQZx�t�����'��U+��^�+"K?�|�]�56V7m�,�&����Ǟx���J�ȷ�T�|�%��_|�Q��7w�8��R+iNZ��h����&�ʊE�SQ���Ȭ������(�.���z8�D�Y'��?����p_�r)�Ͽ�F��Ax�W֯=��o����wB���^M�����|aP�'�������,��2W+�/�M��?�0\C�)͜9s�ڵ�����
����?���Pap����}
� $����Y~��SO��
9b:�wVS��J��24-�B�r�M�p�O?i<��.Z0�Ưk�����[5��
�^�6��a��'-)�b).¡N�iq�E�R)P��*&�����z,ݐ%��5� 텚a$ �p�����RV�)��3;�ɺ�E��j��+
TY��V*�.�G$ʐ�K��A����i����6�f���;�C6�1u6�Y���`���T����HuK��w�:ܭ����z�D<0u`` ~��l��� �*H?���՜��<-e&�c�4��t$�g��٧4���1%l�j�9kV{{�x����#Y�[@^]��N6�H�P��=ߎ�~���"��y�	0BU�/����x/>�?]ǦD�B?����Ƣ�kh?�dŦ�=J`{�bؔ���Q�l>��%�8"sĸO��h
�T,:�n�͟�Ϙ�55�D��F�����):%D���$�[0wv����I�K�qw� r{��M=����M�To��:žKS��Y��\bޒ���Y�HϘN6�
l��Ү��L������S���i-�}]�fW�e5]Wa��i�zl�������G�ʚ��E����A�����&p�:�;_V�~�{Xƍ��[�®k>U��x�'foD9���7�Q5�=�/n� 63-�Q$����`��2x⎃�k����)��1���·P��
��i����r�:`���K����G������u�������݃�S��f5�ؒC(u�jIn �U�S��w+·<��E�T��
�˟��㗞vɌ3�4:4<^�Q�NK<J�]j9�� ��x40.��`gdә�W�5>>����kb��*q��j�(��������	�F�E�{؟��	��x�	�s�0��@&���'�n�r���R�§�V؊���Z+��Pك��,*��]Oq
B�K%6b�����C�Z�_��6uY֨�u��	�<V��DI��N
rLg����43Q�x��+S��TJ��{bv*2MOyV��T_,��h����P��
}���\5^w�1F&���	L�u��˚��ɏBP�"��D����_�[�k�ة�j9Տ�y5�9���Nj�'e,#����l}�u���
\P�-�� &B"�T�$��AڊG�KX8���V��qcAm�PW�+�%�7��7�`��*ǼС!��e1X&�W}�����|A�2�r�u�y{��\&3�iCCD?D0��|NWy:ei\ۆ��6�I<��%���"
c#ӦO�/��+�����a�As��������T*b[��A��ũnst/Fc�=ݙƜm�-�IoL���NL�Lq�	r����sr{������(��r5��P�+o�<���E+5Gwߎ;�#���{ ���\x�sέs�i4�^,ɖl�nl0��I�pL�$@�?yy�$/ɟ��Ix����ac;��M�,YViꭧ����>�;3�G���ܽ�h�̹��귾5>����-j�!���F�T�B=���?㌷ڀ��R#��p���n�H�-$�]IA�� D.9$��*��9�n���P����4�/�C�vQs1���?��T�
ʘ��G�O�K�~�/��9�su$���.%FE�|�(	�L���<��}�*��qz�[�h��xr�!
#	$f�e��/X�__=:x�k&Fؾ'�IA�B:���f��*��""ů��BlJ�F���!�N�uD�Np�pE�lS�"m�uV�c�k/Ιd�"	�J�+F/7��N<�o1���x���%1�4I�@�W� �"��<E/K_�!x��"�Ev<u1�T缊ŗn�$G@$#Z]2W��BD^�2�B�@��csJc[<�p�}.��0��
�{�/��ӉMㄆ1M�aR}\���F���[��z�����0l5(��	�����c8�M������I����y|xx�R*U�F��n�r���}{������j����z�v��^�Z=����9��G��W�㛷ܩ�ȼ ���D�m%��Z<��b6�3��,J� �D��\��]�q�榧ss[O;m�櫯���G�������$mZ�`�}j.@�_��}���x���� ����k8;W7�e|�����(����ckS�k[�<A�c�%RW�8��G
�1ۋ�H-�6D\	���+�+J�G���(ID K�L��tJ~�F�a�����ѯ���Ja> Dz�ͤL7�"�2�)l�����0Df	$/�i|����ꊱNԜ�����}����E�C(8�uhh��9�8��@�#l�4=��
�����/�9Vp���k#��̟�c�g��ǘ� w0�� ɌS���ʆ|6���K��G� >ڒ�O�Ie�DR�wBV4��H5%Q��"V�1�gHƞ$��_��N�YGZP1�s�C��8�B��h�YJ�	?adlnP��Y����t�8�]tٙ�H�xAq�ҫ-bR�r�G��= ���)V��h*E���e2�~���1�\���N������}�6yl�5�jEtx����÷�r�g?����ß�j�����������ݏ>�ϟ������g>;::�T��ι��nٺ��_��M���S{���-o����Y��4��4ۡy�f^:.)XOt]�v4`�=xnf7!�E���	,�v(�$|����n�$i7��j��fʹ͒|���mo{�s/���ޏ}�c���xU��J$����h>;7748p��a�%�mިUd�jG�'�l:m�#/<��p^��.E�r%�oq��Ř0r�pܨ��
�իW7��<� ]�u��p�=����ȘU�ˁ���4��7���`8�S7T�O������\$V�A^� l�|�Pv���`Tև��Ч�ĉ�|�J|�(�NN~�_���d�*�k�0z�yU��7��Q�
���$�}
!�0Z���i�¯-�"��z&�b���E%��r�	�"{h��<���?�Dk�B��
�5��l\���@�>6����v?�f�ۍf��0V)? {��;~�y���C���n�H0G�i�bM��i��4��)��`�Lh
�?߼2�Þ�Pl��䨀�$��;Ӆd�5��-��J!�Xf�F�:�]�����ʭ�&f+�� � 4X��R�W2���VYp ��!����i�R�#�=�MBS�X� LoP1����/�n[���"�s�X�_����r���6�����f����կ~�/8������o_�����w�s�o�Ο��mo��׿����S�'�oش%N�sϽ��z�{v���-��~�_��M����{ff�ӟ��_�Ó��D܉b� �QBj�`�pTȮ
TvQA�S�	|�,k~�n*ǔ�He��fM%O��U*۶��y�ƨ�=~�8fk�ʭG q�	�hxdx��Uł�q�&���3��T;Bvb=�����X��]�}#���t�^�e��<�9Ӷ�p��gWJ��?�җ~�?���96�#��Yl��Y*�@�{�Ns�Y�C������v����A�2�����ģ�!~_P�a�=Ӎpk�h�Q��@,�xÍ�����u���}�w�(����C�2��h�йP��R���ٵ8�-�Pb���6E�Ⱦ�V�l
�hŎ �@����d7�8��aP3{5D�Ұ2P�?tx���]�M��S�����{���Κ�G�a��=8(�����3�ع}[�V����G��+���4�8�m5�\`�DP�DiBv``�F�od�[���^�ӂ&~�<�!P�7�S"-�u���h��ゥ��HN���O�F�5	]@��)B��������hΚFZ�3�d��Gh��"�Z�b�RшGA��Ʃ���$�pb\z�B�^�)
i{q�B�B�@jg�1/�q��
��B�Dy�}�>�K׼�C��.{�E/��v����/��E�𡱕�##l�������������gl;W��_���w=<>��ɽi�tbc���Ax�y�y!�G��\��
�I�Ĭ����ϭVJC�V_��ˮ��Ʀ���B9P�fq���3�2��3�?��ٺe˱#��~����Ч>@��A���I�|e��}��a��p�B��Dm�Z}���^r=??;;=C�Q��L��<�A#Q!�_��W�3��sv�y�լ�Dy&P�"�+��������&,�Y�x$(���pT7�ַ�U�/��Ƒ�ĸ��E��9���n���K�����*s|��]���^t��M�)�;�R
��R���x�i�����<w�T:�h��qbE��Uc*������5XZ�D�:b�=T*6G+[׏���q�LN�z��o}�Fs�N��k�E��.ƺ�G��������P��n��$	No�s�GB��FY(E(��(�P�u84^�����Tҏ��hXhKm�NƼ��>"j������K�.���$�,c'�tcA����;'J�&駨%�+����Xt�¶��sw����7�CY�MC@�=�~�Bf�4�\�.C���e��p+0�n�������/���?V+�kW��u���5��ؾm��w���K/����eo��=7�����7�ر�V�&�������(�6[Qea��ƪ�
qĞ_ �����a<�}k��
�����@� ��ǥ��Q��#왞b	���G����u�7�y��aX���x��r�L���v�)&��n�j����_��k_ٰf��_�z���Ȅ��2Jw�5D�����A&p�ă��%ȇ+������H9�1E���p�߇�d`~1�.>v���N��_>��>*��)Hl��>7[�xP��d�<��0�-���i�`WѰ(�m.#���sA��e  �8I���HƄ�u�]�6n��_~����}{������S��G����4P-�·c�q�[I��B��CЩN��Y�2�mb(�$0���xU8	ҍ0y84��*;w�u����1{��EO5�9���h�����w�˯�tr��pY��jϞ'��;:]*�CG���Z?���.��_�+t�V��D0: ���)�*��+;~��������j{&��Ȕ#�1�LIX��T�Єλ��p��f@�d[��a�ؖ5[X�����֘Y��%�DV���-��(:?�`�f�GB���P�׼�X���ZkA�#����!��m�Xp1��/��Ә<4��?��`��OR%�ꄬ���:��q�g���_����x�~�/*�B�,%�����?�W^��O�����>�{ߚ�UC5sٛ6m^$��=�g�ƍ��A�M&V��x~�\�I1��y��N�>x�f�)No���8�*�]s�+
|�C`݃+X�dz�MM`���0����M���_���B�)>���{衇8�р��=�@�j�ڭ�HY�ȳ�F��*��?���)K�ڨ߆Y�_FQ��nf���.a&A<�n���߇-Y�)������.VȪ ��
�Y��V�X)W�����17��0���|j�\��Pj"�EAc]����8^T+
��]�����w�#(����o�]����y�9g��n�>�����BC�8����4W���l�$���r4TX���c��~��.ӌ�RB@�����WM���y�]7�t��vt1�Ƣ���a�~���/=���RQ����m���=�;aì�N{>`Q����J~�����y�n�VD�9�#�"in)�O��5IUs���Ν�v�����0Ʊ� ��`dZ��a��4Yy�!�����1T��p��^P��!�! T�{Ο��b�$C���K�r։�A�8$�2w��b#��/Q쭴^�"���#�V�t�#�ž�e�d侐�	��p�0�	���_?�f����<&j� �5V�����������_�ʅ�����ox�/�d�{���_��_���=묝Gy���?p�cǏ���ox��޹gx^����-��
��mc�v���fI'l��M�h �@��s�6l`GB�8�!�^
z 9Bdh)ޙD���<i%���-��px#��ῠv��X�l*���Lfݨ��K�3Y�X������P�є��-R��q����N8& m������m۶���;����9�2�=pKr�U#�Ÿl�![��m�d2�Ų1I��,��sY1�6N"`� \%u�I,r���0�0#�θ)�B8�d�jՁ������z�g���W�j�ѧ>�����%_����nZ;:::;uT��f6%�N��Pl6tvs�i���#'Y^��(!M��I�3�d���;��۶'B$j�G�*�2�Ј~��w�.���� #R�)�j���.{^�].{��c�gl\���l9�j���c��񹤣t���g&�@�Ma��
^YT,6¤����^���ۍ@�)��yfO��[��iF�,�:�}7���A(�(޵R]�'|*���l�)2�)c����D�t)�����Xb[�%�#���	�J�"�#�;^�!(g��gD˓�V���š��o���ifA-ږ���ɝ�1��փ��T��	Xa�l%�=a)�uR��}2�|�_�S͹#c�#�~כ>�g��C�vl;��w�7�������؞�����6�����7<��/���� 8�3^���q�mo�擟������o���5�Ҋ�*S�m�Bl�$2F+1A����em�!��|��B�/�St����V �]�^����q[�GG��l�>� ��W�0Rl��Q�9��%� D2e�+��Txv�N嵣h��ͥb�Î���Jl�?>��)KC,@U5ͷ������c��(N%m�2O���L������A�8�A�1`���<�y 
ƓA�4�f��ر��t��ə�j	/��U��~�^�����vໃ���PàZ��f�\i�xh�x�={�\��_r�URx���7\��n���ɿ���۷oúU;�<k�X��F�1m��$�$a1 �a¸F��v+4Q�W^�
g��Ө���dq��
k6f̭p��D���W^)���b���1�ڪ]���V�4�����g�1�8�C�4N�|�T,����ER�����ʂGA���=-Ԍ��OR-���Ɔ�9t�(�K�h�}v C���d���o1�dAѱ'�z�!���2L8 |C�:IQ�w������^S��aǎ쁭�Ur��]Qyk���q�,��c6Tb�9��d��������)�%c��P��m@u�o��_{��mB��Y?�q�؟�����`�Ng��a�m�����o�g*W\�|�ǜg~~vllt�ؤ��k���?ܬϙXJ%�Qkf|��˚�����c� ���,)5J�bh�4������)��U����$��q[��B
�$�Rt�^7[�[)�I���Yv1�#zڱ�I(l�54�,z������� Z9������S��(��3O��&�suW}�xf��f��0�R�W� yH�0�а�0	��G�B&bVj��j���3�:c͚��#zd�����˦@������izb�6Xm��ؖn�!�Oa�hv�o.�X�+FO��<�h�Ī^zi�6d�O��3S����N��?�s�����D瞻�P��vl.�V6W-�� ���T�|>t������(��bh^�4��Ih:̫m'8C�� �Zb)m8T^���&T�Ո=	�6ϖ�;� ��W�}�"��p��D(�{��*߂�(�f>*`�0�&�����`�0�	�֑����%���B�&�S�q�ph�au2-���Q���\2;{�(Gs���3&NT�ϯ[�������(	�����'��M�w���Y
��/�4�����4-�Z@J���7;0��tT�i�Jaؿoj�8�fks��������ЊrQL�LW�`�1V�J$��r�@�I-s,�N��K��4��E�<t�W�i	�=�vb����m^�o�(�|������Y�j���A�Q}�C&ټ���v��Pq�
��n�����k���2	��r9� �C� Q�:���k�/Ȣg��KX1�5BK��5�:+<y?:6v�y��{���G:q+��6c�T�8�x�8����T�	���b�ln9��F�%+#qC/#P-��bɼ���C��+`?����8Cxʒ�̔j��mZ��4A��Ͼ�駟�=�3��|P�f�_:4Z&��3$�3^"����-���Ay�6�nxt㊱�F�����	1���	,`>yJ���<t��|�a�F�)9�_��Ev(8 .5���"�E�%��B�P��3�bbth�����8���
�!�v�و?(��)m���yɠ}�=�����",@g�5D,xO���>7��Iہs� jQ���O����X�h��۱��X,4�w�$�l���wݔo��Eֺ�5���3�>�T)�lo¸!I��v���p���j�7��xj+��k�.Z` {��YS
���tX�NѰ��]��,��̅��N::�#��c�C�P�z�U;�a�2b�0��j��w��573�j����&�<�ʱN'���>~�y��+'J�e�Q�6y
"%�N;-N��˩-�,�iZ��`P/�{�� ���f�>ĺ�U�m��je�G��|�p���ӈ3_���,Q�53;CBځـf�o%��OH�F*����`�X��ֱ�TJ`���p�tΥ��H���&.���J��AcAm��)h`>}�Mk�����GiV��Ȉ����}{��F�Y�j�,��r�<p`��W\u�7n���hHY,�Eq�g�?��)�-�P}���0/Tq`,Juemt�J^k���p:����`�\�~��+� �C�'��~q�Ƽ3s\�۝�7�8����{D���X�,��TG֮�ԉ;�Fø�	��Q��0XMn�c``pt��c�
�Ay@�>pdޗE��¸��?M|c�M�LU�WU�2 ӡ��"Ϲ�FJw�'z�:�GH7���s�Th��r��T���O��G��3xj_��{�Ke���,�vE����F�`��1�/��`�]�����G0���EI$ BKm�}\�ڭB8o���+�F������{����j�D���Q�e(����!�������P���ZtMI�Uw�;d'��2	<]���5ٌ����;Oz�a�4�s3��F�T6o9�W��U�n����j��}���v?��2������(y���j��h��` ��i���,�30��Ќ
O�0�Y������jH�(��9�d?=�7Q�cǆ��[�vmp��֔D�N|�EZ���l|ǝ�r����M@ El���7������<�G�$R3in�4p�,���c��7!���0Z=9���WoX�b8D�n�\��
S�<��ck���3u�����|l	�Ը�*�a���}�|Q�TWՆTw&<b-�6M��zvG��	��-�Wo����Q|�s;�Y;���q����dd��[��&;qt����S���ܱ��X
��G�F[ŝ�CO]�P���;<}p��-O<�j�j�`"E>nN^*����0���|@_F),-|X�OcXZ��Q'4I1%�~�>.Kϡ͓S��>bYA+�<�;���DxRB�rM��n�$���SPm-� #ɸ&�5�����,b���9|�@�#V{M>5"�:�z�e�G�
a�b8;2\.W�!U�~�'�|�#=t�ȡr!* �	:a�zb���+FP�6^ ����ߦP@��s��)�����Q��8jp��yŉ��e�ՊB"�@�^��V��+0�
�" ��;a�H�d||�T��ַ���+^�yPK��x_T%e?$Y�wNzdχ�)b)O���D}Yn����N��J�xT�~0d?=b����СN���.�=�r������J�<C/�-4߅��tQ���m���_��׿�%/����\'/0�w�ހ�⣇
Em�m�	ۭvP*�]f�@�@��Y��J@�=a�O�j&��/u� M@iL��ݜ��,�]�D�P�d��*ڸy�	�̮$Έ���(�����{�%�s3�f��̀Nz��|�N��'��ЀAbT0c��|a��`�Z�T�hyR��St�Uy�&",���a�9������s���b��#�S�9���~Pb2گ���Z9Q���_{5W�#F�B�hn���5�����ӂ���z�G���D�_/R[�4G".�S|��_]L�L� R5�o�ӒԆb����gs0o6)�J�RP,#AR,''���K�"�w�e2��r|�S���+�B�E l�$�Cj,sX;��8E�G����Y���@�T���T4�Zu`~~>Q��n�oxd�Tm4[�J�_
8��:{O�T�3Y��uK�i�����_u���|o��B�hT��9�1GOMNS�i��Ou֬,�BPH�8艍!�ؙ�?���,	h����\�6!u50��w�W2��ᡡ���hd�4bZ�W�C���X��^��Ӊ����~�e//�q;,@!J���Y��̲|��5�uO�Ts��f�G���/s�8���u�7?��9����6.b�I	@eh�7Ѡ\�f�����FW 	"��H�\H������j���|U ���B�[m0q��9��r�<��V�m���4���7'�E��AK��tat@�Ƙ�2%�3���D�P�q��TE���0k$J�Q�ah�Iw8D9�}n�1E��F�x�-�LX�'�?� Z��
��5Q�L���r���"��d�T<eAL!*q$�~�O���֍9�b�M"X6v�NP���{8Z��RN�a)6O`��l�]a��qa�G��XPfЈۦQl�����|�,�+�$�ڞ����[4�i��7C��Q	pxCw^���V�X100����l�G� ��j#+fg�'���)w塧�#U1to��(�Fc��Ag4Q�13�6���Ȉ��
0��f���L]kF�UF����j��Y�=����y�CC/��̘�X)�Rrb�O#Xп��i��؆�U/|����-�E�s|܂|�DU�U̓�.��&��f5b�r;A�=��v
���m[���2��|L6��[0��D�5��Ӊ�{Q*����Jv����:����������ÇO۶��;؉��e��2~���� ��C����A*�Z{�/?69e,J$1�F�݁]�2�h7�jxdЬR��!�	[D�
m,Fd���\44U�+�=J@��ԮDEK���
����H,�+�.�	�Z�����	��A&`�Z�OL��$��s��֭ی�kuZ��P?eɥa���W��=%"A8l�D[�� j��D*��� �F��ø��Rأ�V}�58�I	0��(jWk��Z�V���2�P������¶������U�+�D�������"B�Cx���J���Ty��N�t�o��$pc+t,�;U5��h�؄b�� ZNo���A	����Tk|W5�l�L��4X�T���ou��������?63=7�bdpdE�T(����n�Q;�`������!",�%�R�oF����塡�R�,��uc��=3O?����^|֙[��xr��r���HE==�n��p���3w��=���v��m���kW�E*�Y�wSݶ
A5�l"_��_J�����<��}�����J&p-v�#4��X*�r�p��B#)�q X �n�@�R����K������4ː>0B{B�o��gf�C��f�"L���v��kn�9�G�Nd�͛~��3v쀁_aǓ�n��'2����`�i��e�<s����=�+&!�Xʬ�K���q��#S�k5֘�иP���U�����j��V��-x�:�k`����䱦G�Mf���>�f�����02�bI�ł���8�EH殐�\`'3����1z��YV�⌸ ��B�F��+F��x�����W�!<5)�C!ȏȔFљJ���i�"6�A�A�D3��$N&�HF4�N��H��k�'8![�T���� P=�� c���@��h��	3�K�s��O�Sy�H��<�t
�`S'�i	h���#�^j��L_�`e�ȹ�z!0�Iǘ�2��PK�+�� Vȷ�1og�V��(��PE4��!�"�ff�����={^u�+_�W�\������ǎ�_������?���7�|�����ֶ�����>�oz��a��q�����+W��[��Tv���w}�K_���;~�g~�.�袋����O�O~�߯��s���G�W���:�ܭw�s��>{Q4�j��͓���|�P����'��>��;7�_{����6��K^��+//W|L �?@���4E3;oA�(YP�<�j�أ��խV���b�b;��>� Z���������
1�Q x�]�s0�̻�H!�6]
�L�%�r��Y-����+eXKa��e_�.E��H���U��2FtjvZ���'5��i��F�uV�?mF��q*���(���VJy�R?~FOgN;NU�^(�jF��P�/ ��@ B+�8c6�_,��yA$�Ľ &V{���'���Y+3_��P*�Z����GD�i�OE�5e` �!���"sv�-�����"��@�
����͏�8C�,ɶ�QLx�82�V^d|*�2^�#C��{��XR��X3'�i�@-�����&�>0��Grx���.��N�H	YD>��r��V��#����b�2�
���ͅJc&�`")Kcv �h *���nд�Q��A/x�Y��єb����t��w>z�s~Qx�&̅��������t͞���ц)�b�)���&\�8�fǷ�s�k_��:���.��;\ܲ��	ܫG��o��߃ɦZ�x�-�]wӺ5�/>m��L����}��G<wp+V�%�L��O��3���?��[n��������+^�����>��ۮ��7nZw�M����G���t��w��]>�4�=O>���׼��Ǧ��*����Uk���'޽b|�Yo|�3���O]�z������9F���#Wu�!҇�C����I57T(Dz.��^1��:�M-#�&��Bn4��v�۬�*03�#�S�M̌D��?n&���ԑ+�M�)-C���iC�+�� o�� d����g�t� ($�4����z�����X�"�\���p3�w�Z�Z����ټ%ً��z�H�2<�dsQ�e�?=��ˠːaN�O��鴛�R�Ӊ"$�-��3Ȟ14�`���`"T%�I����T��	����B�o5;�|hb�ʉ�	�h�@��j"�g��_Hu	 2x�UG�Y�nWh�Ehq9[�fn��gD#����!��2���\D�d�p�����t+l���4��V��*Eċ3�b�pb�"�6F5%q�.���y0'�9�Ua΄�����N?b�U��AT(��M�����݅�V>4�U@�;B��B&�Yh 򆒍��q�;���,���:��2�����e?5�~�����u󹗼�R�>6]*U�OBjQP��k��#I�@�@�,��0T�S���S<��Y��bL���?v�Xk�x43��U6<��R���gˀu:lժ���������vڍ�}��+���H\��h�8��
=��w�y�Z��<�>�駞>��ZZӭq�h��niܭ	���q��=4��Cpw���!x`g}W�/௣�hԬ�Y�)�Ϳ��9�7cy�w>Ӷ�3�]-���I�Ǎx�J������n�N�Eߡ�?|�K��o�VOOLO��M�j�����C�n��z��I1(U��X*��i��o�,IQ��p��/Lh�Q�(:��l�ŏ[��f.�x��l0p�}#0=j8&p���7�>���?&�5ib�\��b c|0����cZ�?r�-��̓$��%��g4rt$��Z)�q����.����,��p�s.�ǲ�,ROճ�"|��������WhO!�٦6��F�ć��x�A��Pqb&��l �L� >_9B���cA9:lj���^��ٝR��1��� -��L�J��I7�+v�|��Ft |"��R�5�ؚN�B��{_�%�.f�Oqk��X��6������?	RW�O��h��Y#�³%���"��C�pnla�V����j��͘.`����ƕ��k-�i�о�C6�_r�	Ã��Ϯ��Y�1�C�e���� ���ڧ�{zUAu�����G�/�"˦9��'� Cq�����`}"m�R^G�h����H��8�	������f���ԧ���לU�ն������(����Oh1�k��oS���˭u���>�5�^��^��2�pd&��Y���荄���'�7�g$�����b�~7Z��Y�<�ѿ��8	�K��o%E泳���a%�Ν��������o���b�s�\癬���{?������,Kh�Y�S���|�bI�8).ԆU�����"����j���,�� ��^2YA}�<�)�=2��̡I�sZ�0x�:WhH�"��$�g?�d��i8�ЈRw��%���]6�0N�i*���9E
˪�|^h����i���U��^9:wDE�aKFL9��	�o�2h#?��	}9�@a�!~("���*=v�<���FK���,�F����Ǣ]p`e��I�ǈ�v�_����T�P�9���q@XZ�������M��#��ΡI% f�O�&����	_*¾�b��@��!�d��g��H����i&�%����A8�Z1'�U�$���J�^�T����B�q`UEFb��!8Ƅqt9���d���ꟕ��;����l3������T�<l��i���9[x�tQQ��u���!Dh��������z���]��_6�J��JWL[Ռ�ݵE��<)~1 ��t����<l}7l��~��W�
�18]�s5��
�Z�訨���dx��&�����V`gjQ��=�����Gc����Λ�o���f�_⹧�]�%�O�y.m&��GSs��}����g�U����N�KNX[6:\��T��}k7sQc&���[���s"��Q_<�h���������Ӧa���Y�9�A'6�[w�����8��_=�f��Yb��Q�a?�7��H��W��ң�,�|��s�/���D�;I
 ��D3 y�8�GU�Xh�ͮ�4�LX*ؖ��H_3��K��*�7���_5؈�
�&9�B�n!H|���	���s�ې��ޑs�1sI!�)�4
�_	(<�G����:��k�D����BM�ĳ���N�������g�;*��AܗN#��P"+~�y�^R�;S_F�6�H@�YH��)W젺$��g��R,}��6�]�^+�#A�=<L�[ �6��og}5�`���g3��O��u����E�&K�!�%g{��q��JL�Ukl�c6����4z�H{�s}U�cY�@e�rE��H��G� $z2K������P�=�$����C�RK��X�T�O���)r��P�v���e����&k�k���&._@�N9*o4��}p�4�w]�ldaQ�~�N·gc���?��e�N�e��=�����?d=$��x��u�fF�܋
>���l����~�m�3�ZDB�>ٳf�<+d�jgf��(s&��M�?�4����]u\>�|�����
Hy��o�nx��=Ə���eu��?��|:�惐��e�"=�o��D�݇���P��fU0�qb�����V�(���#��k�o Qg��.�h:�k��=)έ�F鱾u�g�,�����g�9��k�B(�(H���K�9��Z����>Cx�h*ÕE#��5�Vj��%Y���aHq��|�3ǹ���d"��a.*.�����(.m���6����#(C�6�s%�ܜ2n�פ[]!*�@�9G"Q�e���T)/q��k�~�ܓ_���ނ��]���e�%-`�q/�x�J��ᜒ�@dZ ���I�-V�� `7�Y{4(Ǒ ����Q(���Y-������uSWG�׭�H�����cpT��6��,�t��ږD~��nX��бxD��&;aD��:�t+W�@hc�$C2��'����X��2�.�S0RՁ=Y:�n���r�>k�����6�J�@��1�X�65RK{nI�����E8%>���߶)U��(kG)"P�}�������4�f��;)F�H%)�[�]H���19��4i���<u�f����,�6����2�5D_���ZN2:L�%���~�����3K�^s~��]̜�`�x񫫮�i�v�uwv����@҆E<���1W�G��V�a�n���V�L��5�:P�i��[�/��e�Ox*�1�U�M��ǻ����-\���(�Ro��&p^%�k�e�m�~2_�Ж۩��xv%}` �@�v^>��H ��J��b�>Y0V�)����O�\A4i�щ[Ѓ�����|1p��#�,�"8W
��O�!
	���,ݙ�C�\����<�*��RchU�$�f	:����c���!:h{��5�.\���Gu�.D���� 2u�ADS�(Z��2�{�E'�z��F��B?K�c�A�a��
��2�z��u�I�QH�S�k���}��Yxx����{�Y�I��L	\k��,mKn��0eHOBڞF�+��g�Lv*�,�u�y�Y�A��/F-�"o���t$}R�T�)E�G^����qH�DGȿz�fz�r�BY���8�����o��u���R�6s�h�k�E��9¡�h1���V�ڝX��Z��:lW8��f�4�V	A�!P�U�Y��u���׌��[�ZT�j��r�On����#W>��N<fY��[Hq�����㺾��X�n׉VM�dI$f�����|�p�|.�n�:�3����04ђ�\��nRu�l��%��<��ʟ j��m�7a��X��5�{g��Y�v!i�˹�v�e�6ˏ"]̀S�0}D��|����1 ���;<b�t���'J�F�W�
'_.�d3.�B!<"o�������2C�+�.��)���`g�0v2�Q!-�P�Ò��a-&��� *�ܫo���M~�k���/;�z�bw�+��b�5>��1��i8�I"�Xtݱr(ު6���7ĺ?�9A�k t��#h��덌k�*C��j_}��'�ϚT�})����r�J�=*�Q�xUU�SWs�^f��>�˶��<�Ď#҉�{Re�+P#�Is���)��pg"on����|��ԋ1��vd�Z�3�u�����ʳ���e�ʡ�7�"ᄒDSY_���fn�ԁUV\NV=�_�l��G �u���&�gA$'�OҞ��j�6���b�^b�y�"lv"�+���jm���Ĉ^>p���~�.�uOôP�����EBq/^�H�0J6SVV���ޏ����9f��2�UU�/�[8ܿ=�՘Wh���s��퍞�O�/п?ԍR'�݌8z����!ON.��<��?��8�G8���k�v�g��T�\�;�E��:�6_�0]�v��;ov�6v��i�\���~��A� %� #�GY�dS�7��/W����V6l��z޳IF"U���Yql[$j�T�m2M��q�k��E�?����^��p��9�̖:X؃lX@%�C�rZ���� ѤB9�[Ȯ���2�b#��?�A}Zu�+D� ( �õ�lQ�5
��5	Qb���[B}�L��߰Q����:�B�ߒ}���|$|j�.�7lGR�`���5;~�%�W�-{�x�Sz�(���T�n�-�)6��>q���?��+����tUBS�_��r$�'���]/Uף���N��ɌO�4�`#�M_)t/�Ч�`��fuCO��`�+hL���:��߃ VH��^To�C#<��ge�r�=ɳt�uHɇ�ɚ�V�,�MBI��{����-����I�e�u��B�wZ&�����E:J]tf�ѝ���'Hu�VͲrO�G�.�q��[^���f'�?c�كݽ�C��}Ӕ������F��^"e��r���~l�s�*����"AQ:%�><��~Rً
�9��ɸ�o��:��0����|�y�x�/���7a��K�~�KSv��I펳2�ͶV^k�>���4aN`/⡜E=��}81�����AV�e��AVVE��/.oO��[�!mun�M���E6iqDr$wiW���D�uc��'Ha���#ڄiFCܟ0e�֌��G���]�uº�G2��+�љnC��ɞ�[p(2��ʜS��_
d R7����M�v�2��D!'{@��**K��n*���t��#۝�s���S��;M߅��a���S@��0�)#g�m�ـ���>_ut9��e�uSjvk�v�nT��dx5E�h����<*?��_'4���!C����K�5�>����'�8�5E��P0<���O�z�'��D����2w&�%j��D�~��I)�I�ʘ�����/!�0/��9�ID�5s+���  ��)Zs��_]��:@��O��"��XPBP�,�x��=B�R�$#EAz�;E"����̎�2c;�7-���i�0K�C�
��=�lD�z���V�a��Wї*F�k��l�<.*�����Պv�-��{@W���|DS6���W
��!���l����� n4�`�͒H���cZK�������~���-�9�J��^�߻���h���|�O� F�C�L~�(�L}����̯��m�t��gsvE_*!���+�|[��F� ��������d�LF|;���X���G��'������̎�!5���z��;�u��`�Uߙ�(M`���0䰰��-��f����y�m8�#���'@���/0^M�c��<�d�ȑ|���B���#pS���\�+�s�ŭ�?ig+hp�pw>���2���҅�"�$��'�~�8�ܸ��4�-��?��G,��j�Ad�)�����('i�a͛c;��W'�G���~aK"?V1�B��MpuO �^��uz���˲c�|.�qr�D�"���<�vB\8��x��8l�������_�@�=��WF@��.K���B�V]�f��������*���E�FU$��:�Y�+!k�X7/>�Ə��!���hvn;+�ۻ��MzAHJ�j�kq ˂#x�&�	�%W6Zc�5u�쾇��E�f/zoh/�!��L�,��	^����Iǅx���9�D��a%
�	��0�E�4s���D�aeSq�:3Ra� �R�v�}�-ea�E�6iߜǥ��]^�f�^J��,*l�u�jI0c�ts��+T��#I0�l݋I�M< ^-~u�8 �G���;a?��@MwD������f�~��y�����s2ah��0 ���d�{�^TB�M�n��ɾuϤ�4���V�̳��Q���p�i�b4WݮJ�(���J���X�hx2I�=�
:�����.1�s��PR�d�-ZK����j����Ǡ�4��Q��L*���3.^aK�?�W���wP�ّ�r���;�&SM5q���/�Ԩ��m�՘0�]������>;,;��>MDcLL�>�2Nqvi5��3��u���R[������>RV�F�Ǐ��pJ�O9t2�	Y�n��9�"�Ly��%�,�0Y\��l��S3��ݯhO���/�w��8�{��x
y�&}<����o_�ZA,���!I�S支hք0�xÿ�4�Wa`|��ȣZ,�M�k���8v�dv1Ue�t_�K^w	f)���+0�;�*��T��*�_�c�(ԝ�ke��7Jq/B�s��Ɋ,��øn�],y�����v��ǰ�Iĉ��E���)�p7��^�l�#78�����l�2JS�����|33X6����Q�H�rf1!��,�5Q�t�],��p��$W���Iz�d*��X,�(��� �jW�*���
O��F}Ħ<�a�
#��Շ�(�������s�j��t��<K�IOe�8��E�o�A
-թ�ӎ�������!�=�A��� ������&Tw�]�;���k��JP���5�P��[R�f�V�[����F�H+,���Zb����_�C!��7n!CR�_�8A�|:�Bb�9�1��}�݄7?^��kV��,�bM�aC�,?�JR�3��uz{ۀ]h�Δ1$;T��ж����ĮGs8�r&���6gqpZ���R��ue��Z�0E�8J�~L�?W��y`�nа}���PܙH�b�^Բ�s��gx �t�ѝ�g�:�Ϯ��=` %7[0a���K�^��O�_�&���)�΁C4���n'"�V9���(�2�~�����R�=)��KS�FHf�*�6�R"�q�ᾜ�0qÙ��\_3����b���G��^�k� �+C�V_X���s9ِ��η�����2+��73�48�}�%}&��eEb�墳�nTBSGS�!Ŭ��i��:H,V���p��ա�?*�Y��e�(���CFqW�؞&���P��=y�Btݓ�p�MA㗛�%D����ȂC��5}�_����*j;u��&e��%KT�$���J��m��Sd%4Qٰ[Дd $ގ�H�U�1�� �'E�Z�S��^��z����/�+��P��.흆�?
��Qݺ,���FG�}���2�\[�}.��/�s��h(������Q��m' �����'I"t�z�;�>v(8���K���۵*��L;�{H8��2����#��,P�J�P����
f�F�t��e�*�6�/,xFZɺ]�=_!b;�Y���JK�����9x���uC(���*��	�_������V+�]���Zܿ#qs����&K%N`��ԑ�4�l�h��X@�V0��LF��Z�;A��_N=J��kFշ�dЌ��_��-/�F��p�� `��`���*
T�:$�,��>�K�����!-�@�6ޯ�<��������3=!ivI�0��F�.���L$25��>'�ִEx:1ED������B'�G���^xq`�-^|�֚e�ŰD�a�
J9��C�\/~�o�qѲF���~�\��-��$��޼;E��6m����L,��9=��_B��Hd
e����k�K���8b������z�Ҭ`C�N'#c�����Y�A��ؚ LW�U Gι�c��Ʒ���#C�L��q+�D�q9HT[@D�	~����?T�+�c7�FF�m��IT:���tm���
���	����S��hN��h?��FK��OZEϏ��3� D:)�3�\��Xϑ��P=i�|�j�Ũ�� �X�\�ٯ����A����i�S�l(���6~u|�*�>�9fv�_Q��2�7mҙӔ?��C��*.���0i���^|e՘��ZJPI��}}�/0�?"ծ���G�Jϒ8 �D�� �(��Q�6~&*`�0?�<�3�..���s��>�3�0穌�)76��ph�B�9�t���]'�(hHhGR�hh������� �s����?�Cx���EH%9p��D!�ȕ(�8�R�P�xЂ���	�������fS7j@��I�D�W�#�ţ�X:ψ�Ey]U=�>_«mY�@���ڟ<1��B3�D��!������������Y�W�=G�ZUBH����|a\�=Z����\�++�%��;�����3���w��[�{�y�B۬]dT�!<C!�R�v�U=���صI�d.��|btq�׸Z�-2{�����ﱈ�#��/��c�36��j����=�_]#��T�[���S������inRy?о�mAT��㲊�I�0�Mm����}"����uJT�J�F�w���4�}���̸�����}R�
c��*+9vn+{PDs RH#���m�Z��J��V����l/`���F���nk�ucL�.n��X�F�ŗ$�����ۓ*"�0eN����z�2�R�J�'���@��	-4�n�2U�E��]��
z���dQ�W�X(ܦ�?��e��^:�<x�o|+d��&(�h;6��@.�$���]�R�Vi 
��-�����[�/�fJSh?��6�r��C�Q�x�#��2a�B�;�Ί�Y��H��\���/���/~z1�����R�օ���������:>x�
Ry�,l��R���.��D }���]���x/7F�u�TpO����+��)�L�R��DÍK��M?��:ɥ�˟�i�ɿ��*���*�A�lW�TM�,��<����05Ł���s�sD�V���"Y��� wC���z������ʜ^�h� �MûE�䎦O`���fޒD��~�j���z��<���s�%�T�S�5m�(Ija9p�.J)�(�ez��0n�-o)>��Z�gz����m!�
�F:�i�d�m˄���on�S
ǰR�B���(�z3����?�B�#���Rd��D}�ŭ�W�6�{�r��GC	d���G�C��D9O��$H�m{[�����W�M�=����F�VP*V&Z���c��*)�r?�*g�7�j�DA�J2trgf L�ȋSL[y�5�6��q�����K`�,�X���kӿ�㡬�*61��!����uN}���ڸ�M�5�XK���T)����3�8�Z���T�2�K/Uv�]��t�+�W?y���17a1��eP�o9�
E�29"}-����Xr)�z�*�^oI�z\�ao|a�b�c|m��7z����,��V�ϼ�_�	*�oӀ����ї�R��Gc<j�S��ߘG������v���`�)�eqЇ{�����.��4����Q��+��Д�E<Va	�iy��&�H�O>��-b���
�,f�1��X�i�4ƾ�L��1p�9~�[O!��m$���,����z3ŊH�	B�P� ˇ�+��le�Ӂ��X�׾(ud����K2�v��-
���
��!x��:�6�!�2�ܻ����:8�fX�<NJ;�����jk�h6�M]��8���cqDxG�5��rI���P��˧ি � �T%�ׯ�f�x�Iw�O�KVbx
ymO�~l���o@.4�z�&0��/,����Nq��o���?�g�� zq;׈�h<z�]�������������M\!���E`��#��c��T����f�H�����(�OC������O��K�)��j϶��/�U�~ MB�PK   �m�X��
��� � /   images/728f499b-3713-4da6-8795-3b437d35f612.png 6@ɿ�PNG

   IHDR  Y  �   �ZN�   gAMA  ���a   	pHYs  t  t�fx   ]tEXtSnipMetadata {"clipPoints":[{"x":0,"y":0},{"x":858,"y":0},{"x":858,"y":422},{"x":0,"y":422}]}��U�  ��IDATx�佉vɑ-h�a%��E�����꧞���9�{�R�U,n �#���{��#U��o4���	0���nnv�m޴}���RN�_�S¯��E����%�i�N�Oڏ\m_����+e�?�+�{����O����}�����>��UU���׼����@����Ux���Oɮ�2������2�Ǘ���������p�õ��J0���2|�+��u��nφ�/���v5NL�H�����}bֆ�j��[V��$W�#�E�3d��e���?DR?TO~��:�����Ru�%����T��J�4�x-��L'�2ɐ�"��s�'#̒n��o���x��U��k���~�1z������nK~g��2/g��o����jʬ��W?��G��>DV��4up��Ԝ*}�-��^I���w,3#��k��A��hi��C�ь��2��P+��C�n�A�WRe�1&��X��Y�{��7f*���|u������x���_�o��u���;��m�������;�V��5c�F�������K����g{��it��I�����Ϸ��ǐ�������?Q0�Y_���\��k����!����+|���;e3������_���l�j��ڜ����o];���htÿ5�:�y��:3��ܧ�,��d��2b�w�O�6�W���}�_%�Е��i��Z�yD���,@��!��Σ����ikf�����L�� ($f1i@��;�� ���O�5�������N�m�b�F�ݺ]v�#o_;v0�^��Y�T�7��[7�y�a�J��x���z��xAo�ڸ���0Z�i���ץ�r�ܶ��6k���=>_��%+�#xLΣ�Y~&	e.]�Go�~�0���������[�h��=cY������5�Ð}\���h�ӭ� 6.Uݭy��(+���������.<�@�㮾�ጧC~[s�2������.5��^K$XE��f�J�:Q��;��fb4X�4���-����1S�/��l�����׿�x.�W��{���.s���T���3����_���o�M�I�w|CU%	���(~������/�TU��d�������sT'i��Û~��z5ү��:�2��2���-78^��JUQ�rQ�I���cs7ec�!�o��ݐ�������*4&D`ܶ����kdPj�S��Žs~��a
K�VU��g<U#ŝ��q������Qhs�_�:3�Y52�>_cei��ބr�ԗ�b�d�xx^���a��6".���9S�ʮ����e��x���u�����:º@��ac����F����T�� ����A=�m/�-�7�S�0�֮ϭ��sh�ڤ�-p3���o�K�8��n�m���L������~�+��*`��M*ʧ��U �n�+:�!�*F��V��G�sa������H�덪8V�\ma�<���ǧ��gFύ����޶k]��2G����=�4>�/�m��L�C�f��^���d�?c����gS���t����F�	�;m&�/���`��N6���{�t@� Tz/L�X�@�7�V���o�o�S����~���z�����M��l>Uթ�S?�u-瑟�	�P|�7�=J�(4SD流k�s<�N�
�	�o��{��z��Z��^�W�o��	����׾�6:�<�5]��z-�T�Y�.ج ��ƒ�n˨�5L����Mn��6��Z����C�Mk���7�Л�����4��tlf��=��e=�ڽ�Y��x��QY�N��� �k*��i�3g���7��������o�7ڴ-�Z�:G��j����|�<
]E|�}��t-/���ax���d��U����j^�:�oU�rX�pgz�ܪk3�Kxn�f�g8�����9BG�YF����RZy�	ޱ�v#�FO9�%e���ߡ��5�|ZO��Cf�Ɓu~�g���F��n0LcV���"��*��Zs�\�m�1[.-�V���#�Fm�G�����77�k�eff��tfg6��>�y�(C������u5�^7e9��+��ɱ�r�1�7RाS����/z3<d{���e�v_�fd�PV��x��1*�)ckx˸���_/�n�g�*�3'�wo����?ĳ�.������l�����AO��ha�{m͠��<=�z�:�ƅy���xB�j�BOT��,T���_�������6c
]2���v؇z �2i�X��j�r��5gx�l��M&�2�tK�Q�ہ�|��[�8��?s�ς��Ua\��Ѕ��aO'���?i�Sq��9;�P���h?� ��L���q@W���d���"V=�[s�F�j�eǽeɨw���9��WB>�wW
�W�������D}�G���4�Z��DI�2�y����$b_V�,�m�mt���{u4�r�8��پ]��4�G��<�I7�X�ny�9��6��6��І�">ΔV2�p.�4�zW.+e72c���{�ОT�U!�}6eJC�b ��}��4�߲i�GyW��*��,��F)WA**�XUn���y�9�el���A!� ɯ78l<U���Udq,7U�����'��U6��W�ʯ���値��h�QI[!��%c��H����/��2�){e����%=�g�zһ�:�r&U(g(�ʍ�};��\�C^nyϝK�ߤ�E��1q{��D�)����IO����~����e����c�@�$�[��I	 �lM�+���f�6�����b:�\�>.��q���lu�֍Do��M�Or��� ���@�Hua^ ��$�}����Z�^��cf�Hb�������^�n&�p��3ڹ�m��'�����ǘ�[�<1�w>��2栧.��sy�@1��2O&����ib�@���F�`�������X���kn���/��>���	߇� �4#cBmΙ��ɠ���M�T|C��lep�ޢ( � �S�T��R�fsH �m
��ovԛ8>�y�����8�2�S���a�v>�z��1��.�+Y)��T���ľ����@����'��_��|�\WN�!���9�Vei�Z���J�k�2 �����kB�F������$���4��{>�Fu}ѫR�g%3Ȅ��W�ŝ�A��ER�� �&כ�RA��E��Øj�0	H��I�@�d`�U۵��Dy��g�ҮpYUF�Ai����5��+]#���o��`��F�(+�@������*X��&w�����Ƒ
����k��7� |A�� z-֠3�P�lñx�6���s��Z������uV0���ӫ�^���2���ڕ���a�6 H||�Ҵ{e���IK����S������=�$iZW��L֚�n$�ح��;#н,�S�X���Q�B�����	Hf���'v@{���ռ���樓q���h�{:4���u��l	IK�ا&SL����QҾF��g4	����z]�)�K�2�s%�-l�H��ρd	����[�k�����3a����z�	8F�cN����..�+|�|�g�ڜ���/���b-�1\��c*�s��C��"0pҔ�vqKkΆIel�!�W��W�	��gz\k'P:]|�*^'l,f���Dd�l��)�a�}��k]��~� l�Q2�8� Se����hE�ǀ��Xn9=�W�������,�K����6AL#��NO��`�C����zaF��~D>B�/���J���h��2�b�s��k,W�p��>z���	��1����4�Pb|�*���M�o1�}�ђ�xo��R�xݦ)؟G(h��$��tE)RY91lj'&�:�@�2�1����=��q�dF	�v��.�p ��M��7���hk�M��2׃�j��T)�Ir#��2��4�c�D,����u����T�k_"Aq[<E�Ƽ=��� !I[�7~�B|�Hӳ�����!*��Tmr�ݶ.Z7p�,iD��gh��&��Wi�; 6���" "��( ��»7��o=Ҕmn�<�s�?'37�8㳈Û���>-�!����2����f��!���q��l!;����@6���u���־6�%��fc�Z_���D�۵{:3�s��+�R�?]smaqZFٌ��;�mUÜ�����B賽�"���u�����B/r�k�����l�3�l���ʄD�10�srkεҿM�#;�ϸV$)񹦳N_k�|0�S���u!�Ie2
۷٬IL6:O��B�¨��}f�&�j9G��u�/:�<�}q�0����p*쩵�����X#�ս��Y�~�uWd����Z�{�\:��p�Fw�*(�m&���('�r]Hǝ$F�jN�;�ʍ�����d�K�c��~6�o�^�h��@cQ�JX`���-t���ۧbk�M�:� t��[�ߨS�ì�g��/�/��dี�ŞX�����8���� 4 IvS���=ӽL#���4ِȘ.��V�Ъ�"�хJ��U�v �^|���,IVD1r��E7���E;���f�2Ss���X�#��vloo_ǿ��:+�o����
yż`���T�=I��u�bk-Z��?Y�T�Nu��=z�Z2z�Y ��(w�U�BFN��K%���] ���	��6�YU�`ٰ��.�I�o�j��E2,dv�d<�C�5�{�&S�s�>	N�����b���V�~�	:	�k�yf�{cJ�l���`�)�6�D��e��&�a�oY.Վ,7#�kD΁ɤ�=�i�����Ȇ�{�ۊ:���������@�W�9�+s��-�GA��ǝ�7L��nF�0O$��i���:�Y����*Nd	��sL��>�~�EeiA�]���/\o�zk�t%E��Hxp��ޘ^v����N�$���w�p�!��PRc�_�N\�K!Z�����ţ ���G`��>z-� j��Xo
25`ԁ�����"t�,�,^������m�HSߧ�J�g��t�sA	���5HT�)w����r��KcF��#�zָJ6	��F��&5�s0�����t�T��k�i˃B���}����(sc�c�>���y�aۺD�]�����%���r��ic�ʟ^����+�L*݄��n�3=@}e� [��̈����#�p6e��ez������ �JذxvR#[��n�^���Gu���g���8<����PHx�܇ǱW�[F�YQDO7%0�K�>�4���Tú��A�(�ύ�'� H�ZZ�8�5"jxV�{�'zrj\1'^�&��������	}�����=�`yjQ��~ ��{	Ol3z�ނ��w7��x���Pm]�#ˮ�D���	�$#�	Qˉ^[��5fD���\ؗޢ� m������u?��A�:��9ȏ��vS�5T�TN�1��y̌$�&�x�Y_0�;�Pg���U
�X�D`�XO[�e�;���Fܯ��JV���Ή�y�����T��2J���םE�peDk���c��ul��۶��rd`m%����0ð[Ze���(��R���HOz�M�"K���sg�{/.���N'^�W���]��k#*����S}��M�ib[~pj Х��bQ�u�!�X(4	O���m��Y딭& ]�	R��p��S����K��]g���,;ʈ9�*��s�=*�y�='M�'�h��ֲ$L)�R�m���G�N�:c�a#T��
�M�X�!�6��$A�1O�<M��KE��=��1_���D]��4���뙮��u>�� ���Y�=���Ʋ�q�5!I��ڴ%J`+�2�`�/u?!�����+;��]�rM��(P[�ޮ #�Eq�~�^]�=WԡW�\/$5 ����΁�F�1�)��sp ��ҷEv;`���N�S������[*D��Z� ���5�P1ʴ�t���%��L:s��}!�7�7��u�����m|v�߭��\,u�r ��$��YXs'̙�����,�Y��L&��u&�m:��̱c��L�-�7���ฆ�0	s�=�&�zK��J��|>#����L�K�)���`�� ����{j&R˂�H`!~���2W=��J�XjdQ�4DF���FdR����*ө�3�"�a����9����U%�+"�creN�ʯ�`��y�=�����w�!}n�cו�z�A�>��B? �d�@$dT����9�	�*����<�YId1�iI��Yd�
F�L��\!Ud�o��%|5��X�Hx3q�g�?#�v=���α�X��ĺ��O.� �̞`=���ҕ�D��ڙ�	F���q"}7G���F�RL����J�..��f%*�!+Pk���eOը
i�}��"� u�8��y8+g��B=�lA�x��$x@F(R����iՕhP`֭ �@D��AG)L��4�*�bۄ�~�4&=�;>g�"��
��Wx(��R�� Yy�-ϑ	`��9��#�J�!��O�Ј��Hn��!|u��Vi��ke�l"�gӹ��rk�d1�Y�H�7��/Lo��֜����l�9¿j�APڪ@��E0��{R:���±���Hix�� L" P�h���nd�R�j1�	�h��ޮ��$a�A�1�K��R1"Yu�ź�z(�l�0�yw�{e�)HQd�C�|x'l����d�,���!�*�Aʵ�H���)�E�LZ~���:�I�8XP�Խ�>����j{*z�G�G`�û���l�.��V�Ӻ2l�`HY��7�7�Y\�z�o66W ;��14$kH�}�fH9!hH���2%�{�[��\m�g�H
��==i�D�Q���%�%xB�ϊ�%I�H!Y�Zg6w����5=�)2	�L�Kv/a�3��@j�f�BS�h��V�v}�)�L�h��A"�J�J���`pl0Bτ
��Z�⺸/�Q�fT���w��1�>X���u�TP��!0�뾝d�+u=�cP��nX��b�l��攩s��޽�$%�2��(H��5^r'�$tC�n� �D)kg�H�úTn�x�:O�څ���:%,��؍ j����Ե���|6�$���S{j}��R�2�y��/P�y��(�Z�	:�HL]�Y̗��̈�T*˓��.皑��e�m����=�桅��辮U>��i��}hL��kH�� ú��]%�9Җ��4:� 8�j��V����5�I��e�EQc��R���t��e�7�Ӳ��Z�d�98f45�+B��Je�l���w"�nЯ��N�vE�I� B���=��j�Ys�;���vl�y���Wv���kV�?C$��:Zsrt���<�S�А5o�[&�~N�XA-"aH����Jp-�X�)h�k%Y��a�Ĉ�奁ڳ�,;�iS>���D�����fZcO`�X,�==#}7��ru}��H��#%ē�����0n=���h����憑-ڮ(1s�>K%*��&45��R����f��I���#�j�)�$\�~;d	�1���\���fW��n����m�d�z�1����u	���D����E����K��i&sx��5X�:�K�/uJm��XWfz��,����D<��x��闺&7\|b
��=�Z�$�,5I��֪��	u]�آ����������X.1��v'@��c�H���;�{#jàs�E])��H5� �N�ˌu�������-�d3�Q��5N&#�dw�Dt�=6�bZg]�"�̲�Z'm��tR�/��Zv�=�u��g�.n���^�/^ʻ�rv�m��r�-�&�lo7��ë,ԁ-5HV=����g"ZSH���-�f��ϱ���{`[3�%�G���R$������4 'qE�����"�`��1p�uFV�i7u1�ŋ���˟uf������Hu�B˧��2O�b1)���bc�7�cà6R��v_��w�H �D�u�R�TB߽y�!Le5j���3��B���0X�b����ɦ"&*#U�^��<c�x�R�v��=��A�����bg�g�{��}��� 1�S0�s�as#�E&˯R�$�Ǎhx��N�(M7���ƪ�oӔ2	��K}�����G�� ������4���#��tb��j?���9(�:7R!��|[�s�'�i��A<wȩ�p5�����+�)�J+�7�J<�8�x��&C�(ӭ\���q8}J���)SRQ<�Ϯ?��y���:�pO!cBC'R��䘯���	�8������뛕�jɰL@u��Ŝn�_Y~�U��37�S����Z.�o����&�+��T�M?�g3Rp�A�L�s8�ϵ����҄��d��H���#ɽܐ��tf�b+K�;<<��wt�;� Ui�4�ݩ���U}>��\^1�����ܰغc�P�$�!��� R�$cc*�@BO�a=O�	j6�2XR�<���Bc�����D�y������<
$w��Xm�� ��w�7���S�W9	���l4%���D*}�q�;O1�ݗs<{�D2!ԢE^�m�ZǬ2@}��N��Qץ�ό����ޛ�$�+�ĭ)���d���t YZX�����Dz�<0��:#Ő�:ى��/�m�Jj�V�����}�$���z0���aQ���Pk^��^�=+&:��Zq�h�jȗ��#۔8֧��J�g-���J��=��w�#{�ٙ1� ��>D�;�ik�&˞
�9�~��Y�|�M8�3��^nn�ryz&oN�q@��?��룮j�$�gj��������.,�;ܥ�7�������)�I�ƒuZ&��I��{cMz�� Y �h�4ԛk:ڨ�lj�CK�s����^R@��i���#���j]���cZUy}��ǃ4E�*8��¾�yUnz�������j(���$�2b�Ѭ��#��%��1���}�-`J�X-�D��um�7��A����	��1����=љ�3�܏��и, ���`_\^\r���{�m8nwOn"��MV0_��Ret]"B�|T2���t.��,QB3&d�w��� �����t�l^s����i8��cK��f��d-�x�)u���c�1���T�������6�fZt�y�M45�GA����+Β�I���M�=1����s�'�;:S%�r�:��٥|��K��_��/�迭�n��X7��jEτ�V>��ۃ�F��t��Z���@���j�yt^�3D�L�:D��o��!ԩ�LEW#�8c#�G�W��H-
�fE��
6�kt)�s�OtvJ[d*o��oM��FJ	�T)�6�5%U�x\@�$�1�($kT7ƍ[�%��hl��S���� 	�*W4C�C���%���N]������.:��o>�f���t|m ����0�,L�D��4�1�
Rr�,���Yl�����0"�]�Ec�j 1Q?D��X�4��2÷ՙo�˳�̧4�m8A������G~t�)� �e��X��vUt��k8��)C�Zԧ���*�p���Se�� �}ldt��b�ɴ]�5.��F{p ӣ(dۍ��)N��ac���%w���@��78<l^��F��*:�=U�}�P���T��,S�Zy����{�t��DnV�d��a�d���=�=!��pw.��ߑ������G��P`ݽ;�7���/���S:ȫ�h�~�Ƣ�3�ֆGz�D��K'�}�&9G�� ���$y�i����#Ll�U�e��O�����ݥ\.�$&0F���ۧ��������K}��͛wL�BvER# L� F�_O�NR���bZf�k�Z�	��2/�1��J"J�r	i��׵X.WL���Z0��iD9M� b�z�o)�f�'wsn��|�@�����,��G纁z��\ߙݠ�ځ�9.�����G:t��*�����A�7Sq��v�bցg������kѤ�}R;����d��-u+���&�ڸ�U�r+�@�۝�1B�N�=�ʌA��C�GiB�H�=��"u+7�����d�<0�X������t>4�R�DVR������Od���<���4e$
�'�f�Z׽���5� �^�����2!D�9g�dSD�֯�������$'���U�Zs
@wT!��B��[ɇ�֎"u�������5��n���O�F�X����ق���]�z�k�و�w�`#Cs�\���c��G�l�>Y�tc��,�����"Y!S�qx��h�a� ,����A�����>� 0��H4����s�wĕҐ����fD��>ZG�T���u��BFӃݑ=��}_H�ךͦ�ҷN|H���6�����)؈j�P�e�hL���g���4#}T�'h|�qg��	ÿ��7�[����F��3��y!�wx�6Q�둸fЁ�ϵ�%�n9�ǣ0�oLg���ұr+�l�9�#�j�E;B �ތ,=q,��&2��ұ�xO����;������ޡ ��D��2�7�������ݏ���9r�g|��>n4�y�F���ϣ(y �cE�2U�<�"����t �~�:4�� �f�G����L~�q�E����e�8��� �JqejD
���E��ݦ	B��(����Svͪ�@lC��MƑ���cr��^E�!l[*�5:#Z��(D�����x�^��/�pP@/��Z'Y W�@B��F14�z9�@�M2E=Ȓ}UNBj_ϊ@'��IT��_̸vb�`�,c�P~����c��2��!�҆G]�kaS�;��r�@�F��T�_d8!/D�w��X���-�<���Q��@���F.w�J*�Ĺ�z&'X�ƅ�8�ޡax����(�y��<�C�GJ눴��2�ﻁ(GS�����p�>��R���{%-]a�U�E�jw����s�kA��Ǐȝ���%C�D�W>y~&_}󍜼;���
6LS��-ݶ���H�ܝ������W�4���L���k�G�7��rrr*���/��b)Hk�)#!��,X�E�V��K���WV�U�x%!�-%���&{�ʺ=�Xհ������<{�X�=�˚��|�z(��`��NX?��=�^�ʫ7o����_��o�gÀ����!�
�٠�qm6歬͞`ݖ�ݒω����]A=�5�1вX�
C�'�mmX'�y�Hr�g����$��b{�ZZ���G�A�Pʽ��Fi�]ou�]�UnlXM�(��:*Yv��at�D�˂5�����C��0��6�o�h��)�b���d��Gg�`%��i[�ފi��:&�V���A��X�c �K$�N�G��8���z�#�r���Z�_x�[�F�R��\h��ca�6i_�ޓǏ�ѓǲ� w�����]����ӱ]_uru��Ԗ�7�?V�x�_/��S�4���mwv�$WJ�nV:����}�^���9=?7XY�A*$�t�P�YZaK�����w.MV���z�ѵ�0�֕h&����2��I�:��0���+�E6�i,S�(�S�ű�D�Q�u�X��d/Y�S�g�{�3�������9PrDS�<r�C�5�{��l�3�eoX֒Gӹ��n��:Gk��S��j#���4�l�m<���cjbt0���k�
a��m�B͑��q�V��	}���_`
w�4u8b#:o8"����'`p�4���7�lj1���z"Q�����ױbάOR�a��Nk�AqAK�t��-gs�6�*�NХ��ۢ��6�xt�Kg���#�L{�=�����V��׺�/U\oP�a�=}:���F�����뭿G���2|c�k:�sg��,�Y���@�̻��g]�"��HO_nT�b[��/C�,"2&)�J[Қ~��^ ���K�L�,?������4�%9nλ�^�mL`��6T!�^��,2���hsm�&M�&���B퇭X<@�I��c�#������f�쾕y�Ҳ0��e�q���d���a�vyH[���X���0"$�EJ4��J�+�=�*u�h�܁���g��J��ʀ�(�O<�+��`h7��Y5��aʻ%��iS�đ78��"�����s{�[o3]��p��@~d�G����C��q�u�ޮ��Rw��gW6����(E1>�ī�$�D��ƥ�._}�1���>�8`ة��Gw��\��J���SwW�Ffg3v����+������E�Ux�P��L��Yׅ���J�w&�3G3�'�h�=��<���)�Z�Zu���������5�jf��ڥ9	]1�R�8��;�!H;��Gq7����&֠#R��wi;�^���������GQ���Vɜz��H�x~��$��(�Ł�A]c������FEz�u��ܬ����5vr��=����+y��9�:�g;#�"�K)����#�$#� ��[�䆹��>X��foj�J竪q6��,���2�*����9J�ю9���Z��Kѭ=-�S��1�� ���~g� ��=ѹ��5�[ZV��W�dk��WLQ4ǒ�y�C4+;GAj
{0&Daqn\�Xj����ݶ�}��$-,���洎uUA���o�4Ǩ\i�@x���,�.���Ys$;{����GJ�>��c%X;;�0
�F?�W�uyu#g7�HTY��r)�X�C����rg��e)�V����{��U��J�wvyn2C���3�p�ys �]� UCw<?`���s ��ƎuD��/��KkyO[��-MI"MS<q�}HGi!����a����;���ΊȽ��t/�� S!����s��>a�_S�����5�_X~ ����!��t�5��YP$АȏWq��c���N)��"�*:��ɜ���w%�c5ȃ��)v�ܛ��<��g�t���`����x�L��m����증�gN��ӿ�)D��%n�#��ě�uv:���^��p���1Dǲ�-��J��R;A����e+�hy������#��$�|��� ����1}�� �g!tH�sg�ǎ#`zsekM�!F�_X��ĳ)�ܨ�ͬ��^Z)���
r�0]k"���#zU�ɂ*?����Ɋ[�CK��^F7V�Y�[;RW���B�M�Ж�� ����DA @I�E��Q�OQ�����H�)��A�aoS�5X����WD7��|��
��� �����q�l��L6��d�R���=�F9����ps�y��pt����c�������jdh�Z�r�P�� �kt��R4��-�8X��M�Z����	B�i����
��&��(Ma۠�����E����?��U��1�w�?�C�9�ͽ!U��_[�q�E�07y���떷7��}x��hkx���R瘬YI���F�(W}��ܫ��v��- $��<
W�$�!>w�D�$*�2t��{$����s᷍J8/��X��k\�!2DU�s�Z�؛�\�v��=�@�ù�M�#݅��@�{{�'-mdo��_]_�ۓ�rvv��k��9k����kF<�10};#H���II�²�nbg�CB�^�r~v�&+�IV@h�"��#���US�w�
�䩻d��X#�$��E��!��N2ݡ�� �c�;�[�,oNN����ՕKy���<|xO?���)�@E�.;Sie휑�:Al�"��]�m�#��3�gEyjH[[i :���ή<x�P>��W���Oyß^��/���,��A���Ү{;��#WHC�4� ƺ�u����vei�USGV���W������+t����{GPk-^3FJ�)��|g5f��H弿��g~	F�?�6��l����A�LA�>�@JY��u�,e��#���s5�A���d�~�[<F�@��H��xK�늻q8�hp�������"5��G)�q�H��?��UaԐ���$S`��Z�!��m#i��5�Fgւ����O?�'O?���9��{W�"Z���L^��I~|�VA׆]�К���b�v=|�������ɖ.�������#�Ƿ_˛�'�F��:OS�Ȣզ b۷��Y":�A�6`u�����.�L�2o�T��9H��;4��Z�Sb3oT���֮�:�z���r1)l��2��*����%:ej "����TH����%
��v�N�$&Eڥ��G`�ث��R�����d�Yu��'��z$�ϊUx�M��T��/��T�tAۥ�֚LC�Fc�d�ds"�&C���!�q�Xo8)���Y���-�k��lb`9��>�@��W^׏����Eo+�&H	��;�m����.<�:)��C�[�XĴ4��-M%���A�e-�ӹ��5v��ͣծ2K)�Y��r�P�7�I�`�0F�<��N��2a�[w���72)�|��p�����HSD��Y�Xd�:�RѬrӭ�<Z��x�<֖&cBA�����u#��C�ۧ��)/K�ѲF�[�a�]��x⑩H����>*�Ô7O���a�Ѭ7}4�5��"ׅ����mj��@���B��;̅�$��56����X��5R��]�1�F����Z���iʣy ��u���6�!1E�.Pr�a9p��=���$/H��  1�=^�A/�b�O�P�D����9�u[�6�/1���*7���٪�b�%�9�b�{���x�����3��F���c�(�L#Ńy2�TBJ�	�����6���`�
�������Ÿ�ѓ�/�X׻f x|n�t����P��f����R�:����J���x
kG�^�X�G-�j�/��i0���)
�'���GA��gK�+�>�/�U"�z@�hܹt@�N�B�����#7�/k�Qz9��~�׋�3N�������q�ߤP��O<,S"%��������aduAon?�I�fS5�s�+��ћ�L��c�s�H�
4ή�@��P߷PW�Q0v؂�ݵ�]�����=9�w(����2
ۼ��,��2�I��Xmd����s�Hf�KU�͊�k?�ke��J��<���z��*3j����q��P`K��1�0OUb��ɫӷ���/�����O����9:��ݻ�L�ژ��R���tG��Ρߗ�s�͡T�=v�����,�0�h xa� �l��^�o�h�H>~�����N��o��J���������)]o�s06�6W�Ԛ	��΍��\{$�2�`]�
;O�sO��f+���M1B�[�Ա
�J�.ȩ�zA�,N� �3�*w�Y�\���]�=��DezBr���@�����z/�Gj�bg!�Ǉr_e��,�_����� ���"� �w���Κ^����i���m��=��7bw14���T�԰�?��zgJ�x�;�Y�Ԕ�M��`�w:�[7Lz�Y�'l����E��7�E{1�م0�BDvL* 7""V�cz�G��,ekvAm�h��@w�ʝG�d�h��7�5�"7JX�]��W�'�����/߱Ex�i�0��9>�#/NNe�{���/d�P���T�Zefq����W�^�d��L�.�2��6x�	�82 洩}2����!��uF��=�h�{���p��j����N,0W�.G��xY�}^t��9���>C���~����w����{g��W�L�rq�����8��? �����V���s W�Mo6� }1�a������aP�6����b�:s�����kA�
�k��l��5��Z��,�u\s6�!�Le`��C��[����uN��s�{8��\V:<��e0}g���~��<�-��~�U�m��±�yy��kh��V<��R'��5�{��õ��g�!F�qlǦ���>�����/�[h3�yR���or�X��%�NMH�ʀ�r���>��:dGl����9���b/OѼ.YԖu�8Ƨ��k��,�*������HT�H����V��#+�8iGZĎ�T�����<���XwƮBc��w�r�6�3/�<����B,�z��J�ElU�C] S���\Y�$+�'����0jy������N�3��0�x�;���-���� m�/']�4��	ue�ʣnL"�$����	,Q���0��Iȣu�p&Li	�q��Hð���1V|)���0H��ę.���#~��]f�?ad���� ���:���in�#���i�u��v�D"��Q��s*h���"P}2�5*{�b9a(ڌ.s8���C�v��@�IL��������r5��a���8�����į @�Eb�k���㰴�h����7M�C������\"G�t��CG�q5��kx��N�����2�."��~�Ӑ+���r�)!g9������,1����[��ɨ~�
�vx�<W�w���j RC�G����/�h��O#=�N��Z��PLT������`ڵ��iP������Oxs�7<�q�����ٍ�+$v�<�LYS(��LK�?8��[3�v��r~q� 劎/4t���'H���:��=���+;x{M�bQ����_j5�)-l�s��w��!��F�u"����w1C�s|&S�^(�<?���J��y���>��M�n]MK�#�/�^ۙ>K3]�����f��4����������4~8G�ѣ{����J���?ʿ�_���]��9��~����ˮs;61�~5��LVЛ�_�9\<29�sw���2�����$������0i��[��Z����ᗖ�inQ��W�H֫�荂6�	f�:�V�f�����0M��%��6ܹ����"X�g3�������S��q�jek���GA6��u=��{��n�\vp@o����_)���`�d�g��S���l�S����>�d�A��5r�w�b�QC�6�[��i}F��1�^��@��{��*2�a��.~�hW��k;iMK%�+�8���_� ��K��_���|����Ӊ��T�~v�{z��_�Dh���gO)� �77��Z���%�
��G
̙�֗�f��c�o�"���9Stֆ�!����R.W7r��#��gv�6�֩�OL��2j�yݰ�e>kd�~�G<�aN[:o"%x�����Grxp��{zv��CM�ңm�5�;'٢>A�j�V3��~�C���PGK���ct ��e�bs�)e��c�I����ruqi7I���Xv\�&&�%pJy��wvt ����>��}nG�`�&v�%��CV]���� ��f���^��F�l��9��.Ku�dQ�H;�Y�]�z����1e�3���cJ&v�0�@���'�}pg�)�7�V��\�q�2�QX=<�����,�;hoa&b;�0��|����*W����|C�lUtJ��}��x��>D�G�񁨱�7��.����,$�Pdg���j�F����Yoc���d���o�.����t#l�W;��xp$P�����r�a$�0�7���<3.��`�'[�;w4(���Й���R����y����@��6���v�G��y���5 hL�:��~�>���J9 `!Y����wZOJt�^��vmW<�*��CX%��/�;"�c ������8�rpmc�ƾ������ ����u�m����S*a�ډqɧ��� u�%��4���e��(�b�(��4��i��S��+���m,�%Yg�(|�R.������J���Z�Ax���!:��YO��*�Vc K��AȘ+���b�S#�c2����o7?��x1�H�x�U4�H&VRE��aM+��ީ)
<�DykR��v�(i �U���%R��Z_�
�-�sh�zo��E��)�}��}rCٖ녂�h�[���q_2�6�47��	��Fd-��kU�g�;�%�1�Iְo�Hԑ��o$�GN�<4$����r~~!g���sWA���,ņ^ԝ]�^��>�����m0n��pǄ��;r��C%	��lU�Z�0�=y'/_�b$d�
ʺTY���9��z�5u��u ��X���/RW./���� 0�������A�¼�s⾨�w�꺓w�O�͛7Jl�队��oS�\�lO]����� O �ZC�r49 �a�����٬x蟵5G$dޱ��ǟ<������_x:�<{�@>zz_�����e����tK��RE��ĢT,��������R�ը9�������-x~<�7�K���4e��$k��ưq����h_nְכN=���y���Lm:٥��"Z�tU�;��bCF���:ef�ଟ�����F�P��\a�t�7K��->V����&<�5�l ��ݙ��֝����Q@������������+�sbj �8L�^k�{��-�-k]�d�9A�:!�<g��^���f���v�gg$������Z��$IyO*O=������0��͵�~w"w�Z�iv�d������/����_��Z��ᅼ;����INYo����g-un_�y'ӿ|�Ը�Wtf]_��<A�·o��޾$��"�PM�eI�yÚcÞF�g�����#2��\�9���w��u}OTg������%�#��j�����i�a�b 2^y�"�����{��ﲣ�t>%��`!j����ߓ�����ށꓥ�|5�Cr�cE�\^ܰ�8jV?l,	���K�T[z0�@�{�*�;<�#a�T�����b��Ip���\^\��7'J��,�'�,��̸U�q�������;���\[�V�2�x�f�D�����stH�Ǿ�ٝ�9w3��ԵCD���Rn����j/��\��s_�ry�sp�d�������ñ3!�j�L�Νs�w��g<�
������F��N�fM�����y��X�=ƌ����}ϥ^��~A��3��g��ݕ���&E-޶�8��I�;&�� �0Lӫ̱O%��v�|��1B� Q���;��rdK2'�Lo��X�]��2[z%k��B�w�L;�.�u-�KZ�a';Gփt#�����x S�>j<���l��=��Xuj����B����+K#陇ٽ�]�4&�pK�Q����w Z1z�b)<����=G)uq�9}e'4�2�E:Æ9R� F7�P�I�P�(ܧ.�"����R�N_D`�-�?|; �W��oR���V�4�%0 �2����!H���F�8�h\4H]��m��s�h-o��ҭ��r_x�D$`xm�5%�����,ŀs^E�Q�q�gzZP���OP�ʽ�����;mE0���,���MA�[�̾�B���{��`F|�Y���yaQ_E%kYQ�ɟ��&q�9u��9u�+-X��m��Y�Xx�x0o�]�<+WՋÃ`�Ϩ�)�
"1I�H������
��_�H�~ʂR1�Ld�̵gN���[�i�d������̾����ż�Ö��6!�7![�S��s0���[Goy��d�#3� ��HS5v�����W{�3e���@E���ݽC98����Z^�k� v�}���z��ʟ��j����3�J��|+ ���f ��*���%��Q����;F}��V< ��](��-��:�����ӣ:�;a*�R�)�{���\����Ts� \�()���7�0���u]���ճ����ƙuw�����s7Sy��<W�ut�K�ho[�������=���Hί�t��{��J�ֲ���Q:A7?tKg{�;�Hi�g������=y��<xpW�"�x������@�����~A���z���
��<���siFw=ը�V�j�D���|���Ƚ�{z��
x�|�c <�  ���[9=��7v5:8��`oJ}�&#�b���~��ߧXkf
���PԗVQh����z;��<�$Gwv��h�]��EcAZ,j�ޝ���^��Be �{Φ;
�j9y�����/�I�&̠���� �n�mwm�����,a-�W��G5��9@����Wnv��TE/�t��^^�듷���A4"�Hc{q&���|��7��w?(�z/+�Y�|(#�tޡ���Gs����╬�W2���a�����8/���Q=D����$�-Vp�AoN��s��ܻwW��ﰥ4�'����=�w� �MR }%�'
���r�<`�Ӎ�w'�����t��S)d]�tDz�Nf��O���u�(�9�nA�Y�	~wv�z�����c��rY��4��C��ְ'''�мU�s���BV�g�'6�h����sf�x�Q�u��꣏�˓'����#9�������>�q�l1-��$��J����B�tޜ�gE��]��F Z�ߜ��Ǘ:/�r��P챲���JX2�����g'�O?�D���q��y(����7+8�T�����w����R�J�^�P���ky�sqq�bd��M8��,3'�L���h_��y��^i�K9}��x%?�x��?1ҸG��ۓOU/�淟ɽ�wU�����H����e������Oo%��k:
q <y�|�^t�Tt��F8�(�fQ"�=���\���5�2���J'<.��z5����v:��ǆ��١<۱f�|dBu�@B�CFg7J�,��
��6I��N�M��8��V?g9�m�>�d�f��bB��੃LU0�a�����W���=zzJ��Q���d+�.YPf���׌T�$Nޢ[�M��h����e���z�� �B'���q�:.���v����!{��h����n�%��#cf*@|.鑖��F�[���GB;D�JL���PQ���:�k8�Bܰx:�����g0�n b ~l��k�.�{�����ɗ5���qc��~udFfᵢt����A��rmDὰ�z;���_�N�VY�v Ȗm[��+(r�K�Q�BI�1F�Bܾ���O)t�GSEa�7����+�~�c��$��7m�Xl�ۨe9�6��W�
"{jL�F!�٬gIa�W�$E���5V̟F]Ҭ)�L��˕��H��e�$�����)iY��[vF� �����U��J���4��������.(����×��z#���J��${m(�
���^���T~��'
�����k�0wo�Ōq�쬬����.�.�g�����9��z�TB<8R�6�����y{�$����ZY>�a�����gJ�Ը+y�`쐭�-@ti] Ch� ��T����M����7�	��Y'�?��4-=�-T���x��oⵂ��''
&�z
���u�
���>h�q����%Z+���k+ �)MCP�no�>�t!��C4�_���<���<>>��w�o���8N��ߗ?��g<��B��\	��O?����%S���sؙbR:vn��*�=�h R�>�����7�ȧ�}"O�=�g���T�(xр.�!��O�f��ݹ|��w�����^�����MӅ���F��/H/���l�>���F�<|"�<} ����X�\p���ں_�x�'/^�P��8���X���IgH�Zлr��W_ɾ�7of�m�n�́� )���*����f�}������|,?���S��m-
&O��<~yHy@
:�`>��y���o������]|���|g_Ƕ˨���X���s���K��Gv
3)�jƇH�;��)뀬��ˤ���M<�c_5�*����~���^����S���HnK�I"�k���^�~���T��P{J$u�t/�&�~�h�OJl���� b �k��.��#�w�ۄ�Vy]ޱ�$Ϟ=���� ��}^�c� N���N�����x�i���:�o��/޾�����J���nk8��q�@���ټ�now��dH�BT��ΕX�M=R��ݷ7��ֲ�����}%f3Ց�J��	�O޾����k������˳�JHnH��%S�Pȳ��p Μ{������o��L	�G���1��"�4��3�S{�.T#d��z_�ݱC��,I�ԅswJg��K}��K�P����_�ܯxx��k{�I�h�4��+�<}(�����GG쮺Gg���{���38 6�^�wW���NЉ�����/�ȗ�^�z+o�Θ���_`T�7D���4= ��ݯ���?ᳮ�W���/�?tmo���8��=�k}�_�ꉾ�S�կ?&)�[D��2�>�7t ���W?0�����Ҏ�`c���Ȝq���f�|�-�{�di�9����Tl/�I40�4l��#YmN�� �g��6v��jE'���Ӭ�+��qSY�Q;%ñ5�Y�N��-�,тs,�1<Z����6mc�i�j��)m�OMr�mX9[�>;�8_�p|5	�j��!y�J�����)��+>x�J�{k�Q�u���{=�Ȑ3]�?�+E(��)Q��_���kH��4y�2���k-ԧ�C�xx�88�m���N���tNUy������؁78 �Z�䭳;Π��0ÿ}Be W%Z�d����+���g�YC�ո�����X�X�BW3pvm��x�~T���A�1T#^}�-^�@f��w���C���sl17%]${��<��4�R�BלmR)�#R+�R��F��Ȃ�.��������MԺ�������\��.gq�hP������[���_]'�8|�X~������qAAE]L=JA��FU--��Yδ�^���M�Ѷ�"��KdBGG/z�<����9�&Y{�W���Ĕ�]���-6��C2�k�0) �U��+r�Vd��j�a8'D����8�<���@�P�uyy!��LyA:���B�H��ϵ��
���ѥ��ҨC7�KX�CK7j�8��^ɻ��D\�ݗ=�C�7��8CѠĚ��s��a� ����?�/�����g
�i�� p!�4�!��)�o޾WC���Yv$Y��.��;��7���{fʃ2�|C�`ެ���g����)Id�_�c�lH�����&xށ|5$Y-��$t��b�:�)P[�z/�o�)ƙE�|�����ik<�
��^���| Ȟ�T<~��x�^���AD���hj�iēa�	�(��5���H�v�>H�'��\>��?z4�H_^�(�ە��{L�`D��&_�|-���shþ�a�S��9��Y���w�k�R`� ��]��˿����ӏ���]q-�8�c��l��΅�́�;���A��.������k�����û�BI�o���6�e�\�M6�\��&��S O?���G����J~�ґf�G�s�6��n�={*��H{�߿ù@�u�U�<��ɻ3H}�1���;0�_���c�K]T�y��5�%� lD�z����I�@Y�h�v_������W��#��B:*RWAbpF������U�Q��յ�7�y�bm<�H��z�{��9�A�';��D�;R�@�q/6�@+~F����/wq���J2>e'OD�vTVJf�8�&�ҵ+�Ҟ���H��)Yp� �5A���\ޟ��a���g�_t��N�|���ɑ���'���>����r� ��x�K�ab��v�����������w���OD�.�u��
��,�8<\��|i��6Wl a��vl��̿���/T�>����K`G�T����s����ߵ�ddZO�	��#sB
���>z,��kݯ˛F��;��$����)���|���W�2j>�#�����@,ʨ�KH'ߟ)6>�tH��O�G��������w/��ﾗ��NO�*{k��A�w�#��D��~���)�<�n�t�d%���ߙq�?z�L����ٯ>�G:?p��y�zt�k����Yf:�Q�������R���E큍������ '��Ą���:;FC�Ȉ1gqc�ٔ)��1���3� ��8S��)8�ܱ���voxHqσ���/X�f;��ӏX�`�+D��_��;���V����b�M'F�,�Ϻ�#�f;�ڎ}�zw�͵$ݿ�q��fK���x8�*� ��hypl�'Qo����s�Ar*i~�k��Ҧ�\�h_ι�݃e(`���׽�$��ӹy�;	��Y��`7J;ߨ���	âֺ�Z���l2WH��6�B:ۄmQ�v*����Q�H���hl��5�܊LE����Oe����`�4Dk��e�ء�p1ƷE0JT�C���ϊ�S�b��m��9����!�Ԓ�{�q�Gl�R�бF,7������8.�M�V������d2��M�g.!`����9A�1��Q���|c�6����/v�La��5EM��6gHQ�w=��DXRL�F� �@�=�>�G��?2<GW"Pɣ2�g�8<x��E�A���0�].F�1'81���%�r�h�B�����v�6������R��P���ĳ��.Q���G����*�W�T�"¦����R�5h O;<Rz+�u����"X#��us4Ei�x{k�띣H+�&�6�e΢�9�h�Lg��ry����]ZJXۛ��������� ����L'}�A����W'�����j����A��; w�_ۚ/W���+�`�1�T����7�?�N>�����l�s��,��g�Y�׌���|�1�uzv!��ߪ\�P�0�&Woau3l�LDgʄ���+͕y�2�Je54�t�Q�\��հ�	=��Be�2��/����\���]e�F��̈>_A����Ã�T3�[D�&�Ou}��X��߰U�	�����=��9�s�������?���?����+���G:�s�4�TA֑���������7�Y�weg���w8�u9�o��A�S`��j�I�����gp�����Q�tW�����_�����TAٽ�s8O ��q��(��]�1R� �3�y� ��u-�	��|B�~��������߿7�c�6����\e������'�o~����w�˓���33	?&l�		�>ǡ�ό����O�==yxOI��؝�G���߿����7�)wJ�f����c��8H�mlA)C4�Y7��<v~.�Z+����� �t̙��x6��Zë���N�NO�8ܛ���>��x��>����S���N��l>۬z��I�$�?���F����`�X#�Y@� �b6Qb���ޑ<zpO	�#����L���h��f�ؘ9k��ِ	Rg�4�H3t�*�3�|�gUD�Wz������L';{��Γ��#{;���G��_��$3PL�5�-�$�x�x ��7A�&�TM���s
l[�F<J8���ן?��6����g?��{%?��J^�|�s~�5D��O�)�z&_(�����ӏ�3}�(�!:�^�_��Պvbo��3�����Jv���l��h�r��w��z"O��X~x�:�k%��݈�<zxG�={�H�'�<#��S�8׉Fg���Zg�iy�L�J��Zc�bH��=%������'���G�����_�L����t�n��:G��T�*�>d/ ��F��X��7J�v�[�3˱���{Ǻ?���ʘ��}�3��}f࠺���ɑ���'��)Bm\�j���\�n�³�:sN�w�g�a�C/�f�w�l#8L�gP�
��xG�:G�V`����J�n�/���./����w�?Q�3%�e�uSԔ�z���yF2�nϦ�$Cf�72zx�^��9b�����9��/<rU��ʧ)y�������j,��n�(D8�m-���E�J2�t0�#�R��82�5��_�b�V��H��ԃQw�8$�G���o������ �`4[�|�"x[�s���}�*�0��P���ut󓷙�2��ZMm�X����#h� =��r��u$�X���&YJ�_ D4��Ϊ�D�\@,����指
�����<yKo����5���Řؙ�f7��:[,^�>�3����Ľ�eg�عg� ���Qc�4���1ԾFh$D��v�P����yh� Y@����g܇��[;�xS�އT������χȖn�m\A�H��F�mjk#G��3�1� �����1���<�6_0��<¬��>��(A.���3�J�0Ǎ�ɎY0R�`Q2u��t��]n��r��ᨹ����%�$�H&;�."��7i|���]�B"-��A3�)�8�Һ�D
,���ժpM�YKDxhgom�Q��&�ѻ�ڽ:��s,���v�"�����=HT��}�Ƅؼۦ|�\��:���r�Ho)�C�皨a�{|W��]z|1�(~�S`���%���U� ���r����n���;�]^ޓ�����[�>E,�׌��v J p������	���g���UFQd+Sc7�k6�0c��%x�
�',�7G�ru������}��������FCz]��Іr�������"�	N|t�;ؑ;
������Յu��օS<�À/�\-k�Pp^Ցڛ؍��|��8�]��NAf���k3;m�5H�C��g*��'�8 Ҩ�� k��)��xﺉ���O쨆�ԏ=��8R=�H��V/�Lҽ;�����+�S�mVrW��'���T:oY�Ĉ<�HO�1� ��`W>S@���-��/��_=�;w���8Ev�p���Z����>A\rߞٍL0���<�P���h�[���O��䅥��8��?Ps���?�?������'ϟ�׽���x�ioځ���Ab2G�k|�O�꾹�?�˗_�Hߙ.�Ņ�U��<��>�G�l�ؓ��%R?�4��w�y!^�)���(0���)*�;u2qt�AD���Wr����ZrdG���J-JKh���4�ͼs����p�l�(��Z�xn�~���O�U����us77�?��n�%�{Xϟ>��1�D�@uE
t����R��x��K�WT�g���͖	C�TnP�9��b|�(��᡼y�L^jb0!�}M�ё�y !��l�I)��P 1 4�k��ڬ5�=��PmU
g��ލt����4vM��9k���������K9�u?CA�p�")~�����r?�f|�$2���vv�uZ��M���ݞז�y��������!��H�7<���w��� ?��Gy��y��X�y��S�)P�p8�O��r7�L:�{����. �b˙kt��Tc�d:ѿg<�:�mM3�u���%c�@}�E�?+��{����^��7aLaT�L�hWm�1@_�Vz��<���k�y�hed��c�L�r�!���rx� i[�����f���9;}]��bΏ����^��߫��vP��ya�T&O�%NaG!lMv�U�yV�-uХ�f���W,��l�!�[7�7D ��l[��ɒJ�����f"A��#'pВz.��E}�+�@9�7�����ٴd��	�1gN��<6��5Oحb.eE'愈�N��?�.����YX����͕[��8	�#�R:`%�s�Ȼr)�ɢl�CZң<:YT�P	Y݇8(����+��c0�Y�$� T���5Z8��g���S��`� 0nV�i8���%�PA��(�E���%<��c�r�d �8��V�Frm]T�r1����"�E&?jU㬒&��N�`��ܫ��%���)�ě���!<���n�mEdnҡ�̜�#�*��q���u�4a�@���b�NB�(�4&�It;�BB�V�n�V[W[�!7���k��Z���5�!� �	^; 9k�P�|�a���m�0�f��@ �NN��"h�q
*�1*�=&����9�T?�L�+>(�� ��l��u��D6`��Éo������$HE��b �1���8�Lx��"-�<���p���k&b����H��Q��ˤ��ǽ�b��R9�iK�*�$������ ��
]�hB�?�Ӥ��Pכ�R���%~G|�BQ��M�&˼��&oE�2)i~�{��M���KO� 7�۲��s�:��0i1�u& ֑AB���%�pnE��c#.�nwQ�"0r�"��!GAR�G���/� ,�K�E�a,��dE"�`Q�"!�n�j�L��� ܽ�}?u~��|��݉����#�@V䉟��ֽ����n�@��S.ޓCt���2���
ݜ�ݮ�������W����i"rD�!��r�3�[.�Dc��B)�^�o���U�z� �9}�#O����y_C��-8#�y�7��K�aƃo�*I�D'���fh���j��&;;ݸ�'\7	�
�c���7Zh��� e��	z���z�u�h�ѬyU4%%��.(b�B��Pc���T>��(�g2P Z}yH���F�?qd4�u��P�qy����>N�	��:W`���Dvw��p���t9gx�lTC���~Oz
lzH�4 q��v���Ɛ�,������ʓ'�
�����o����}V�Am�|�Ro�"����jLv��D-��y�/>`'u�ܠhYo��{��*x�Z�з~n����S��&��ˏ�lq,��/��z͋�� V=c|	� kRl�������di"�$�������"i�C858����
��8�r<��c�}��myEޱB8,�ƞ0Y�a�����h� �����r���HNK�G���N��`�k��Q�[ ��7(�/�gH£ʊ�q�@ʥ�Kpw��;"�Ȋ���)g'ѹz� @k_�f.��`]k1����5�:x߽�CJ��w[�"�<Ȇp�u��� ��7��tl���ܡ����˹��.�H�;�������MDs�e�!��AF�/*�iaZ �v&����g,�i;���VG�E�׏"B�֔-]��
.�]���?��~�����P������?*p:М ��i���u?�}������{���� �f�T�&O�P��Ç�|��vv~&�77\;�������~��{�q�:�:>ړi�������t��BJ{�����'[b��u�h���s�l�==�8�k�j)����*��v&ݭ��P�/�Ӈ�\_^����8;S�-�u�q��@����ּ�D�� ���AJX��B"�3h��7ry}'�يs�&2Qg�fl��f��̰kd�����6��b���9� ��{�{S瞏��>C|M���*���&����;�Ma7�D���z�
�K�n9)kI2��9�.�G�3����~�'�V�
3�։��	���y3���:�
H$�9���d��]�z����V���{�ʱŧ� V�[�%-�e�ɾ�C ��ϡ�Xw�ӀPP5DKKҸ���eO�WD�vs�0G�^��A2��>��屧N�C/�:X�`3����ht2�(gY�����A\濓��TܤX8�̧?�B��(�D�]�҄X,�6��F �D'�p�x���D��&�B��ϝ�jY�G�1���;�i� úQ�Iу��mN�KS�אzE@���t4��� �`A4b� ����'E�D�* Pi�n���EU���ڠ%�6C	�|*4���\.���͖t5a�B%]�je`��r k~/x���Y�z�7�4�2�n��D��z%�y��4�K$,�<k�wF�*�XӠq��3��h&h\u>��Z�\�uH�v��Q�,9�o�֥�����V����
�&�W�{���֫��|�����y�}�V�y��4���QVV��8�\���5�|��+��� hU����)�����'} �S��uO��b`]�&;�
>7�\�6�|�hi���bPP��wY��%���D�[A���D.�����.�x�*p������+vʠ������ _�!�V��
��ho�NWv4	��=@ER��S]5Q�C37x�U������*3t��s2f��,���DXY=��qN�5���ѡ�z�D^�:U��Z�>9`���1�P�XA��A�9Tmq1��4#x����RL�1#���IJ ���[�ΗT:�@�a�D��.zm Zsr�!�0��ڛ�)����\O9����̅ᏤI[���c��I"�K��Ϣ����r� ���3^�r9�՛c99���ܠ����ş�d$grvy'o�}fR��-'#7�� ^1��8��?7�ji�%�U]_]˻w���otO*�YLY�����gO��tM �jt	׋�@��
�q��F,��DT���;���ރ&��r}}#��}m�0�h2���KM�~��޼��&D 0H���&��cv���d1�QL �x4�S���{}Mh��vI����)���fhQ�?�$�}��;��'�u�+P�g���pC���A��:���L���+@ۖ���*���]9:ܣJ�I�s�edb(��z��Zq��7�3=��[������	�̓ �;Xx��mO������*����Dy��i���OFT� ���Ãc�/6WE5�8��Č	Y\Xgɤ���K�# X����r>����#y��^�פ��`O��Xӭ�- �|��|D��/�?�׫������zz�n5ܫzM��p��Q��<�����
��X��罼�*s�6�Q��#ɬh[��rU� P�\�d�դq4�L��K�#9W0qH���w�<������'�vmA$����4t�NO�����
Mܙ��J�De>��"o� �C]���Y�- 0C�Q뉂Vv�q����!������?��u�ϰ�ݣ���/�)�c!fwoK^(���O�^<"[��u��z��;��y<����Z>|��q� ���������r����
��z�@���|����P)���uF,uL%����� .��:1��IQ� ���3 �w�?�
��F9��RҸN*5@lE�$6
v����T �I=�̕��c�zJm��
L�qN,g���ǰч�e�s_o9Y[V����S�֒j#H��X�{'v9�<�d9q���p���XED��v/b2�T�.����c�kYTE)�����L]��5��&R��T�8�U�F�����q�ع��U�P��D���CP$��	���Z�`���:���F����,l����^e#��~EU2p�+�;�>�2X"��1Al1�'VF0%u$O��*T�7�����5����3p��|b��3���"$�\P{YNEa�4����
�&70��.�$�ݘx��0;!����U<8��8"�kJ�VJ33���j"�ј�,�|,������ª�̺B����ʥnL�����ŧ�y�/Cb�Ġ�Z��ll�yt�(���[�����\��\�'
�fz��f�)�S������Q�no���Zf�+�|P)O��L�ID�U�qAЊ5���	�	���L�EDzhIz�~d)����ps�͋�$���K��P�*��WcKh��$%o9�(6y�N5:TkZSI	�6����G��3S�,�+�krZ�m�� �s'VT0 �ׄ�����҃�JV�;�;x��*%)+��jD?̀p����uX%i�O5i3Hu����y��-+��6�[��d�A�������@�,%1'�5_���k`1�5���1׋���"�h8�
��N��sMP�M��o�0�n��+�Q��U]7'��P��{V3n8=V��l!���(��ӻgR����e��`�������;H�@�3A���%�1⡂,����]�ҼL껀���-��"�O����TF��Pe 8Ei��+*Ai����<��s��Y1I�2P�&�4u5�:�������+&���M
$�쪉F��M��ۏ���g=\x /A7�l�&Q����SA��@�ݣcP�z(=�`gO^>{.�7w2�̸ؐqi��g�N�p��@�t-�x�,m �!���.����ŽQ�zk�����C�X�0ph�@������G���P~x�L��������3��k�����߿����r��>�����U��ʙ��Bࡢ�1�]��D�&����T��o����˵>������/����NϢ6��M����=?���铺�wƃ{KA�|.�ݺ|�ɯ�~f%�vp����n��7O�/�^�����Lz���=�V5�܌�j���;�m}���{��5@����阀��ͺ&��������,�f��آ�������ءI�>�CM����O�y/Ot}u,$A�b���9�4)��D����d���B7l)㙂���U�^O��k���?�Q;�Vf�TT޼|�@�\c�ON�N�:#�M�J]�o����U��3��*�}��2*K���C� [7,Dh|�"t�j2]Try��g��*`M:�E*Q8DAC�OA6�y�Q�f�a!�M���It�`���ic
��d	���i��Q���7��{WG���^�9�3?��n��˹������Gvz���������T�pw��J��t�*|�c]K�2}�
���~jupx"G�r�� �3h�o�eW�$h��O��J!�r۠R�֬�u4�Mi9���E��=�g���<�Nd��g�q
t�I	59+��~G�J��g������\�XG�e=��w���������3��NGϤ�އ�
�z̍2�����J�~�{��BA�-��Y_���g���d
(O��u$;������ٱl��Cxb͟c	l!�O�L5� �sd�����\���ļ��%�~i��:(�ʦ��Y��=�՛�{(���
��k�ΑV�Ti�8��te"�5��$�y��� @�dy-m�T�*3��5��v%���s����`�d\A���<b�mC�l�1�AᏊ{+D �xi�Рe65F�
�AG�tB�Z��X�/d���k��I�܌�`�ր��+L��q +ƫ��=�{S(�D5&�%��� P��f(�b�2�s��zZ���/����@��?3N)	b�(�ƅiX��Yj��c�CI���gY<�nJ��,�6���K�d}#���2q���C�R=*z�&,��������%�B�����H,i���� �Xُ���45�����9��sT+޸8��5g���b�*�*�Ea��غ`�e7�.�
,��t��	�h@��\iR��Ć��tS�)�`��IF":��&�+�!�4UE�*`h�	E Ό�\Ę�#�L�U��+T2r�-60��@	��X�
�z��M��(,�OL���Č��	ȇ�B	�st�p:@j'Σ�wrg�1�M�Q�ǥLZ���&��YkA�p='�{�Iy��jgx~e�L9-a�qJ3��\��~,�Xs��A��|.l����z=u
߂�4�FhuCN�$���}AQ 3J%�����{Ea���,�x$\l]����������	�Lv�E�4b[�@��(�\K&��^�;����f�O$��IQ��G,j�R�s3/�]�>���Uɢ8�W^L9P����"����@
����_j�,H�(���L� T��x(���������^�~�guv��D�����@ǰ��8�lA)�N�Ry�ݻ�U�1F7���K�Kղ%�� cJ�[��f|H�m^�^W�+���f".����O�!m����F7�ꕞ��ր	q�bt���-J��)5eq���ߵ�%�h	�N��v�����qH�4MY�@l*����U^t� 0��M���rv;��qν8.YI}���������4���㳴����vv���0����I(�ˀ9$鵉^W� ������,5�����a�ϻ����޳[Z^��/	v|��(
�x0�#u����<��՘]��Յ&�C�529zr ��۔o_, �<�k}?�>�*�𦙣C���:��P�7�=>W��Q]{����h���X��bJ�&��\�4aCRA��ق���m&����k���=����!�Z��ޫHn�������Q���`<99�C���p�TL������������ ���4�i�) ҵ������X��ݧ"bjo�m"VcN����`����u��%�ǧ��{��
ܩ���}���+MT?����v2�M�!�<� [k4�?�}����<VG4?���s�`�Dv��4!]3I�},}_z/qq�IK6s��$�0I�[ɕw�6�����x:>��r��b^�Y�/_�٭�s=}rHe?�@ДMp2M9sE�0F��f��n���i�=9:T����`8��lE5R��q���h�8��%�L�Ny�B�t�0�����������2o���9'���'�W ����~O����x�p��M��u���j`��y`*+�5.&�<��O_>J��%5�=:�dH�O�-�p�XG7�������!
�P�KF���3�iw�K;���`�[Ø7����
ߛ}��}��&��8vY�69��L���A���71c:��AA�DzOG�1��9�򄪣E11C�h���Z,��3C��P�[!g���r�CM��|�0�����{u� ���Ls�9���)tm�~O�x����4,�=�����r?x�{���_p�g�5B�v�)�~|�	\\��D;@p�!nr=��{���ʿ�p&�wC%3��Au��@���)y������_�xG��0u�p��>.bφ����/+Y�6l/�`��Z(N8M�k�AD.M<r�S�c�k ��ܺr�ќq-vR�C�Mxe8#wQ;Qa���G���"�t�Օ��Sy�h9]й�v�<�i���0�PC��6����${��Sq��Lb�qHTd�X
R���Ng<K�Ib��R��P>{�䗮�1� �`�֊� �pmH�ᗂ� ��ϊ��m=lN���H�<��d,���N�P�N9��פ��@��\Y�U���FK� m;\l.U�O�Z�t
�2���jT�ݜ��f
]��P��Zw�Ò�2�EA���b�f����4�;�W'@>3�{ܲR����-gi�Y���t��s&�P�A7,�g��1��LqɂS���'(4��D6��%���6�1�:hX�,t H���T�`v��z�n�	=��+�u��b���c�q�u�wBm���ې�Q�L�q8�!�2a�EXgk{� ����d���� r��D�u^�3���(�<�>MM�
��LA��
�w����`3Bk&f��J�:b7�NJ�����!��U��[qI!�L%�7��П�4���٣6 AeE ��w�֐6f�0�/��sy)�&�I�:H܄!���j.MfIK����8#���y��Ƕ�H��g5=p������o��U�P��x�7*ͦz�b�,�0�T���>'I�-R,&d�V��M�v4�$U���8U���e�q���T�誕8ИU$p�6�vjk��ڀ9��@!��8�C{�c����c|~��
R��R./����>�o�����'*vA�ԉb�U��E$f�us�X��O��Z��z�����  �>�J���,�?�ipE0�ne�����)�W� ����_��s>?,F�h�t������9�B6V��La���@t�`G���m_��MƦTm�'6�� ��˯r�I�ln�2��!Ϯ*YͲgL(��%���`
Ք+21��1c6��n1�8�ej���S�~�$�J��Ӯ���H0�mR���ohҹMCW�Bܨ����4JO������ӻs���&��^>~�Bzj�hl�-V�Fe���n[��s��g�H���@`CRT|+�k-��Ge�������Ky���>���q@�U�Q�sx-����RϪŬ��P<:�����o��ړnƺw�CTT���Xśt'
�Fm�U�T=��o����%��+�d��]=��)x.�ލ�sy��g}�c
a��������j��2J_����=����l1��]�\(�*�J+v0���rtT�3�����;6�KRC�}�[4���Z���p8��|�g�l�Lp��o(v���q�^F9&��Y�dN�ԘJ�x2�����b+�
+��	�Ld{���"胀�A o�$66�@(���GXWTQ��淵�w�o^=���J�gT�.�:FH_���%�j��:���|���A:4
�)���޾�։>�)�#c;����]��Fhjpn1�~4������)�$zP�кD�	(��{"��,r�+�H�}�,]�~h����; ��)��{܏��a:X��]�B�����F�ק���^��%D�����Fd<�{�����4�O�>r�,�Lr��s��w��|:����a�=��Jj��e(�"W��#�x���x3+�}��ý�]���f(�X����½p�@|7E����k4��4�:t:���s{)20FlL!��)w?*#{��t���ͭer��v�q�ȺϠ]{>�aÈ�g:6�|f��ll�d=;���U���O���P��`�&$��T�8�N����XI����F[�x��)ܰ0�
 ��
��jb�ȥ��m��p�������%έ�7�Z���Һe���Cƹ&ɏ*!r_�Y���Y���̙��4�~r�/?��'/�Ç!h��pe4'\�r������5M8��mmi@�0	��9c�����5�g�M�� �4#G�a������ݑ�[Yq�����k>;����l���а����Xy�`>i�T7L����s��%���m�%�V��I�����Ti�ֺ.�ԫE5R��;��#0cE�Z�ilp�������A��։jPI-K��
(^�����M�u�1� f��N�b��9��jS!I;�=>���D��y�d��=���Lf��v;kX����z��ݽ���)&~�Uk2&L��@� �tcDT�G�:���C�$UT���؂�@�؆~o::�s��R�3����0+�z����Լ�h5-	
� dЙ0�?�D��K����v��e���b��A������0�NF�J[(��Aǳ�Ȏ�lmt��!9�ý�X|���I��O�d�zC��������1���?Tk��;T^l�e"�G�"����dx��"�`F	�`�IB� ����Ʊ�,�X��j�fPsQ��̡6��҈ ��<�l�R!��Fs�A������v|
���DYI�PGG��t_� (L�		/�/X�(�L�cL`ĸZ�C@�Eb��oo�����|�x.��J��c�bϑ�Ai=� ݍ��.�����s�[ݔjp[��lo�^h7m~tWRB��S�Y���u�]�s�� u���ŗsg���{a��&&
`t��Γʔ� ���(��c&Nb��{���?��>�L��D�H�	�&�n��؃�^bUHS͵!�|��능��T�@ᙀV�PN v��r&�U�8Y��&���$k��5!���z��i�:�3��9˙��} L��U@�L�n�
b+����w|T �����hN*��qN73�/k�U�A�l��s{^4�w�ܾ����x��l��!���
�J*�U��DG�������
<��3�n�q�&�ؿ�irvk:[�#�z�_��&TR�=Ik<�$x��M��?�a^hx�����_FЉ6�+
�����|�L���A���H�*P�Q�U�RZY�������z��lg�ma�iG��N�����{*�N�C ������O���Z���t
B�K����	@���3�;Bp
�)����I���h2���M2=Z�ڦ�4�c��"YM�� �$���V�̵�&��k͙#(2�����v����Y��T�m��9im |8�@�ì���a����,u��G���'(��Y�`�J�����*���O���99�������5?>tײ���n�k����,�^��^��e��f#'���<vf|�����N hx�M'���ۼ9��L�Pl��^>�������=0�@^,�I!��W�7r3�P�a�ߒ�~S�V�k�ȱ>*�5��y��9VPq�V�� +`/L�A��������������9��uɬ3���P����X���/b����x��a�ʔI@���j�樋��%�m�*t���X�]�<a;Yp��,<��
�(Ys�@�N0��U<@7���7����%�����f����	��]z�,�(}?����'@X���1��| P�`@f�˪6߷?�1�b��.6�L�̈ӋԜ7�p*g�rs�����v�p����8b���o�k���3�ׂ�(���X�4�ϱr$&'n�
~��=�� �0��S5j]�IN�fb�C�S$%��=���s���/u��ȳ�1���6%�AU�������k��gg����\\��  ��������:u �n���XeA�p����W\jJ/�����$��N_q ]@��/}��ՠ|Ik故�y����s���ȣ�j�xڝ���qsY׍C��n��{�� 3
c���qp�����|1a{�`����á�k��������%)G :��:�9����V��ʘ��j͍��V�0�$�T��(Yei��Nt�������]l>\*����z@��Y���O������J	&�b�0[h�w2x�a��ς�n�	 *p8`�҂�(��C���s^�|fE�7��V��`�N�2��� �z���7��*Mv� �E���	�����~J���4Q���חrA�\�a�`���s�(Tmk�*����s%��`A�C�
A>?�~ ;�Zo�,+e+.�[��#D�Δcv����XxNH������	NFq����@c݅�Qt~�>v���|��8��(���Ѕ�,�sF����Z���su��W�f��L�!�B�-h������dt@�����`b<��]k�*]*���������*�7�3Az`���*a�����>c����&Aw5��t�~��Ԡ)�
ЉA���z�p+.�T��A��'A�{���h(zO�v�º��U�)��@GEe�5$wc7>]s���G� �I<̑�g��ݣWP]�2Uͺ�Oa}ЅP�S�㊳��[�X2���|�A��L�w�X��u�L����u������3.�2Y� ���g��	� 
���B����^�WM��4�p��f�`̧���5ά�<W�:���LF�Cx���-Ίԓc�q�^�P�Al�ޢ�`[�%���|�}��`pw��7�g�X@�>H>�>��5ku���b�����UgQ �������"Y�G1�+k\�Ӑ���P��DS6SR��h�#lP�Ѫ�0��])��s��G2��ߣЅĲ���w��QY\�?:��)I��`gc���x�/cj�׺���}�Z�z��v�.wO'�'�P�i_�k�?�&�O�zN����8V*(�~��p�9���8W ���6g=����π�%6��n�Zc�1ju����/i���r	����0�sꗦ<�!����&;>��8Gnx���*X;P@5����̊���[]��\��z*�_/)�tp�-����A������xex}�
 !��@���]cc_�|�g殼ze����
��5�X�P}=�ܓ���ԯ��?��=��\�H��/9�ys����"+���k�b���s���wr��V&3PE���Ἢ%&�����s[
���Ŏ5��m�ts�{�`���BN����ua4��H����?{�yćO��_��/���wΨ����f�6��.���i݁��ҹ� �Ŀ��c�9�{^��Nb�+��s��>���_��:�i��*xV��Y� ��MdϺU���v� �i�����ֈ�$6�8���_Ì̓��F��U	p�7	��I�h\m��G�|D*t�xOȪ�����yg�h��W��<\�����qءU�޸�U��O7�7$=�V9��\c�|�U�i/��c+�f%����c
%��� �1�u./��7U+9,�|f6H�B�������Ej�p�)zP��T�hx��׉��0���p�j.��a���k�z��b���RM[rx��j��F���Ɛ�HY�5C���W9���](mA��|�����=:��0�v����}�u뤆!P�� 0�/�!(!y�tzf(�$���Ni�ZT{��f4����7����"�G� k4��ה��=(ʹXm�&��
\��{��A�\���2E����u:�,����X���� ��	���uFG��z�$	�b毐{'��,���\� Y�mH۶��O��%�F�ej���@�9�ܣ��������G�&��drX�; hn*��¾E6���9dA�c�}���n�iҌ�
%�hTFHp����h�͵��w�����CEs:���R�������TTD	��r��\Gf ��A�ܳ�{��n)7M��CfK,���� :�h��$^����fC��ٓ;�zT0�|A��e	�%12��>'L>@{�vxgaV�
���葁!r�JWՊI���L֤��X���U|DL�ss@̀��8 *Qm�V��(��YGkS�[N����k����<q*�'�\?���\�7?�̙lQ����y��F��i��}�L�d2�k�s��s[i4k��4���Ip  ��С��)jK�^�Thй�6	�$�_x�ļ����G�T��ݱ9J=y�8ׅ*�|3�rJx=q�.�uq��h��ঠ�����l/ ��M�a���������뫯
/�1����d�uΙ�<&��}Ib�����n�����|��b��=��9:<�ӣ=zf!N*����_̴����ťQ>�5@��o�9�}�9r��������u������hib������|V��m�(4��/�(�V0mI�F���s�5�Xd	A�r1����{v�����-MD5�,I=�b�U����|��+ʹ[ ��a���0�o�-�.�̑4�5�m��
@��q���<�3�G1�����dIh����8}pC�|�8��@VRBy��8��[�#p�6晏σ�W��tm]��^`��p|�b:z�ӧJ/
#~A.|t�+0�����/s�boC��^w�f�,eH'�WhJ�9�^�k��y�6�Q S��}ҷWT��	��;S�l����i�(҇tB�m ?���w]���ݸU�)������4柸�0����3��@O�|(� k�P�a�jEYyZT��lő�l�p��M�TVΣF��=���s)�\vmL�� w�?�s�ۜ��J�h6k�����׻�)�q�W0?����i[�=��3#�c�}J ��nEf�@0p���B�}F��f9�.�ـ���F���k-r��pTE�+�i�R��(��9ݎ���}��6sl4`�̐ójAK�?�}����P����f��C��Қ lF�jkD�����˃*������nƊ���/Թ�Q`*�㱏"�|��k\�$���4e
63ޡ�z��4rz�3��7@,�����]�	f��0���?=bS��Ҭ�AY��1��am�G�c!���$�dE.����&�[���D�f�<x���RC'*��$2Ie�,�8�t �3��s����m�0Ț-C ���I�I���lߙ���������y囎\�U1SP� �
��Z�Z��_�p$V2�Z�='�]y�����NJX+i�!��v�y��T��x ��,s.�,���_>�t��E�G�֒�����I�w[|#�j�bєe	OGևF��g�q�BY�7J��!�t1ș�{zط��Ψ�G����&�_PEL�	��y�B
�w��es��n7�G�)*a=�[&-�*i��bե�Y�bk+�x	�c���H��n�����?����n��9gf!��˅񈻝:_��6
L8Ȓ0��;l�&]K�O�����=��)��$v�#���zƙ�����z��n�q����g����
�}]��NI1q��)0���h�NB�����-�)!��M�9x�������hb3�0:�k{��у�i��M3��/��2��p�M��`�n_Q��A���]�S�Hl(�홬V������@�	J^x�0�L����zh���#oh�}k��V�?��1)+,��Z���GE7���1(f-@�P�[s��^�'�V�L�=������S���;�]��(�A%wLJ�@0Dc�r��������k���_����'���KJ6���k>���Hn4���V�5���v��>eL�p���yph@���O��̧k5�u�VN��ld�X9���r��k�A`�]9�'�v��M1�{E��`D�f�@3\($��v�8��|O^�x"_�*ؿ��B��)�u��,�M0�Y6�	!RR��KRD��P�آg�vw�LH0�e@���@kz��� f�r~�k�(墓��3fM�����t䕞��{���b`2���n ��BLdL��E H�ˍ�
�~݄Vbɡ�IR��t�9���QBװ�2�4�������S�-�i�/xA�Z�6q��ʵ�EG}��n�*�H�[�ܧh��)��I��z��g���s�|� �7'��z��)�
dIQ���88^��"�`���H�1�����;z��
�ZR��X\	r�Xc���E(�����q.�oq�&���{�^*��_l�+�Y�;�
O���&��E����@�b5��D'ne�{2���o��Pc�`-�����RO������8�_����c��5��	� x(��yފWS�U�%>+`�`t���y^k\�z@�v>[�P������( ҕ��5�ĭ�LۺV����n��p�v[��Eu>D8q�Ik�y(l5�.ϩ��������h\���cW*��|!��ڣp�+tߗ,�,(_^��罯r�����Zש�ԅ������S�{2wL�j(�Ġ�g��a]s:=�t͡�������ɬ���%·�ҏF��̗�Ǉ���1�0��|���m]�4�[���gTs�ӳ������� �H�NS������'��;�c���"��	�����
a� �t��ZG�F��d]����@�9	�'��z��m������g�i��G��>rŐ�G�2+����~�c��A=4�'F?|܏�k4�>j��
��آp�*�J/��0[��	��/t��/�������m6��=q�+�����#����2���6��9�(D��AL�xqLb�r���x����{l�#ky��S�%�����_��M�ҕ�62�.�Q���oUK�3O�M�p�qz#��k���̦�Vq���9#�^>��~|C�����v��b,Q��X�*i
����)�bV5ʲJ�6�$
�GċES9ǝ�1�L/��'�Б��U�$9���F?�M�^(��@^>(���[��-����X��[�޹'��D�ٴcvt2���&�,k�>�Qu�(�*`FO�ɏ�W�ӇMk��9��F�a̅&�S�-��ڑ ���e��h�L��\����7�MD��!eu���sp��=nf̱soM�����7�[��
��X�jhT�y&M�;5��>n����Ȕå^Q���Y^kz�A^ q��P�y��  s-�#��-���9m�YՇ��~k*�,y��P�	w�؎}�Y��em U��$�o�CϠ>��R�zh�� H��T7���wm�]�Ue�ssl�'���eC���(�i��ú�%�X��� �3+���Q���ԓ�����K���N��͝\(88�J�K�m#�Â�D�x|_����TPD������~�HU��1n̓ʙy5�N�.OO��y#���?ɏ?��gOO�\�ἃw?Ⱥ�:q�{{�J����2��Ж�z�T>~:�[�y�'VL���$��|y�y0�t���R'u����vON��ox.H�Y%3�H	_�b��n3�%𛩪�<}z���P>���)a���܏�<�`93BB�l�֪(��[�����=~�n����YG�����v�M��~P���������]��j*��P���<"���������7��`F-�E�BL�B-v�YaĊ{xt 5T���	��L8�Uz��~[S�fцQ�!N�5��ɉ�m&7ibq�cP2���aB5�-	ޓ���Ok���J�]	;?{m(�
�! }�I�t|"���r�e������ڡtT���F���:-�
j���u�8�ą� �J�R�������6���s������Ͻ�9o^q����I�o�xe��J�	��N6yQ�/�� ks�H��^��\
�?������� ."�F� m6a�b���>v�󗕌W7s���nweg�'�[[fUPZ��
�2}�V֥�(���|#X`��BE��"�=o���(�jE7����`�A���^�������p�2ԯ����3�`�l��I��f�ۇ��M=9����&��xbL� �;|�bA�*��`����Sy��EvZ0�gV�2z�Up5v�*6����w�#����W�J�+�� ���,�[�2�(bA���Zۗ�~x� oN� 0n0o���g9;���_���u�{q	q��`f�����BahM��&i��>�Fj � �L |���NNN�5��m�Q�	��[�In���c�<[�n�@�MAk�:�b�/�2 ��U�����`-0�F��p��u��aF�3u�+iދBMe-����GVKF�Y��� 1���uGQ$.\��96r�؅���
�� ���(h:�a�j��:_T��3��Q����0���|igA�u�P��,�yp�3gvѸ������y��Է�?�A�c��E� ��]���o�7h遺z�,4e��L�6�4�!A�F)L���=��AZ�kD�7򇏭�0O:Z|h��H6��&#_���Y���0�uV6?�{w$�R=RBk��۸ %gljz@w���:}�z�L����&<$�9��s�z�Ip�H��  �>*���"y$O�^'P#�)dӒ�u����'
C��{c����	!6ɗ(�:��/á�>-�9�Z���N��[���UW���%����d�Ō��Cl�f3fŊ���+�psU�^g������K\兜]<OdVN1��E�>�k��A�̰uz Wlz-n��(��ґ���C̗<PI�z(t�ޠÕy���(�+x��9�Z�mۼ�Z��\�B�o�֙��zw��ftʸ�,��ȧ��>VPi�����(��:�	�6f�M��^�~H�[���#<4p�"���� s`Hz0���k撍z�f����mp�q�Q����H�fV�R�`�Jv=<"}����sM�TX�=�D~2�������TW��z��l^���%����)� �L�p_$��G�:;r�ua�)T�ؽD�.5z%n��%I)I�ށu"~�)���X�Eԕ''��D��g��kK�����@�a�V"�g��W}R������Y����cE1�=���޶&�/�?��o���gv��4Ƕn<�(^p�"�>��'�O���5����ى����דf;#��F���l���S�R����5I����,%�:<ܗ��)�Ll+s��I�9�� Hf�iE/���-v�С�����IXTS�B�L*{�p0G������P'�h0N�Ks�������m99�����l�IB`���⌋��k���ں��h�O���o���������-~N(��H|C�7:�8�$2oIRW���8Uegc)������l�Y��}~��<�L��vܶÞ7$��8ZU۔GyV�F��Z%;������ �*�L��J0s���|����/�[�ON��ٳc�����-���)j��hA����eeF�H�ҧ����@�G#ڊ�?X� ��ZG��}M��Y��\ι>�y�z�SU� �ҷ��op���z��P���� z�	� ���N��ӧ�7�Wr~����*����sV���(��l�\�tQL)����Վt]M���07�\�g�����ٛch����q���KS=�sT��a�s��k��-hT��=����L��(H��X��םI����������뻧�f�!|�������{��x��1f��C�£~�U���4Т��8�.P��v`��W�^r��{"%��hEp��b�[	t�����������z6Ayp1��� r�^�k
�����v��W[󽚭H�����HF��o�������~Yi�b�zg��n4
+��-x�t:v�w��2�d���Ŕ8����7t�K�]��/4�|��j�G'k��� �б���HL��(��_(Hp*��n'b;b6����Xg,��l����(��UnP�1:�D���Z���KP�s�����E� ,6e�o�Ȭ�ې�¿��:! ¼�u��si��9٘��D�6�����(H�0��x"�>өj������Yn�}����|��|Vm�5��n(�G��-f	8(P������@뱠��"��o[g��+PCݻ^�; �r�j.K���Ɵ5��ܗ$$DQRΣ5�D�iP��a����8~���0D� <�[6���T�@ eͩF�6bF��%+��9S��	Г�#99�Ʒ�j���3LfS���� K��ki�jC�W�Ҹ�n�?ȸ)x ��g!�:q%\;�77?���G�s҄b{�����-�`aI��K��"��<x��J�#	�?��w b�����	7�Q�l���3W~ӱ�&#��̙����:Ws����}#h�s�\	��
,�sVm�,��|{׆I�̪o��ӕ�9����F�	w����Wp�ͬ�9�����٥||�I��m�~�B��9�; i1?~�L5E
Z����VU.co����91���RbO��J#d�{�Xw�\��<q bM��	�7 :�$+tqЀr��d
xAEgU�^��of<��� �:>:�D�H -���nD�uEA���zu�FX7ir�k � Y������{������+=Mޑ�%���P�	&�&w
-�9a���b2��&e	��-?<����36����r�	�����H�k��@If�Z�AU~��.�  �Lf�Q㡺2����ٽ��T��K�S���I�C��9a}��l��O1��*�m*�Ӊ�-��x���㺷���X~��wM��I��{ʫ��I���Wz�>Ѥ�3o� 4��B
��E ���3s�Ǉ��Hy���]���9�/@�P�q�%���[�ǜS̟���u�8E�� 0OQ�'��i�ߠiFF˱���+����=u�e���[fr��l*p~.aNI+�4.�d^&���@���-4��v��6�۳���D�D�7V�i��Gb�&�#�r���������~�N��h��-H�?������O����0�/֌�c�O�ocM��Ln�+�[@{��G�%�VY0C�]2��8j5S����&���Uh���d[w�@se���ͤ���j�k��2��ܺO�dF�⩛~�M^o��ǂf�T> �Z�I��ß��,H�C�ʳ���W�z�o:CUQc��Q^�]-~N�6�o�T�p���@�<����u5�M3Ŀ��|y*�����

P�y����1$��up�,	�@�稲į���fkRq_M���{����ѩ	7��P���2!���@�fp����x>a."��f� �\��"��\�9�0RH���s>hޒ�k̺�,6~޽�,��
�V��v�=7�m�����Ӻ�~v�
0kH�+��
�]��&�/K�Х}��	gN1cDS]�a��
���@���ci�ʠ8^�_�Gp6jnt&Ϟ*��XW	:Bq��'z�(�����(��'2�j��ǁ��}=K�q6�}x����s�4����O��	����c�ܨ�1�%llf�v����/�|+XE�8ـ/$,�MY{�H�@�^���"�Gu`���]�V��nZ�	@6��Y�]AT�,.@,ř��9��R���J.@vx�s
���,Ź��Y��	�Z�֞�G����#h��>,;HQvFE�0#�y����)��7�օ_"O����� P�]Q�W�U���ͧr�iP�i��-7\�Y���,P �@�`�` �J�5Wώ���8b)�"gU�fP��ͧ-z�!iY�:Y���uo���2�Q��B'��B;�#l%���Ԅ\G^�/y�o�L�7�h���5Y\�}Y��#I���:w�%f�@�	:8CpL�sW؋X�7��h��qÐ��b�0	J + vS�q�������FJ� <��rJ9O����ډ`�j�!���恙$�����^ɻ�_���-WT���EU�J�����6�끛;�B%+�M������\V���T��m!�T"ʟU�I�kMWN� :�.$��/��(�}$�A2���+�I���q��2o�@�A�~�_���\�'dS���c�6}��m�ɄPM������k�`�<���4�c�=�<)�[
g�L��������I��ޞ<y���A�	7�ى^�U�FP��v�T%�K$W���>�hT��͍������)���G�PY��q�8 ����k���� 3T�D�~tp�σhg;e�A��gOh�����-�.��A%�^�h3s� 3�?̽���۱\���-C&�6�ݾ���;v�$EY�_t����J3�1����SJ����S�m�l>/�����}���}� �>{��7������*@�ځ���D>~��_��|��He�gϟ�R����%˨A�A��5o�V|F�?����>)3l@����6't����4��Ɣ���)��$��	EI&z4�n�!�Rh%&e ����XM1�]+��[���;G�K����p��@��o*R��VЄzEsH�iK�R��ئ�Z��P��w��|Z�����}�G5v������p+_M5n.�CC�vvt_���? @���O���ҩ�6���HЄ�:u�{����N��A_�۶�j�Q�\1~IP34�� )��9�hՁ�ٌtIT	���']�M��g��)a����Id3EP�T@��	��U5�S���m>��ݕu/�A9���d1^�z����D'�C�]���P�+�������U�C�f~��Jн�0�d<�Z����w�|6�&���4�v�i1YA�q� :/�؈�]�Ğ1��ڶ�����ק���S9<�"؝,׼��&�6t����+����Y8�'��� i��0Ca<���ҳ��gC�=���.����
�[ s�����џo����7�V?#�I�@�QԌv�]�Ͱ�(�`���dD���zI	}|P�1?�?�`?�FT��o���^[��w ,� ެ*2(Z�΃>��ƭEAT� ����gm�B�8�����gЇ��?(�1s��m�;r'6�)n[��i��E� ��S쳙L��N��oYW� 7�*�T`qrБ?�p(�ˑ�yu�bUg̴�$�TYřk�T�*�(b�&���)mKF���pЭ�Y�5��sMj�[4q'�ɢ�ͅ~���hd��	�T�T�|�ǯ�/�h#f����<)��2��>#�!z�<��~��x�{��U�"�A���@���b�ב����@�]�<}�o�p��i�r����<I
+��͌9\�÷����@�{{[Rkf�5 ����j�ݗv��*�`]�l�����z��
����^C�`Ȼ�(CYs5��X�XiPHع�" B^�Ad�*�����6�pS�g~Ԗ�����n�x�%?������~򎴱��TAq��B���l5:d�to�Y��K4)�&���4�ל��睞�=�����-kN ��8�^���ߚ5|�4��d��~9������Ҩn9{9���e��Y�Ydj $A�O�&#�[0�P�F����%�Qi�F�jK{e4x`%�����؊j�ߙb/
�ȋ ���fj�Y��&RQpe /����n���Me���v�ޤun����a���3@��t�} z�^���\��Δ��#��Y:'W��O���k�So�.�����dfa����Ty����X��e�T]Ο��U��Z���d�~�9���q�+�@�&�;��hyBE&Z'9�g��tC��j��.Q|��,F>�4]��h�b���6v�m	�$>[��D�2�Ve��|�ڒ:к(ɎR�v*�
%��	om?�sPQa�>fU]O(	}��Y�����|�D������QanQ���1 ӝ0��P
i�RI�n� �7P$B�d���!�������noL��A���49���(�C���qտ��'7�
$tx���Ϻ10�C"~����/�h��D�9��(�a�Ƃ�~ss/WW�� 5 ��l�|D����Uȼ�l�{6����y<��k��z�JF*�fw ��R�+���5�����'��R j6�ى��+�J�8���+�Lh�g�6�00܊��C�o=$ �
/�/_�l��c������w&����`�����d��0�B��J-(��@<�،���Z��5�~���o�&H�?ؕ/���ݦ)����#�w�i��=D5����m�R��f���ϟ�������ω�L/�$��a,�.�mTPR�����I~���|��Ax0��h������W�V(�V�|~��;?� �*]�"��TC�^�ٽ!�F���x(���y<�T̈́��_M�)f�ń���עG*r0>�|@�.�5AK�w�f�s�@�b�-���4���)���MvH+�d�ɳ����H,��d�����P�Ov4f�4O�X��=xt�+��R;��xB>; ���/��S]˚������mq�|6+X�������'�ǆ����#N*�w���P�=bZ�7��S��NhBÐf���1�u`�����6��NQ�DP�	�d<��H�ҚJ`ww7�	��@�m�L:��KR@U��(̇���N��3wU(36�ܔ�y\�j������"�3�A��"�1�|��n�{J�?�A<qK��Ju�mأ������Iq����CA����\2�!^_�rmG0��%)�%�y;]Pwvh��,�.N�ȭN ���,�Fv}\}��j�ʾ��5u�qc[>|<cWe2�2슲�y��f���(.�\Er����L����}M�	0�Բ�|`��qp@cZ�'(Vx�.Pq�B�@�a��i=)),p�� ����i�؁�A��i2��E\G��ٹ�h��k�f�ks�a�(pm(�M�	P�*FA���5�`�қ�x�S=��f�b���\tD0���R�ɩ&��7��|K5�����ጝ9�C����?��|:�guzr,߿y���sv��tx=#����K�s2k���� ��������,~�^�ᳳ3�"�쿾�`�>J��Ln���v@�`n(��FP�� 	T��]�{�p�)0����J�>qm�T�H���5�ك�H;F�jIkS�#�������>��sIl���{Z�8��hn�^�J϶�͂��K�>��añ��� R��d&/^=���O��f�f�,N?�%���aq=�
5\��:'(��5`���l_����Md��Z�1Ss��˯z�"&���OKݟ�[�٘]d�����g8w\1'�}�"̦q#�n�ٽ&��9�������*g}�p�JPB�i������#��e�2��be9|�^u��8��VlsI�Ox/�}�里������q<�Ԥ�b`ܿTȣ�>飂Ϸ���G�\{�tA�8�������߬��rX6p�M����H	�G����]���󾽁�V�����Ax�8��� I�p�y���M�������XG��c���P�1�2�-(WImU{/7?�EUy��_x�Ea�8@*G�A�"uM��a�y"�v��e�Fk��+&8�	��!�����9ݜ�퀣���׫y������#�PA�����i ��A�hb��cnxH ���5�,K�A �P� ��8C�3Cp���rMdF����,N���c ���V����7��{��]}}���z���{*Μ?�a��%~���R�/b�����r6a�[��q�~��J��wwwD.��/;7����!�%�`�`xw;�����,�P�4���eA���w��LW��뻹k ���� ���̙���yq�����f2Ś��{0�� ��{iL:#�	���P?���a-�Z
�`��{�_

��u�`�@�^�xĠ�^*�YV&�-���~B��4�a�| �����!�Ʈ��������>@:���Ӭ�|�"a�� ��5��(���ْ�����W���:�5	�g�H��y�\>Y��D����A/�m#*ۥ�>?���mw�ב��!�&<�f��u���P�N�����)�Yp/2��NJ�������O�hǑ{��L���ߝ���_�	�}t���1���I�E�����}�M|�6�^K0����?����n�X� Y�5�::D�$z��iltS
D8���맜�",��AC�u)L`�y�*%�g4Z곺���8a.��H��
 ~��e@�*q�����>{v"/_>�
]q�{�`׽֨���Uu���h���w��R��i�{��j3b�Ui���3p�C2�#��x�v5;�sSOdӳ���%A&�0s���]�$Hsd�?& ��cw41��Ȼ�[�[ήZ�o��G�G�#Hɿ|�	$m0�F�2e'��",Okv{��� �vaM�(OO�#O�����o߲�����h��=�5��-�z�+��t-����@l���f9�4.�3���&_�-R�r�N�Hc됾����� �Ϛ�C:xd3t>P�]�mM��ܓ�A0JtJv	�O�%+������F����b2���3�������Xt
�c���G����l�����g�I�,h$YqT�4��N����ݓ�p"����[63=�npZ�Y�`�j���}�0R��BUfd������*�XßON��o�ۧ��L3R̤�0)��s�ԅe�XM)��Iݬ��N�I��rV�󛠵�ϰq>F�D�� |Ji����E�c�ݰ�$���ƆGY�C���ƺq-<z|���o�<���zĬ&f�11�����`���!�>M�YH�c.���<�Tamx_qO%p0`G�t�ϟO�I=���F�Wv��xFB��l�}Ft�a�=��:�7r�p���sJEn�C�'���R�I=�'.�5pu��E�R���zq��g�L(�'�+&�3��qnF�� lQ@�l���h���a��U�|k��3}>7�v�^�[�.x�b3d��X:5M�:�:�?�y�ӆ�v���J��ؿ6{��Q|��YNG��;�g�)Y#����et�r~2�bs�ƽ���v�X@Ц!��55��'�B�|�y*�1~��Q���� �����P�&w��߳�b?1/��#XP�\\��؋KA�u���Nj��А��g�g�1��XXoQ��i5ZRЀ<8�H�WB�q��c�2���}�0��>�P5��<��yL[t�u|� ��b���\��^�o%*��\E�����J�J����.�K��΁P?����0�Pd����;��t������?�@oz������M�x	~;K��,����,[���A�CV�
��Qy�MK��:�t�4ar��M0�/,��)�\��ă
8����������P�&CT��fAþ6�-]FB���"H�>��uC���\��Ԝ����51�;/����T���3-�br�1Y������Y��9�J�P�8��S��':�I��~��C_lZب��D�k=?�9(��@���,��\>h��\�����U�fĳY�K�Ko��5U���A��Κ�~�ȝ�c�����M%�Ҍ^98Hr�  O��a��eY�����U�5��?�RE�e'
�jF��>A �8^]!�_p������0��W�Z�]	ս���"޻��Ʀ3��6\r=����I�����>���A�ڋ����YL&�w
&(�(��	~>��M<f1���,�������jG�8�����~�îs��C>�$��Ku�}F k�u8a�f;�a�1N$����p��~R\e:e���d�������-U�(B��~@z��y.vR�݃c��'� ńh|@JEAq�9�9������v��n��{>@�Y=%� Y�7�<(Au�x�YUA>�W��������#�w?��m�np���I|�{��0�nZ��b�
�GA��sYd��^�5{j�����˿����/��Q����g��W7�`#�������v���74��=���ȵ
�it�H��>O�~����~��{HeAP�I��h��7A6���u��ݨ�H��=�wo����p�í�5��ݡR�����f�س��$��+��^�k���,��'�E0���x2P܇�^�X�׵~7������d`��Q�ν�R�de@<h�f%��A~ wl�$%<ce�<��쏭�m�ۆ��ݘ|Y��*]ƓԚ�zH�1�9g����˸����W���ή
/9��
��>|��~��{��||�xȄ����s�N<�2�����9�c��S5"7 Y�c�a:>9#hd��A�服�ac̓���>9��������w����)|#��@r��}��b�o|]t�K�v3��)Z��<��tJ��c5\��Sm�;$ڠ��)��,�Y����hW��.)&�����ͦml�L);���E��ɮ�]ю �A���9����9">cOMc\:���#Q.�nÇ1V��:":Q����IP܀��xm��=xHn�8ҷq�y���2�W��g���l0�U6P>)f2���B^��o <P��,A�JI%�3�[/h�{	j�Ѝ��k����fd�&U���\�Z����:�`w\�\�Ȱ������C��;�v��pYjV�H3��5��=_�"��a����m�<O͜���X�)xmg�(0\QmtH�\|�W/�P\��'K2T0G޿��=���a|�螽z��^�z��:~���=�x���T]�La]��6�����������_ �Ψ��*AL�܁��Lʔ���8@ـ�_CD����/�����*+K̃֒X�P:��_+�+����)�1�Ub�I��(~�{\�����;X�Z�||�^��V��dĄ���K��gpd�B��]�y�Z }�q?��VΔ7I|E��X��L�׺pR�q$@�=/U&\ޛ���fYY�H��Dw��_�D��űE?G��r�Afg���+�?$!���d\8�4 Kp��������V� ip�K;.2�7L��$4)6%���:�X(��xY�՚�2�
�,&��Wq�]q��3�9U�Pa@�M�U8�t�⍃���;U/��u�ZbޢM�==X����!�� �jV�!䱈����:^╒��TݥT1 Ii��|Br��%����bU�sU�Nk�ز��h�����.���`�{>w���'����Սr#$���0__�1���WsTA����&�"���<Pĉ���9�peP
 Mڥ������b�x:=�I�?6k��� �}��$B�
p�N��\�������ZL�����Ν�6��6��b(q��XO����>X���ݽ�M%[u�������� �g#Xz|>�Q�g�)RI�@�5�������l��E^2�H�`�:�%�����$�������#�pp���ò�>Qhf�߯m`�X�@ᬎ_�3���v7����x�A�b�>`W�D�\s�"��1�`���d-���[U�r��%�?�����߻��a�RFC�C<AWA*�KZ���M�丷�=V����Q����5G���� �8�ءPsY�u�ơ��ᣮ�?����!̸�<�Ҧ�:����Ͽ���Y\�O����Q����87��Bt�߂Zk�'�UZ��r?]���/ya�����iz>`uq��M>~:���۾�͙�t�2Z�o�>&`+>ۧ�?qƏŕ���V��ȯ�~m�E�9�bZ�Rj\�X�X�d� ���Z+u#f�,���}m���?�O?�@?)h�0���с��ۧ��çxo�.1��W������~0~p�^�P")b���kz�K�siL����D�pS�ʹC����&�<Y��!h�H�!�����[&.(�d4H�7]�93���uM�֜4v}q��v���>��A!묞��qc��1�ݸwvwY �Y���I���ߵ�[|�D��o��c]�>x��
�0|�A�?_ ,P�>�P�7�9��}ru���wR7��gTڠ�
�o$�Xp�`�?��`�l�ݘX�\]���-)��Hll�sbm}�@���]����x͇�L�z��h@;�:�Ypp_,�U:��}�ֿ!-#�V�5�e9�o��U��J�@k����;��>����u�Ӈq_܋�%���uY�d��z�h��f���2�n�0�u/��u��<��;���xaI%����i�[�����5�X_E����ݸ����Unqn4T 4x��om�w�����xW��ﳛ�xn��.,4b̸����Yu(��`��/ ��<!��e�S7Y*���f��
~���X7�!��p��P�CNFq�������<�+��~�;�5j�����.�Z���d��s���q�O�i��Ï���Ƅs�dSD ��+�8�\��#��?xp�<�bW��S���
Vr����1���ڧ���G���={�|
��R}��1�2 ���Mtm=�q�~�fx�Yh+�6ޫ��Ճ�%���k7K���]D����>���OX�E~
=���T3Y�Ӈ;��O�9��ai���*�ʰ��3N�)��Z�,ԍ¨�,��4: �Җ�<��sR���p6�\E��#A��b]���������|��BȒ� �Ӕ�=c.�֫湐�%�~� ׌�?��k$�t�,�tMo,��#�k��u�͊ ��>���n�wI,�`)OR�"�֕���-�y������:��s0aZ�SRy�M�p��py����^��X���%���T�L��8��t;��C�7yz8��W�		7(<H��R�M�8��ߜ������*TIz�|@���]Ġwf���X��\O��@�� �z��5)�����qAې���F7�A�V�@�Ԫ�ϙH:�s�p�� @iYT�/ д&.,@��o�!�?Pz��cq�B�gհ�+����$��җ(pc�j�
W�m�z�0c���k��~8�p�11�F^8��q���\�64��= qʾ�k_� |A�_*���/	ԢRu������Ft�:����?lA�pae�n�x �6�k�D�K��)���,���P���$Ű6s^1$�q�5q=��+G�WQ����H!�:��Đ�ZM|����5��C?o����/ȕ_�i�2��ᮮ'�r�ZZ�P�LDh:QL�NC�x�M�g�e#ѓX���_|"���<p����qRQ #��C�x&Rr�D��R���7��$o�e}U��j(b��
Y5t�|�	Ҥ�'TP.l�xK1Mn��WC�����2H�����&�0��}-�t�a$�rP�WPfH͛.d���	(����OCң�c
Ѐ6��A�y/u�ZK^>I��2�cr	5�uU��7���/��?�����o������5վ��pM��c"���G���Ec� �[�Ae��#hI�����ڱ?|�=���kk�3���MX5�dcV�h@W��,�/�ڿ�۟���WvrrƊ!|����R.�ğ~��_��ĥ�KőFː'�������3&A#���g'?_�ˆ���d�H�v��δLϰ[v-Qe���OL> 4�c���`��^��ADb}��?,� V��_��?}<f7�(��La�JP���O��CR��Ɵ݁�\�T��o�2��w���?���O$ʠ�c-=��}�ƣ��aot�8�g�C�sl����}���9�/�w_���%����J3	�s��=v��uˊkHk�U������2"�D���W��'�Ӑ�F��X�����N �?���䣓��	�2׉r���c?|�=E��~���^��<��M��x]�\�������f�3����
vl�� ��l��ՉJ�������4�f�dm�Hs%Ng^a�$f�)��7�W/�R��s�y,��6��Ɏ&͸��Pˤ�&�<����G�GR��P*�R^;�יSg1��-�Y�|�y���	�i7�y��I��cAm7��{�{��J�\Ÿ8��8���AL�{��/�����A��C�w� hA���b��ͭ��8�a%q{�ၽ~��
��"��1�D�����y����*Ʒ���X�d�i��ی�x/ juڴ�������O�����~�`�)՞ѱ* W������ښE�*�-�4������\m�~R9�G1�H�k3�/���g���{�����u�������}8d��q��Y�´���-��E��rgo#^�7���*~t}�c��c�1㸆QQ q���޻��={e>�\G����'��zj���zE�������8����؜r�
��%x7KYr��װvO?�I��)�z�gH9�  1�W��2��!G/�Q������q �R���5��k���CK�d;�o�%���L�J��{�S#}~�v
`F��=����ba��B�1�f�+%���O�CK�͙,���a�Y�:+;�AֵKYw�欆�J�t5cV��|�
7+tN��)҇����t�b�1�'�ai���zd�SKC�T�pwiV~s�[9��۔�!�E�F�'\�Жr�ν]:wЇD�y��e�aG
��W��r|8�*�"�S�f�����#xM��ll)IF�@R����N� ���H��CV�k(���"k ����/��P"�^����F�P�e����ƍɃ��:a�@Hʢ˸Hұ."��O��d���0�}R���3t/@hӎH����$r�cT�u͝g޺Z%�T�5/5r�97����`vIz-�4�=�(�� ��y]�:�	�� o?M��š��z0����f'}ȫ�P�x�|b$+;w.r���H�I������c�~���s߸�Q�Ƌ��*�PhR�ڌ�95���K}&xBnH�d!������fo�<m$jgbе3�K���q��y�j����:S�`C~�M�Ҋ����S`�����qSSz?��?	L��/u6�gsP��uO^e�]d�N_�3߾H?5� �S �U*�T<���3�+��z{� ��{3��[̜�$�*�pH?�]p�#9�����7�`}�u�gT<[�l�e�:l�o7'��������3M�q��F�5m�������1�����xh����N��vo'&�%0�^��hd�6ك��T���|�2%���'�s���J�߸1v����&�����y�g5��lз���?�#b����_Q$`'���\�[��r(�0���#�6����g���������b���]�z��g��ύ�f K����}�c�d�[�e����_�ί����궋��T{�г�P{)WS��ͮgvt|m���#Ȝ��ƙ/�m~���3�94��ܝ�;��|�s�i+Z�d��y���ћ֭���fs�l��Acώ�o���_��Z���0�'8�_,��K�		��_���@T���,ݧ�k��<S����������fD��Ø��̵Q��=��L ��Ҫ A��=������@�B%�����2&�����������6�۬$E�����U�����<�B
+g&�1����g��^�^f5&���P	��=����c�ƽ�bŝ��x��>��f�	�,�\/ ��ba�a��*���1j�Es��鞠��Όs��wA���+>�Vv��N"h����ގ�m�D㽡�6�"���#�1��}?�k�  @�v����K�x�n͍- oR[#��E����"^�x$yy�<!�_^�۫�o��G�QSg%��Zŭ̔ZV(B9�C̩�݅0�ݻ� ��#�:�0K�u� �[t�~�����=�\�����i���ɥ.���?fQt�y����YQ�==��f������=��Aį�+m⺌����u}f�x���܆��-���+�i�CX��K�G� ���=��v��(�����1ć�
��^��?��̞=�����?���Y�)����S�W���UDY#���F������?��a\C7���D��Tn)*$a�:4}>��a���:Hd�/J��S��[�2[o\P�k��F��t�Z��H���@�Ҹ[~B>9�\/��5���l��	޺�TS/������1�C��[}�g�yt����|\�Z���t-){\v����(�|��%�p����:'{&��2��ݭ��J(R�G�^�g�~pP3�9�����rz��g,����s�e�$��+�r�^�)��� 2�I�c)0S�;��bY���Eix �x�el��^�Z|����E�����EbMz�P�f��4!�äq�t�����]1�g��X������+�XJ(��H]�+��r�{�+�rKz �T��i:up���y���H� �$<��2����ɬW��$`��;M_� `s����0�ɣ�u�7�f2M<K����y)����0f�W��KVn,x��Aѿ.��I��ݍId�+𽼕���e2N�?�2�t�8t�k.c�HU��_��ߧ�PI�Kx4м2�3��R�%8�,�0�WIh���#<0$ť��AN
���'<�6A�k�dѸ:WE	��<� l���ܦՍ�l�w��܃���p��*n��䮭�k� �f�
�������V�`N��}m!󘐫�lj�\�p��\{}6�?zH�k(qJ	T�D.>���;��8_h&*$x`�j�d��G~�Uּ��@5Qm���+{��4��#�|��m{qA�=�1��Y�������ۯ��������|�B,8� ��ф@@��~+�G���11x�`��:�{�§�"{d�Bg���vS+z z��Q���T�x���`�_ǃ���]5�9n������?�?��O1>�K-y�e����GB�ͽѦm��jA(:}>9��	͡��\*�F��@c�8jH���
��������l���-�����q� ʀ黭mE����7,?����a��?�rǸ��&׷����g�xpfwbr;ޘ�3��	�B
���,��=�Ǻlۥ����
�x^u�R�f�b�	?��xߧ�۳w��������׸�^Z�A��k�ls�{�-aĒi��S�1i/ƴ��{���	'fQ���z>=�����yL�n��yH%�'���$�����KL��C,��r��p3&��	�a}B��L��4 �!��+`�a+4��BL�z=�R�;���������г	�+A/�,YYG�+�<����:y���>xo[�qo�Y~Կ�|���B�8�@��?���fӘ�`�����>|:��o�88 }J�9����Ѐ�|y~bWg�����#�m�R8hX\�-��zi�I%]��OW�nA�c}��Ɉ���h����#  ��,���FN��o������q�N�@L*m� ����uM�!(���B�����>	ZN�8����)���Fcs[2$(��5_$�R�v�bI�t�R��������Ϝ�=�?����Tk�M]�AHt!����v��������м^�"XA>��3x�7ы�еn3>��Mg�/���O�K��Ϟ��l�U��-��q��g������\���L�Ǹ~�?ͽ{v3�.AB��V2���l*8/��?�T��<���u�d�H�V�<�$$��T��4�ؿT���<_%@èQ&�h�>m��>H*�j�B`����и3��՞;�x���yD����\g��wr�����f�{@���|�\9u�
�/����,�G�P�-�9uc�E>IeF[��Y�S�l�N��4@�I�y	���	��֕CHWD���/͔7SlV��]��8L�t0~��O2��}��W��c�~���S�!�RF]�O�P����>��u��JUsM�*�l�I�+���:�ζ��J�<J����I�;�4�K�Gϭ��O��NT=�����E �-��ҥ��V������|P�|�7`�	%���g<������4���'���Q-s�͙D�0� T1S;Z�5��J ����e5�h]��1�b)�WY���o���Ql��҉�ڸ�V^d>Lٲ����۴�٩i���풯\��Wb ���C��)�=��yA"h���^�h�:��~S���Ќ����/���zоJ�:˗vM�!UY�/�%yV���_s6�3���%���5�$�����^ysݹ���*�0�{L`����*��&�_����h���S3�(Ȃ�IS2�B�yq��g� �:� @ϛF�ܡY�'��_O9{���zA�����2�hf����#%���P�܈�Θ��Z{���&��v��o��O�>^�6Ι������S���wd���F��Y+9l�!e|ȨX�K��Q�����2�"[���jՐ�W���	!lGj7� X�A�	P���l�_���#����U�A9�}e�&���ʉ�Q��bʢN*��{�bD�p��4ǝ;ۜ?}.�.ؙwe�i�JF��q�Ac�b
{���칅ae'����=�ކ����3����fAe���?�8���5�&HY� ~ `����������mX�w&�����J�T!em!7�ZɅ��� ����\��b�b����#zՅnA�6�E�c2ws5�p$���S{����A��R,�~������(_K%���KJ�:�x�q�b�~?>����{&�x� 7�{��+;:�ho?ܳ���叾z@�#(i�̑i����x\p���Е+%���O$��� KTjՁ&�<�Rq����iD��b���i��os/�dYZ^�gg��A����!��� &ֿŽ9FR��X?aB-��^�K/XɃtcWu�w�.8����8_����Y$|0g��R݋O̧�v}������U��i��Ex�mD���Kx�܏�4߳d�7��(����Y����RꊝP��TuK���������Z̨^rrA�;�����n����^�'衐�6s�cs��ei�;\g��q�ͤ�?	�2������b��}���b��딳\���	��%�񖥏�rl��'�mv'��<�����)~��k��I`��{������b�c�jc�G���S����ٝ�mmj�q<*�T�@sfxVeR�Ej�84Ōx����/^}��/���wvx|I���:vKq-�`E�{ppD*���eܯ��`0�k��������8-��a��Vϲ%@��]¼������+̷Uԕe.�I>����������Z��_4k�Ar@���ݐ�⠳/K����	�gP#��[��m;}qJq"Y�t�k���1��wϼ1��;�<�邼a��Ŗ+xPY����	��P.�K��Rg$+�u$�����������낿�PI�>U�)��,�~�
N eٕX�U���{��q�A��#���.'Nh�Y�ȁ��c���l̅�bG��D6Tw��U���G��*�vP�-��]JY�O��X����|�� Nj{Y׭$�ލ���MJn����Z�e��j�2�d��;j�>��.���yݔq��4�3G @p�JҰhL�%�6�W4�ݔ�m�ݜ�^NGmP%���o��\?6(�0��Ҡ�ko�W�4�L7��b	y�%���L�J)\f�<6��nZ@� �9&p�����>qБ\�F�yE���'��eG�i8����Q�Xڌ�K��m�5�� 珥 ƽ�b�$An����
�K��o:�|�3X�vޑ��B��5o%c.��PP�Z�&��/C�h/L>��L�]���r�.F���;mH� ��A��[�C�زN��h�s$K�UI����?���쒒��ڣ���d��,$�G@�d^�-�n�QE�vJ.:\��� ��W(���������m���_ۓ���!��u��kf����$����̾��o��yC)��df;&�����#z� Y�:b�$�io(@��77ش	�ڱ���
4-:�Ò�5�}�ĥjE-ż:hb������>��o>QE����Ŷ�h�r��y6t��A��<(�́:@����Lt�*;����.���*T�CG&�1i��n�Ca�L,��2I��a\�.����ή���������'��;���#��Q����S;���b"���0��i��qa1J�=��p��i���F���J�ސG��(��B�7S�Q�ޑq�̮��@�N�{ɵ������qݼ���J��xN�1����S{�8�ӝm���5lo�u7V'�r�|*�'ye���C��" ���!W�/P�0[xy5ejd��C��������&&y�T8��om￾F?�͘���ΈE���Z �	(��`�p��Y*���(�(nI�B4�l	�`uN�5WE0
�=���I�?�y�㉜B�W��b��d\m�X�"��xϽ:���b��`t,,���3��p�Y̐3~b6���������Wo�k���o?��ѩ<�0�J���ϵ�A����P
A�E�ƫ�����6��# ڎ�!����!�0%t ��y<_�́�?L������b�{HH�����ٍ�(����"��=��au%��ܡ�6I�0?�Z��r�y�tI��At��G`Ϲ;;{̭�={��s��ՙ�t� ���>��|']��?��?;�d�s�����ʉ,Jb\��ǫ$�"�{�~=��/c\{�����{�=�QP����6�����.�Ұ��A'������;���y��������7�<�G����9����[��0��*���U��
����o	�@��|�(���Lj�U�Y���?���sy~��sJ��@J�c 99����+!�͂�ԭi��V1#��)?M,�����R��:�0e��Z��<�[�zg�Л#���=Գfzj�
u�[�0aR:/�&O�́Sk�뱑�4Z����h��Bs���O��B�*�s[6��P.OI
 @�+�n���T�j�פ�$������ÂsTv�������߶JZɁu��1�èi%�I51nH�`uV��������A������t�*��  ��IDATi�MtZKU�$ހ��.�q��V�*�܆�!�	 �,n%s�4����ٓ����������vq3��s�x #�v5��f˳�J!�g��m-�b�N]
�c��}���H��S'P�Hv*�����+��jC���Ց����^���y�XA��@x�p������h:�	H��l���3)���e�ܜ���"f��#殖�c�o�$�ϵ����A!�9��2W�jV��wh��q�11��7�(�94�uH�u�P�����&:j������Pq@���ITT1㔧g��u�L�6>|�	�r��2̣�D��
�B��h՛T�$9_��g*b��_�d�����|�{9�2g|��RW�!��e�ZJ�S�Ȩf	#���sAɰuj�����Z��b��J1Qj�0��0��;���,����ЉZ��/Ak��xPm%���J?���zz`_L���ۄNݟN��=ZƁ��d<�=�������5�ݘ���zf���7vr���̦�Y�? ���v�ark�T��{F���>����ϛ�t�3Ҏ��������͜b�{�نY|V��#��Ԛ�TgVJ��߸� �����3}�bۃ�����[{��q|��:������$9��mms,���L�q�!Ї��ٳg�=�O�H�:�?C	V�̮����o�����O�>���"2���q����YLLo-K��
������o����wL��Ppp>��&�PP������(G�@�;&BSP<-�A�����N���Ǐ19��~����n�Ҏ0_�ۋ�� r�3�s�Z�yb`�)�S\�7 F�s�I������v��#�ݳ����$zfJ0�614�~8�^;H���6u�Z��׿�b��d �e%���Xɿ���˳}ۏ�������ݵ?�����)� *A�p1��n9�9�f���(>��{q�oa�͂o�{L��Cݒ"B0������goƅ��x�������}��+����?����P(B��rܰA�`���@����]�6�]�@Ơ�(kkѩ9�	��ɍ��d&xu�ݬ���i�j��)��)'�/�x1���h�y�\M���p��w�a�R�ܰ ��b-^td!.���NSyΰ���l6� N�cr���ƯOP��$��u�gRP���b�6�S1u�s��v6�<�d�6�Mƾ�����{���~[tɘ���<�o/"�x�VPN��?�ê>'��P2;o��4;��ev]�IiG��fNUexўw������P�@k�&p�AK�]��w�X����
���^zJkγ��0��1�8�Ƙ1��������p?�ɺ�l{k�6��Ha��p|�{��i7l<)�ON�"�<��ޝ���G�.�������u��C�	^c ey�e������9(������(���x�g����.��X�6�w��츎�~b���)j����4�9���K����^ޕy|�5�M�7���*�5��{�|8���_yC������f�ˣ���#"�Qsު	���4/(�C5o����AeRZ�̘Ӥ|���a�V�5ϳF�x�\�l6
=�
�`�$�Z�4�ǁ���}8U+�C�����оo='�@�;����z��ڕ_�l��9���/�y�3�D��WF����Y��8l�h�hĐsԩ�Ǯ�\�/B�'%��Dk]�&�@�m��(�Cr��&���uА�s�ִ:�l����x�e2�[U;T���K�֬��~�#u(�.�s�%�mjK�ƸS��/����Vr�lT��4�o�6�j|��$���~�_O�~H�v`��A�L��[G�� ]�d�&�O��)qB����^v_�R�S?; "_��Q�O��λSX���<(ܝVA�����è�R@���+.���-���ϛ%����98m�@����`N�bѷ���$!��`�u`�k��N����������i<qW�s�+�}5A$S��+9�5��b��W��g�?�[��,��\ M�?��=l=h-�P��F�L��`i�}�s���:��D!��M�[^xU���f��2T�W�Сh��)�J򂃔�N`R*�����vW��D�ܛ,���J��zj^��T]RE�t�v�Q6�l#HC� :�u<�yc}2�wK�g�F�n鉓�Y��p+]-���<�a�@�R��4+X�c��b@�1# ��h.�����D_%��_���%Q������ǯ�a��9��IaOW���?�Y�T�a&�u�
�۔X����.��.d���G�<&S���`��#�dj>��Ól}{-&�1��ߨ�!9�������z��^�|c� ���.fP� I08P�p�}�I�������G����r�7���=( F�W������u��ȳ'D��U���y�*,�S��I���F�"�|vv�p���}ppL��[ʒ�^�2���q�&�"-a����Dv���(���7!egg{���[���yU� Sqq�����م�7������E fY�܂{D�LTn�"�Č��g��L�=ܻ��D\����.�g=��	�,��|Z� ����=���ĄLk�h����x�Itj%��:�xX����G��:�����><|,�>����D�y#�)Ae\�q:���:@4��T������u��R5�˹�t�֗�MV(�=��_��G����~V;"�a�c���?� @a$�f]y��|~h$�o0H"�������;��?9��w��'�'�hj�[��3V�}�B/|������׿aG6p&����ON���8���5�F�� ؟�D�����{K>B2�-�lNoU�n]��jv�!���������S����rp�,�xI��K�p̀E���҇���7��A<�l:S��񈿏�pxp�]�}[������m�.��|��/�=8b�3Uw�l���縲{��.bL��<����m�sn��߰`�2"��0'����"��RF�U~q�g��A������v{����v��A��/��y��ǂ�,J����ݮg�Z��8k�d��h�=�pV'_C(r������n���)��� ���$�%�M���\�#[��bC�ob�g���S����U�a/8����x
�`���U�}���c.�+�xn�ͺ�Uß�kׅ������˔���>ϟ��roj<_�RH8h(�T�0xx�u�b�����Rn ��%��\h����u�����y+��o�ߋ/"I�����(ѩV���)�칙��i>F	���7�b_��3�t����N=ol�'Hs�a��#AD�Vq:ӂ���yVr��~蕅�[]y�^��Ww��#xK��C~�@�m*�ɋ� ����}��o��x(=��b%e��Pm���0���t�	!)�B��NzX��ʝ��(V(��A>X L�z��)cFE�AY�9��T�Ҭ��8ϛ:��˖<`��p0ס&��U�\r߻X�א�Ƶ��|�%���Kp:�`��,�|$w�`0& �5@?&lL$j�����ܙ|� �|���M�ZA5����B�vt�o�7�7����|a�<{��"g��Z��cR]-\$F�iK �[���잌��2�0_�����K<ܰ� ���1�=(�
��C��uڗf!��Oz#�Z�{H��m0�TT��]0&�3�����Yu(��巹9��)Y'z�%��U��B�����$H,��m�+c��TG�/B�.�e8jRG*u����p�U�֊����V�e�H,#W,�A�D+(�~�0���3_訠������:+�=����TC�Q�.P
��ö"pufƘ�p@��`�{U����*��/q���{@L& �J{���9������rk�"���F�0t��fbֶ�m;&�P�C�1"��cP�Y�nf�
�J�ut&�7Ό�{���/�2�~�&&Y���`\:�,`~"{`��*�I
� ,aݰ����:�,�Ob�t�ϴ�L��ԤzT��M�J?�I��W7{��0��+*�!����)b� ̲lФ{��TP���I�:����Zy�M��0��crжP@�<˂�=�{�������]f��*���1����5�[Hո� W5EY	P�)&����wg��UP7�1�I����͜�����Ɲm��.\��g�suwhl�)c�$>	����:&�gT<CU��ra/_p�����[�nF�(��\�N�� ҚS�L�$fIb�$�4��aW�{����Z�XJ�j%�Iqa��������`��M$�d�-"0����Ut�P�_PI\��ʁfG�tg�W�
^�Dvsˢ�Ts�3��i.�FG��PE�q�[*6>�����4# ����v|<����&�<S�C|(���I(�h"zkaIX��s�t���
L��}�q+��U`Z�y�э�J	hHO��c0[pT3�KӸ��yac|!�N�� ��6�[?9��o]Ӣ�����`D��x�=ƫ��3����ZcA��1�m��f�7d�\ö��l3�?��!��yY����,�sGn�r�;3Ϧ�� �2\]�F�uaǇg���kۊ��d(�rЭO��A|׊[�!�N��S���R�iP/��0�1�dY��!��&>�ۛ�< ǐΏg p�q�T�(D��x0����Ĭ+���I�c�[<]HN��MCn1��T�]���r`m]d��+��ȭ���m�U̅�̋�!V�D$�4��Y%-�s���;N��sL�l�瑓�H�L����OW�	dI�^�d�4��l�%~���)K�\�t�e�I��;G��-f+/޻��j�����*vTj��H1���$��J\��ѯ5m�AR�K_i&&i+�Y�~�)��@76x��.O�9m�yuLIR^�4�=
_-�)T�Ơ&��Q�|x�=��g[5�`� ��>�1��Ds�hVu��*�����A�6e�^���a�+��83�� )�½��1ZJ�خ�uA��Zp{8���z���]M_��Bb��<��0`1�ښ%�mK�$�t$ȾA@��]8h+DcC�j������H�N�90k�n�_���'�5���͍��W3���J&� ��{���c��C��~�.v�NV�Jd��J7�{G`}�ϲ1Ywo��?����[P&5K���X 3q]���oܳ ϫDiD�ǁ=�@�h$je3W7�l���N��ݴ���'1x�rވM�u<��l��#A��G�?����#����X�JE ��@���hKv�+H��bߐB\4�qd��Pb�N�IT����s�5g�D���-�*%+�/��ˠ�e��!�*ڭ�aв�eE��RCF��*��l�º�����z�;�k���ٹ�a��%ʡi�/�P
�eHv;E�f�h�`*P�ň�5�(n_'�/�s��6�/���L�A�t��)�G�v�������&�'��"�mL���0O�w6,�O�O}��!L�T�C��h�9����g9�P6~KCΝK�j116bKj��!�OD2P�@�������KŊ����;:f��wV�/�v����5��`Q3�-}\j&.��.s�L�D5=$/=��p��"Ƃs���[}Ř�bM��a�10�t^�J�Q�\Q$#��S�Ms�T\ţǇ�	%�3��>4'1��`QP4Śk��Y+��sHؤ�r�����D��!���d���$���s/�02��S�J$��T���|�Nܘ6���ɼ0!	�@�r���t�7hO]����KyI�Ǹ�����w	�850����--��Z/%�:0�-��Z/�]ԞX.:&��z��r��� ���5���iZ��+��gB��r�];셐��DO�B�����%�h����Q����B?�+Ү����;ϙ1�@�U>�O;�Ҧ�:���|�B5�Q��к��.r/f�ݑ7S�{�z��/�1�
��"P�0�:�.s������16�_G�zL 4���ފk�\� b��nn+���3@��#6p4d}��7�qEne�CK�P����&Q�����S�H@�2~�Tk�ڿ�����)�7cnpgs+����D1	J��A��{By���@�a/W�-8��=d�����y.�#P�8�;n�<Eau�爳�L��X���K0F��n�� �cTlU�}8��M>Ko}##�d��]�M�ֻERٲ���T\���=8���{I$-a��^����%Y�O1�����^T�<[��w%�Ϣ��>�%���7d���4�=!��U�7��xHR��S�CZ_�"��?�dA�H��
V�<��.����hW0!�%%ok�����C�k�Wn^���%�[u��k����+�����d����\T%�噼�����j��0����Ab�Z5��GL����"�ҿg<4��C���V?���Õ�m1-\��cYz��jd��� D;�����Yd��9��0p#U��*�U�5I��y���X��=��O��5S�@�t����N&�Cv�d�I1��l�&�\��K��Il�>����g�A���%�I����N���_%��@��<x��9Ej�oP{��k�wR�]3c���'몚��5SQ�2QغL���ke�߄�#7��4�l3���jV�8���S��q�Q����C_X��C"�'��QX�A���,����K�ܼe�_�O0�^��`c{�pP߲Y%��\�SY	�[�%ڟ��i�w���8?ve��+��.u��b�ՒØ���o`��T���`5I^<0
z��@Eb�Å�(9an����V {b�w���}'�o�ב:��i�Vi˃�(k!Y�4Β�[�6F�c�? ���u�^�4� ��9�4[J7S����Nv@�N��HY�I�I�\\k��1yU%:F���A`����YR�h���L�F�k}~|O"E�����# 9�lRPu���̩:���:��k̆|���+���:�y����-:΍�47F' k�3�7̓�2`�x�E�d0�kUװuN�e��@�h�5��[���������M�����R�p߶N��A��~qy�*�� fT���1�Y-�-�(pس�[$3��VEV�ѥ��,Bv����.rYx�3�@L0IC*��i��&ȼ��ӛU}̹@� �A$u�u��br6$um�>����������g�Ao�jڱӊy����ɰ�|��y����e�,���'�E��U�W5��ϸ�-��L��6y��1kM��{�u��� �
�?�j�z9����������w�9L��?A�9}-��\�wv��H�����Bh��	@,k��bF��Pr�j�4�څ� �;w����kgR�r'�����2�K��������V���a��,j�?kʹ��-��>O��d��X��b�d��Z��U�ͽ��L+�m+0##5Y�f��g9�xsY��m8�9({b,�<7�h(�7^\����p'Ɩ��d�]�ȗE��P%Qʄ��r=Ƶa6�_��TJnX�d�TPBG���K�KjL1��n��q|~7��F�g��:c��	�5^j*�5̙�{:� ��A<�p�P)S�|�HEW'�l������H�F�P|�HK�*g�9
���+���/~hLD�J���5^M����q��{q��ژIp�t1�*�����E���"�N6i���{Q0,� rƂݾ�o���K�oy�}A2ϋiR���DuL��k^8+��En�Y�~I]2��f��v�{���������6	�y7~;a�T{?$MmF��~�#P&�n:,�����%��E��9�i^C�z����Z48��\4�@�n��aB�"�'y�ܿ��J��-ڧ���vQ���	-%s5�S����27_�H�ȝ�W[ݣ[�U�eB��k�P=�� ��}��>ѝ2m|������c��4cTV��	,��֜���nW�b� �媘#�X�� ��\�;�/�ΐ�jc%1( � H�Y �Z# hm#�B� �B�sA��h��4�ۦj��Z��a���8���\�@+O2@oP�)x'$oH�DJW��
�8L�j����y�m�I����M����b�U�����K�#���@����`��xh帤B PbV���S�x��k���c��wm��}J�� C��y�a���e�E�D7��^PX��v�ˍ���bm[�:H�;�{�U=��H��	�8G(�%3B�+k�9���59��Q���'����X��gY���o�";�cb�o�31�_T9����MŒd�K�XJN_�с]��v{���߫� _T���2��,Ni�%��խܪ��l�g�ܒ!P��xx|5�;��H��yl���/����"��f�����煊)^
xx�[Q%���+�&�lV��V,)3[�C3x��S�؉�0o 	��p��6p����kg4R������u[�x�E�N�غ:$�3Pl�;~�o�D�[rG=qZ��t���E1��BB7H� ��"������ u����L���{��|�jv�'�� �sU�}��b�*�:�dı��B^Y�۽���ݽc�(�1���ʝ�Mۋ �������,��3N�ړ�{��޼~� A�;u�ԭM
|�h� �%?-e�Q�/�Yls)�E���
�(���vz��X����ew*c���lr/�����O��j�����2v$���B���X!��{�3Ѯ���)icA/�" l�ٖ2���V�w��Nd\%{mOݳ\�1sJ|��l�����������Xup�R';��ɯ}f7�|R.�g���gLD.@"Ck�0Z)Tn	�D[�lA��n���nT�Uq����F�-&�5C�g��
���2~΀Bĺe�Ahr���Z��_j*�f*�@��l�TZA��6�l�����Yxq��E1#@Θ�옾](�Gu{;e�g�V{�ŹA� k �ك1�]K�^���w^g2V��.缆,��Ш�`���} �l�1
J�N��E.�B�g����� �����D!r˒O/p|&<�:��h}�A�^�Wx>�d�S!��H�{.
jC1+��.�C��</~�\�^�W�c����kk;��V>ǚTS�&��	�k���Bݫ43�r DpY��X�,8�i��3�4��e~��ː���U����+�GI��{j��	FL"�%jK�H&5���I����Z}�,�� ����v�L�R(Նf?�� �̵��l������
 ~��M�p�B2X�V��ZR���DBx�Ñ�ߙ>ӢZ�9կ�Y[VA��Ce�W��a���%�����ʠ��_.P�VIK�Ȋ���ɬ��vd8������ƍ`��!��T�-�5�n�Ե�c�T@O�K M�|��`�3 ��� ��
�{ܔ|��V��R�kP;@�dx��L�[�V:��I���q��t�3�I�!�Vv�vi���Y�o����t��v�r<� ��R4-��ڌ�XP����B'_/uQ'jn��p>�V��F�y⻤�/W�P!a�)`��Ey���$@W16M6lms�6v�E�u��[�<x����l�]#�	��
cq��2e �?�����N}�(hF�In�ƖpF��ڨR��0��yІ���Ö�fYq�!R`���d���Eg|���)�>�h�i�7(?����#�b��pJ�����vcb�ww�&�HL�\` 
����+�t�g�QD@<��g=[��ѕ���Ԓ��f�yV�ohH�i(=8iD-O��(�ܺ�[���N����^�G|h� ���&	��>9�e<Dk�h]� a���{
�Wtcu�X�-�7v���f����Ȯ�<�P��o�-����[��Ц��U�ٍ��i��"�y�Gƚ�"ٱ��g����P%�P�_�$���6���7NE2��i}�P++����
�M=)�m�D�`ObN�'	H�:����w[���:7z�I�Ή� �(���d��g���薷�hc׷7����Ҵ��W�y��1��܉_[��TZC^��Py{��3��_��>Sh " (�P g�^�L^��E��"���6����Ө��
�&�UJ�Y:�~�����`i��]���6�^���r��I���Ye���!|�{�՟ښe�������U�E=c׹��w��E�dّ�l�E3�+*��Hպw�K������W/�t*"���n3����#�{� s[h�˿��^���[�g�*�,Pt.�e=�,f��`�`A���}�p:7�-r�$����1���!T�,U>�z7q6�vˊ9�<��!D!��
��v�R�D�bC춷�7�u�A���$�p@�~���Vs���(�Pw��Q��yN:'�P��0F�6-(0���,ߌgB���2F,��Kjn��N�q�����y�B�����MB�����t�8D�����6o�`c�5i�,XB	O19W�F��D�o��B�l��Z�[�* b ���ns�l�.�C��=����rS���Uԭ�+�zzb%�Vz,Q���SV�u���P�X��:x¿ï��腇*6|��hܫ.s�vF��s	�-���HQ:[6Id�FI�ѢM��Jԏ�k�^diƵ��%�lC�Ұ����P�]��~6��t<���.ޤt��lL�a]�R�!�
��¼� �ƌ�o�B:�ld�U�Qƅ�����q��Ls�j_P����|q���V5�<�30ȋ �f���A+Qͅ} $�E�Ճ�<[��*�aT�²pn+��o(����Z��'yUdhI�IOI��b)5)�j�|>񞣅OJY�T4 �o��R�H��B�.�,nl͎6�&2�&?>1��P�$u��50���� ~���C'Obu��2˼Q����t]ū�H���v��Sh��9��2h�b@R�At�Y6t;8E���O^(nH����D5���%v��ͤp�=�c[�t����=�������{�%, `��N����6vl��m�xúb®<����m=��K��댾qLP�+k	r���4��ҁɨ������$z� �(E��Ü��sK��e;^ϑU�Z���!�M�]�B�����
��ώ��i�V2����ß#|�>ω�&�G�mn���6u�l4�|�,E(Q��}��rPۼJ�5��;V���ص�%w��Ʃ����@��Zk�d6�_��鷪❃'O���tN�L��Lf�� �<N��^��~���	|0���#u�Z>O$��(�Hx�]��^2�{�!��:y��!r�4����q��;�޽欒�y�(�"�}#:R�h��zs�D�M�"�#�B�������3ia�>��#Т�Һ�W�̄4��h���,���,(��C�f�
�lv�����9�f�.�_a�b�d�R�T<%|��Y�cĨ���=������?�O?�h���?�O	�1{��110����\]��鉽}u`�?��^�|n�?���*�A`g	6D�ʝxZ+�3(蔩+/5Q	�4��{�K��_������Γ����T<�=��f������|Xi?���� Z=y�����d��4w� �ȋ��T-.�������{��Z�b��UAUsP�������Zv�:��7-��h�J�T���b"w$
9H��,(���H����F�^ЇE�$s��,�OznW7��&��3/hr��;�u��4��9ɠ�=�5B<�Z�SpU˂�WJ�[��y�-��C؉",E�hA0���LU�U�� ��<g��Ѽ�����4AB�EK�f��R�j�y�p1{��g�[ԭ�P�������֜�z${�M� �[�<��h��5`���dX �s9���BL�$�ٔ暖;<[lA5ԮM�t	���AOӖ9#�%jI��L{]y]*8+���`�n>;��������D*�oX�\���<�3��d�����^`O��A������0	l�nY�kK��rUׅ]��Љ�|O��&�]y<��4���z�}��+�j�Q�7���[_Ѵ>yN�g�'��w�OcX��THOp�IE�JP�m�l�����{;�]����9+�H�m��M-<ݠo �Z4I�ܘ��='R��R"dː�8��N���7)�T��A���{asSU��$��;::����{1s�S� �ΖH��TCF94�8(AB9�Ǫ���^��y�����v?3��ѵW��+���G�-yQq����ȑ��(ix�� �b�U�y��b����1��"�-tM�
=��+������ȥ:5�B�y-0���K���1Ԓ���ws}��u	R��mӯ�����5�@���!tUy����+�5����p�ٶ��;`�l�w��s�rϕ:z-��[H�CrA���[I�z��[�B �!�)TQ�'���$�t!W�����48
*�kVN�-��(��3��yl2��W&Jב+'"i�}`9��97�)% �Yl������B�fE�T�6� �2q�IcY��Ƀ��u�ڸ�;��4�b^���~
�$�Q;�J.�	X�y���h��^wI����[��jgg��
����L(np��C;>9��"�X������墭U~��l��h;�\�5.�c*�dN]�T�V���������0&{��B�9xbÞ�w�ۥ|H@,՟;Ju*�	e��U�;Ո���}h=1N��՞dJ�\���z�g��ԥ��Ү��������)
�7]��n��J�� �RB���T�����|m��V\�*�a�v[��X�H��s%����	���;-����~/�Z "~�������f
�{�����>����ƶ=��k����o~xj���k뛢�jGÒb.�_E����{{�歽~��^���>��[ؗ��7�,}=$0�Nk�����5�5uu0!�}m{�%�ٌ�q�&I�>�_���,� Q�����X_�T}��	�Z=˯��</���;���7Е�����P��X�
<9;gk�@8Ո{�g������g�@L`ڀ8��L�
^Kqj�--Q$���m�{27��D7m\:��c�����}/����X :׹��Mڂ���
�,T�N? ���Ǒ��)������ǿ���BF.J"�Q�3)�"�4�4KK�\4]H�K���E��n�Ә��Pޑj��S����A���g5[�KF�
���(q�9����XH�/N���t�9���t2�<0���oEѢ���`ɼP�u�V�5Ƙ_�Z�S�/�9�;g�����Gg�����!�SQxj���� O�,�E6���\��,�u�L $s����*u}���]`}�k +%���TO-4u������6���w���F6\�Ȥɐ��Wb /�o��wNO$�pFW:+�(ҿ�O�1&��>���]�!�2������.�U�U��j��P��7�Ͳj]���ne5���	硲λ\�QIV|��m^����~hM� 97 :�١�&m��|(���2�T�l�h����7�.����c����f����h2�����}:8����xmH*_u�(C=�+������񢥭�i�A�|dɠ�u��R�$=Y�w�J�h��.��2zcC�A�� ���!����/����  ?]]��o�c[�3a��T��Җ/L\#��>o�y%c�AE=WVA��p��Vh��y4�?��\xeC�����ۦo�l�|���Q���f�Xݨ�a��%4��(�Ӣ���
�p�q����9����8��G�x6���f�|6.�a�Ǚ	hc ה�e:���@�B�0(�]Va�t�z��uҺr�̕����\t��PG�ƫA4[��I*��cs�5h?�U�Ԙ���@4R7؇��^��3U�1q͕R��R��pZC�I �UyOP9��͕du�J�I���R)�KX����l���
�&������1�B#tT�j�.��2�^A�����U��lo�xܨ8s@@���BcG�17���.��B?7*���.��\�D�h��(=�L�ݫj��݊�ȹ1��P0��ʾ��V������Y*�b���#}���|��ÿ-Sw�ݕV�Uj\��I�9M��`��I��ř�-\Y�d�sK��~-���z�=+;Qw�Y|�@+UUYl�kW�3O|�^�֞��;�ijn��a��
��0��D*�P%���yփ�v%a E)82)�y��?���c�k��I<<��f� T��:��g2ٝ�{���}��m��V�g���A��\L(���~}�����?���};>:���)X*FR@�sC�EQToYs,��9�΁�KV�G�{̏Z�,unbJ�ThTL�<��r�	[�h-AU�[��T����`�-��}�x��7:Ɣ����/��s՝
"dj8�@�Jz[��`q�ܥ�eJ�����j�j�W\hf=�Ra;�y���?���y�b�9����f]�ʒ�Nz2�O~�dGd'�W�g}Kz�y�)��I�U�H/�*��.��`R8�a�7຃��?���?mo�,I���GD^磌o�`fK���R�_���H!W+ >, � ���ޑGD8]U��#���jVvx���e���nnj���-G���D�}'�j���}䌣�������O�}�ڤ��or�|s%��L&�6��Z���r�)�� ���D*!�٫����=�^�W!c�'���X�I�M�)G��(|E|Ʃ�̔�� ��;��mR|��cv����SfUy���V\k�M
���
��DZ'�a'=c�9>[L��L�����c��V-&R��10>jbZ|�S�����zّ֣�}�I��F�ɌS�s�}�)�֗v����"D�ru�v*�:U�-[��s¡��0�F�9�|��J��k4k�Cg��Y$K{E� ��r����Iݣ� W��X�gP��veC���|�|`2lX$	�]�Y�xR%E�"*n &:���P��ۭ�'��5��O����uc������k�������?��_Xwc����)jԮ �uw}W���t���(� �IG#Nz�v�+�J3��ꢊ��=�9Ja�~E�bM������.��`���t.��Qe�Gު���4U �(�Q���!�Ū�7�*]��ߋb�������L�sv�E'ǽ��ҹD�k������%qёh�X�b(�d�I(�3[3�I�6��{���`D#'mR)9�iNH�s! õ X�C�z}��"�^�>)�$�o�g��ٶN�(T�� �w<?�8S���8wb@ �8�{L�yP#����5�#�z�F3ȸb���g�XO��<�X}N� 0��O�|ql��bXbe�zF�@H�Q������`O��ax�w�(Z�����M
7�m�� ���#]故g�([Y��큨�GJ���[�mn�5��	",��d$Q,�^ߩ�����[�� �I�R�d�7w�D֖���6��'e�P4=d*�E=P��)�NmA��������m�
8j��������S��6�1^��_'=/�����C��)�1��p�!�����������.��æS���d�*��i�%�+�K�F��arvAǤ��"v�x��@֝\ۗ�;/ڴ�Ӝ�+���0�:g�<�!j���h��l� ���zr�Z���׬��s�r=אTƀK'0�?�վK�2�&�{�r�k�ʑ�,�8>�KIQ���v�Yn���l����u�G��+�kkW�vv��Mk��A��do(@�o��������X��A���0 m;x���(�6�Xo�2�B2��`H�u5�w�Ξ�׻�sv�猒j��-�W�z��s�36�Wm0\�T�>�M!�m�-C>��x�'W�c}�טFC���xF;�h�^)#M]7I�oH����X��v�S�wa?`M�I�k�\�ۈ������%0pԆ� |��P6��.�T�XmeVE�Zr�����~����Rͱ�ɞS�m�zH���
��#��Ҫʩem�h;��@`�����R먨Y�VM�e��iM�^�)J�g_SH����0|���G��c؅���[oP���%j+0"�G @꿦����k�zx1�({�HW�`���Q�X�1	�@f=e����P��"pa%(SY�e-�Z�|$��֧~���l��I�RD�ߌ��#���#��c�AP���/VCeE08[�uV������Rd��3Ɇq�8�q�g��ʘUS:����zk�Vev�
̭�A��
��a#f�b$��=:q�����/�P@3�C����,S5@?�|�Zso%�랤����8�uҠ���<��9��?�00�fuk��)�a�0L��"����u�Ϡ��S�;z]LI4S]̤�-��i -�Ĭ�g���~�YNmX���"B�i�!�ȘR�s�|����䲯hR⊱@��0���ۏo�������!8�X���)�ص�� I%o�i�^�,�=�z�j�D�`�%��� ̛�;���w�s�y��h7�]��k����;j#��H�,W����<�%_�eO�����=�U�����&ё�����F�4S��#[���i��r�|b��O�O� �"�:}j�T��D�FO.������(� ��isQ5���x�5x���V&*�<j�N�T�~5���؍2F6�fb�\|U$�]Osa4�$ +sn�zbl"hS�4�`7�PF\�{au�Hg̟��(��"�Y9n�N��="�&9�ꟃ�4��#k;!�MZ^��E�c�������\9kV]��Ƶ=�7}�5L��"M5������ϼ�472o����O�ZCP��l��:6#�]zA^D�:�����ċ:4>�<׹]#a5:f?��g~b[���򷸆�{����ϡ��Cnv>���'�8��g�Η׸����x�dE��Q��3]L	&9?���	��T�QNqi�%ې�ϋ���<��F��g����=y�߶j����;��e�E$}�����Y{�o���~�����/��[l9�߿���������~��?�Ͻ�T��m����i��bM�'��xr/@���٘e�y�fb��#Hm��Ž�|<���E�t}r��O��z,��.���^����[>[��u�P	Fܐ��T\+;(�,r�F���կ����(�X~�?3���g^��S7K��j��g���; �4�1l13���f���t��Mʤ?;�?9���lSd�OT ��	C����\�'u>���"cs��Ge�HIC@XW7� �3�V���0M��O��U����E"���,z
D�����Tm��6�5�a�9�L/}2�O���3 
y�����AQe�E/5�)R� ��o�}B�`�i�<@HTE�F["9��\Ԇ~rY�U�^�d)���̖׈��k�g<���z<��9��0|��Ӥ�4���� �k�,Ւ%e4��1���H�ȜYͼ���Y՞0���<t���E�*�&%�O��=�U�LNݯ�d͵.(/칥8�����3�ƥ��߲"TxHkQ<
�6�n��;���T��`�ZT 8իHV�u��c)X+����v�U&4$��?tkz:ԟ��)8$���
�\�TĬ��BK��'-t!��5׶�����If{E�&��T�8��zj�o/d2��)՝�N�q�3���H��$ղ�N���;͔97�]��{�X[$��T��4�u�فP\"E���hv���SR>�ፙ��B�skq�+�����4��:r�'�uAa{�\����M���6!�h�Q���+��U��v5���T��g2�f��dvG0�gtI�Y3d�1�:� �i��10c��� +�2}��EqN�[lp���5��<��5�pi�u�M̭FuZ�1�ٝK*?�~�=`���x�]��s�E�������HC��	!6R���R�QOHG�)u�MR19h6�ZN�>�K�.u�_�
�9E�&Q��������J������0q.j�\�a�i��Z�E��7���묬ii9�z���������g�/��g���s����Ի_|�=xF��s�x�����>��G��'�{��G[ 
�����]:���vm^��ȎhO�1�!hBT<�(ȀpG����{���Y;��_�zI�6����ho޼�~��@�_��_��~O���(A��5$�s�@��v�1��Ͷ..p��go6�.>\ip�︽��+����#�:K��u������8�,�g�P�z7�'��3�(��
ij�q��k]7#A�d��)��ҁ���݆z��N�$�4^�#w�����!�5���m�~UP�[��T�m̫�v�ⳅ�h��q����
�۪m�)��u�,�� QB#���g^'Ē�QY�[؛���Z)9��q�w'�%�X�f���Př��{Qu�q<1X��g�޵���tcˑ}��%��^{G��A�h�-;SH �%0��x���%~q��}B"0��@3�9�±��d�t����Hy��93��"^'�m'6AU�3a��h�C	R�KU}Rܑ7J��+����ԼA�%�`�(zrƐcL�W�;�T(!b�NN\�^�y ���P�$��D�G�6n��
n/��4y��̬��=d����U�_(��G���h���6ma���/��jG|����Xi��FY�+�Ȋ�\j�۹0;�V%�7��u�R�֊�av��#�B����H~�y��&%�����%OQ���A�0N8��T/֭���&��Q����t�,n�Vl�����vs��hvW�{��˶�=�}�q� Y���B����8� �49�H��W��S�U��)y}2c����C��qs�T{<�&��@ƍs{�> e�-��W�W��l.������q�U�Z��Q��nȱ�O0+�բu���cS�����)���{K�0wF->���E��6���A|�9qi^_(�v7/�����+)u=K~Ur���.dd�,�)&�H�X���zV�+��)s��P�n#c�5vk����'����Sn}��s�Z�e������It�WA1
��aa�$�c�ؙ��k� 
*XD7�%�r�JZ������ĥb�q�������ДWN+J�� 	�!wڬ��<��s���s�e�;�n�_�ܛ}6y���dV$�*��C�����|5�N�[e��k��PNqvςk���g޼�f��G�����V}�O�:�!�� Zf- cƽ|��*w<���+��� ���;m�`SjASk��������i��Q^�0/�\8�f�����]o;W����ӔЙI��P.כ7?؛�o(���YP����]b�߽'�B�Vʽ؃%�!n�+�{a'ڝ��ٴ�����mr�s�e�-������;���������\���@V �z��t:W+�6p�L�Lo��Դߪy��ݩ*��̝�Pn��g���2f"���;]2ۃ����N(�����{�hR)�y�G�K��
�(��#�����̋���A�ѳ9ǅ�*���k�����k��|52�5��ݜ�sP��HF��#��x쏫�������9[bd �{|`�I����Ȗ�iVe\	���$�]�l_1��k�Q~1�^���䇝��H�E��#�j�P���dj6��Y5��u��T�vr�#w�I't,�����
A��T�t1�KE�*k�G5䵠��[�^C۹P�̹ĤB2�;&��aVO��J=)�u.n�� ���T[/1 ��[I�q�&ܣg[�.���f�A�&��[������	�hF�wGe�n�����۬����:&��V�-�bϰ�03I�c޲�
��.H��H5��Z^%3(U"&�{=��5ԩ%"$�ԲcA=���UdwAQ͚��Ԃ���Kz�U�B]׶Ial���1�F+Bf��0f^ Hq���pFCݪ�į8��i&Wуwy�ot��^�R���Fk}�0�٣.�s��$��[v�Ao�)�jy $��,�\���ۭ����}��o�����_�ۇ2a���g�C�i����K���1a�Д��
��5��ip���su���<*!�qk�9 �dH����9���ҰβT�p�;yt��.I�0��|0.l*�ID�i�AQ��5)�I ���2�@ga���;�0�l�|:�gE]�P�	I'�O��U��wG��8'���b��B����N�`+P�1��j�[�Cwò7 \cSX7��!s��8sU��EA@v[Ef��%Zg��p�e ���s���M��u0���
�R�<��dN���A2��A�1�"��~8X��:&�VFv/��y�����_�M8W��̭���M�FeJ8,�䈙��*B���M$\8�*R���V�'殮��]1�-i��E�����sk�}Nc�]���}��t�����>��{EEǓ
ֹ�w��\z�\t��%��:A.�`r*h�"�a� ��<Z�y�V����3rD��Oj��k�yog�ds�h}.���۽�p��G��#g{U��-��g\`v���JV��
$�e�)F�=�ߨpf�?^�\%�۷��B��hZd�j�#GR����n�*��3g5(F�v�S!j��/|�N}�G�iV1�0�����|6�IP<�_��\̿�~j��8o���sj�:���@���k�Ώ��f����x�K�%�MM��;�F}qZzo��z9��N��'�E
Ĥ�kD]��L�Nr�P���<��vc^�|v���qn"b����vl��l�c%��XZdK9�T�h���ՂM
<%�u��fr�)䊗�C��*��e��o������?@�
�A�����Y.d�)��l^�Ns�j�$|p0\3X
(���_ �'J�r.�A�$ Q3y���>��7)�� �d����Վ�j�ǲ��|A=@	��6.PK^�?�S0���p u�s�Qv���5�Y��+�ӓ��Q-��xb�t��j��5��jǞu�mA�YE@�wK��RO�Z0�a<�&�'�%�f�X�a.�� )t��a��/W����ؠ�X�ۼ��M�w��A�i:r��Xx��]^�Ϥ���F�]��L�c)�����ڋ����k����� �D����ɠ��d�ޗwt-Q��$����xYI�5V^��j��K8��]�򵌾-^���I�B	IAR����7�3=�{E���������<Y�௧�2&���R����(��>o����fgϞ=�HYC��
�����&iP�+;CL�W���-���@��/웿�+{��/m�{Ae��;8d��-��ӱL��mn'�ٌ�5��>R8B SD��"��T��a7uɓ��,i\���H$�9�P���(xpEGDA���y����bD���HA��+�h��u��4[N*0�C1�� P/��y��)����q�,ea�p�Y�x��l-s@Ys���1J����37�26+(�ាW�����g@fw�UD�2�rW\��rp�I<��� �A��P�A}�)gEh�'i�}0��W��*p/ ������ۜw?Σ+'���*����Ξ�xn��w���n�ڣY�w�?>z��Я;�
|x�W��f/��S��5���_=|�q�\���9"1yDF�����*]��tϙY�#���lz&N��C`F E��J�\�:�<���̥M�;:8�r]�~�A�kNn3J^��S���e��'�Q1��0�[�lxc���,ݮ��l�v]=c�%6������9���A�M��N��h�o��Z��`�y^|���L���T�t�ζ�"5����c�$��Y����N���!��9�\U<�V���f�,hRqm��\Y�,� ���9,i|�y=��>sVϚ�G�Tg��Ng���-�.����^����ހ�������;	�DNU����p�ϕ2�!�A�t6�"r1�L�%;���s�/2�97p졀 ��W������$:�����)��x0��+��p@��D��3s��h,�gg����F��8>Ɂ���KD)��_��,fX~�os��7��MN'"5�����'"�r��	Uf�D���:?���T{�1ɋ��Nv�J�=D"��z١n
��-�ǘ��xKL��u���u}�S7��Ϊ]�T��]�pe����|���32��;���"�j����^�f�u��>1�����T���H&P?�P�.�����3�m�o������J��@�����+9Zd��6>un���X\��Nc��
�Do��� xD��T �t�8���\�^#ޫ5H�N��������U�%�Ѽ��sA�v�(����i%��9�@��J99��!R��mqm��3L3}N�i�0��������M{_qG��Sd%D��6������6XWW�
��w�z��&��3�e���I��i�s`�Z�V����w��Es,����Yd���2����]l^�(l�M�,�r��� �2�wh�j+�$��Z7����k]� ���򝫝;*�= �O��T��B�)���/�/��/��=�ԟ7^��x�ۺ��b@���#M��_f���=���io�2�o���bxo�������{3ٻ{(��6wW�� D%�mBF�tl��IR�µ�/�z�j
���:��а>)n3����]���dP�]5��L�5��,���ɉj(JQ��`z��J�|�ӊ �&�bKk�c[��~+�q���~f���;@����������S�� �b(�g�}ԥۛ��l�h6�f�Ã;xƨC7l�oh�t�e^���bolDp̑B��?m��I�퐓�.����
@���� ��XΉszz���,C�ۡ��m1l;H*("���'���,�hW���;{��x�����ʘ����y�փfڌ:�W�S�DQ��X�@'��>�� ���z�΁訩�"��٥4�d�s�E-���.G��i�)�����#� kf��)9^ �Y���)1���C�:IR�^R��sP6�t
IxDYy�\���6'*@W�-��Q�1;�_�,8�ľ+ �xm/�������[{��=�{ε��� ��tĴ��~��)TO��^�t��I���hy�z�;�����X���l��/G4~����I������g��.�����vȸ� z�v�#�~H�K��M
�$���$�Xl'�똝
���%��˃��#Ʃ�$���^���½N�#Nu�_̏Z��.��N�����֞C���=���� ��7�6(�� p��:�et*��Om��_>h��+��0�F/��'��mR��j��I�J�Y{������&���\
0-�kQ��;�	G�l�m�B)�}�Z���.W�IfG�{�-��6P�-Ӽ���Z`�2��7;�Q6ux����<P)��m� �u��¼[��KD�pA@q��:;����+� �O^�L�N�a��@�Y���ű_��N��9�$[�^B0S]������j&߸�J���@�s���dO��A��R���Xs��\}V�lr�Y��k�?`Мz&�&�F�k���vp�ՠ�=����g&����wۖ�;�}�̽裩�$��� �M�͠����2��HM56����]I��A�AJї1ڋ}4��a����sxν��g���HQ��[p��� �!��b'��צV�*0��٣�}�wuhl�%���1Ze�NK$E��Kվ$�A���=�bQ����f�c��X�-"rQv+&���}Fi`0�>MN�[���
"L[?2]*ޭ��G�m 0#Ⱥ* �v�4��~�%)��.��(7���˗_��_c�~�}��7���t��G��@���x�=�=V��T���U�I�Rv�#��������~��#RKA�CY��
 {�)&[:��������V�S�)��Fj;��cT�5�s�l`��qH ���r�l��젋i��v�N��U]8x��n�:��g[]�&�ƍ��#lsv>+�R�
�G��&�u$�̟Ԑ8�e��~�H��y� �,��?둛ǆ���]H���0�W��"�{C𨨬꧘��\��ρ��=b��)��AO-��X��q:��,��(�X�'�����P���p86�٫�0�]�{ϟ?g���@��:�;�w�>�7n���ݕϾ|������k������L& ց�5+�#���Lg���e��'V�[8S2�s�M9�-A憔�]��2�;��k��'�$sڐ��C�˱��T�̞�'�C�߲}�zI��7�H��Q��H�ȳR�z̭�U�ĺ�B�E�I��S}?�c�׾���܀v&8d��O'{�?�����=ج��n���<$�a�+ �S+P�+�%�IǺ���._y룯0��z�������@�Oͬ�!ռ�U��:����V<�vꏿw~�t�>���|�O��_k��KT�<����Y�|1t��ĸ}���;Ug6�M���d�a:�JD�W+���l:�׃zh�<�{g..�j���6gWi���Ƃ6Y�z�v�Qͤ�����I_M��뵜��zи�����A��Yu�!o���D�%��,N^�� �)�14S�<��锫�Bn�w���.;{$<[��P�[������;;C��}&�cQ�1{�����Ȭ)J���QOۧ�v7JFd�h��l������P$Y��U[P��Κy�
�;-մE�S�� ���T�{��lQ���݁O9t�	R��>����}LR����'r�X|%(S7���0��H=O�}���Y ��I2%]u�5�z���t�u- ��q�xn;W���.uފ��10���Y�:��|"y�H L�9����ea�u�>�R�i�AM��{�A�����P�`����ծd��_߰����&�� ���y��ށ���~Cj��a����Z���byv��������!u)1/lpJ~?A�sP��ޱa��}`�lq�fՇ:OV�o����|ɧ
��4�v�ZÃ����M�v�0f/�S�T,
,�pN4�D�3/��H����残�y�#
'_iH<t�������7_i�~��}��wd}k�w/*Ț��w��P.|,N�=��gqh��dGr���?�*�
��d?��Vbd�`�z?��c����[>/9f�8���LƉ�~v'���1��N�P�,S6��8�Ң~r.��#A�����C�c���~�s�(TV֞*UvIY��
�o���C,�S�:|���zokY{���nC��g���B��咱O����N��n	�ny_ ��N�Ll�!�(�ON�ڮ
Ⱥ!�rz!����w�1�mMdb`���ܼPO�r��65���qd��=�	~�
hz��%�Ώs� ������Y�o�kzvgϞ�( �e��S��ov��ᮜ��LଞR/�����vwbo�<�����<^�<+cvg��mq�n�7�j��&���>!�6�[��*t�5�FD��NRD�u�	 ��R]���.i%�����\,�X��e\����H���5pf5���0���,���׍+'k�D?�K/�.��Hq� �Ź*nW�
g��h���b��0�5f�Ԟ�� �g�R:�ןz����̾���{�ϟ?^��K�Q=��9W���?y��?����:���r�5ޕ��/~p5�#� �-��/��!,���j�A���0	����
d�]�7�%]���u��;�qOK��H�`^l�5��mԨm<���.4ڮ-�Vd�"���[���.Dp��N��/�Z�3V�7����>�۵^+�ü���U䮚)��� pZ�Y򀲟���3Qcj.P���b�c�w��р	����β��/��@����y�<��^Z �L���^������ ����T�v1�����$k�lk >�i����q`%�z��0��t�RY�1�+�H�p��J@Q�ʺ�������|�0Z.P�Λ��h�c~P�?���Zqt�l�F�~����Ĺp��7[�W���?<׌��խk����H�d+�����td�����_$7�L������c�iw����-Z��m�p�����Z7�q�z/�U�T�����C��d�A�2}����S���U��,��~�8�ގ�DA���^/�J����^�}b�b�Q1nؓq<��a9{}�I"�2�Tx�m��\E���OX��VkR�y��`���vU�usn��ŭƬ��ӼTLT��#Y����S��R��9�II:_Dѣ�}�I���B�H%�T�����ݭ�x��^�,��g�]�))�p�z6�S�:��nʈf�p�+:�`=�X0
���'{z����@t�z�zEK�ѝ��3�Hg��O���>��w�h^p��=�\�<�B��M)II��݊��)d(�P��KzA�!S�%&�2(���*a��� I@6���QF-�MZ���G���	�"Gm4XQ#7�A�R��Mk�е9�{^���]��@W�>�.Ȉ��'�6Di{Ei��<f�v  �,E6�:"0:�Y̓2�jȺc!'
x뫲�MM�X��"�5����F֯�����^]�ٮ� �	L��5�����C&k�-�qs]����u�ke� K`E`{$mT����&)#�u3e��${�fE�������[��67̮�@�8��˹x�j��H<[>�4yF�'I>
Ի�I]l��H�GJ��<��-��e
�[E�ݩ�1�5H���ò�1r�S�٬E<(G�ӂ�d��t�q�S=`vlveΡ���t[�f����ٝ�.θ���uլF��(`>&���,P��]B����g/;��s����>��~�;L��i��Lf?��\ljէo��^��w�����g���/qAG�=�|�
�\f=Z~1 E��A�yE���g"�}X�Yjm��Yi�y]����[�z���#���g�s����\]�H����R�.�Fs�un�α�:2g�� -�������� Z:C�d2���N�L��s�<qo��Fuq�X�<* ��X���j�G"x�4E��k5�,C�g���ڭNm3j�J�#�D
>!�xz�����&�R0]�ޅ,zoi�����}J�}�-���H1R|�M��,���G��܈;�����?��=6hg��9�R���s�z>��;9�a'%��m��5K�P�2.���l�������N��r�ͤ4,@BeK�Yw�@��H'ͣ�k%A1��<�����q��G��3Y~��8Ùo�<�=Y@�:)�ާ��x�2�������0��z�A�t�}5q0�N���e�{wb��<j�����p߇`�@�CL^L�uJ�>?��_3A�gd�YR� C]��;�T��us`&�,u�ӑl�W�Β�)���p$�m_���n'��]�ף*��x���^Dɪ�\�}\�5n�����s̍f����](�������p<GM�����7\4����L^��	���6Q�`��O� L�|Iq)IE<�t���ŉޗc����6�i궶�wv]��wh=n�
�eϡrΡ�k�u�.I�vN?(�= !
*�=C���<xd���7j�R���=�M� �H%.*U�̥.�����w�נ�mxm����kMiW��G�W�E2�7�~�y�Qh��S��H��B)����Q\b������0�JiԚS'�"i�T�[W�S�lX�Ź�g���X:4��%�Vn�ۭ��r��o��1Mec`�o$R�n8��#� ���� \�3�^q9F?o�x�(���,#��^ۦ̡�>S p۝���{�~� ��P�c;PM�ڦa�Q�r�2��	�X�8��6W���$g
����D����܃��W�bad��0��n���� ����h\�w\/�	I�e��:��]@YX���M'��˃��7g����8�����3��5&Fh'�0/�I<�e����)QO����'W]LTvJ4/8J�B#��O���M,M� O����h�IGEҮ|��ͭ}��}�ꅽ|���%��M�G;==���H�e���(g�5�95KǴ\/ a)�G�c4����-��y%�o8;���v�~�q:�B:��������p|n\ �������>14]Z�F~l�����w��lI���5���$�p�6{� 2����
~?���̩�(F�-��)��
VV���0��M�Bj"��mM"Z��m��[�I���;��{<��%)q�g�ӝ�����Ǧp㗝I��-���~���ھ�۵X��˙���qfe����Pq�1l2�����d jѓ���-3`_`��Yg::�1� ���V�[K�0͒�~8��Ԧf&O#kU��Rȓ�agI~�N�E5T��3ީ���M���XEy*T���ݼ����yPxhR���dU^�)hif�?���Ȁhyʧ��=�~Mp���$�:������H_��{���\  �<���x{�������� ,ڎ`pE5����6"�X�`�(��D���X��SW�-���
��܃�pwؗ�R{�P�a���lPڱ�o���=գ�Ⱦ�����>��h��{b�,Ir�X����{�L����P]r���,z��/�p]��r��J�Y}�������vf�o}}���l�O�>�����wq�y�]���P��u�*c��(�����P�~~�^?������,�_hs���E� +J�K�m'�G������I͐�?��؉w�{�b~6%"(W?����Ԕ��{��y�
����0�lo߽!Ȣ������X\�裗�>2�� rv(��q�T �t"(��y�\Z����������=�`.7�e�3U�v�
ߨet���9#]r�A�Qw�DZk,�a׌(m�"�5�8{�P��A���v�Y�qC]_�pٕ]lS�:��j6IWF�D�\l|s�����˃�����ӱ�*I��r�Sg�(/��A��_�$�[{�?=��͵�_5�c���l�Zd�UZ�ZlLtx�P��G�~#{��4�6�;�|f�![��L{IJ�#�?�����y�!�6~���6��2����Cf�'X���������$e�X�"/pVZ|��K��2 dȠm�͂�:��@"u �0
g���]�v��<�_,RF4�S)j�5�e?t�xY�k�F2S�It��T�M	�Y�֪��s�����*	��G� N�ߘE�$����h�g��.�ʎ2��TW�&�u�4���T�̍R��h����ؾ���j}�5"Q�@P8���8ܒ�E5s���!z���pPƓj�@�d�r���&�Z��pJ�Ήt�x�T�H�P�87W����s��/�/_؋[Χ��2�'H�&Q6�*M
�y��J8����]ʿ��|�*��������Ws��y����k��R�)U�Μ�s�1���wlq,���Q�q}�� ��D�x/��?�:S��@��YÙ��`9F9�����u���QZo����q��E�G�NB��6��I�
g=%l9���b�xr�R.A���@6�k�Hp��u������D���yt�Hq-)T�� ad�:�1e/Y(c�z�eI���y�L����=���mI���2'����V��J�������C����_D=S�k��x֞�"k�$?Ϧ�����X ��A���,8Ȥ�N�T�.�6���j�H4��j���`.�8p�R'%C���8���&��s4J��G]4�^s� !��]=Z�z[Y��4��P��~�Ϣ�ʻ�O�zv<ef\;��؛VL�L���=�2�Ȟͮ��uJ=������	,���&��Ӭ�����,���"8�)�����ww��ژ1+�':�IA���0(���Kh�����Ʃ���n~~Ro�Թ�L�{�=s8��G6�ɷ�v�ѯR<I��<�W�-�S\k�X�]�/�@L"�dy���};�g������Ld�<�0�{ �d��� }6��s�!)��[;�8��
`-~7)�ґA�����.l���l�m�?���mKչ�(��o�̃������Nj4@�����u��蟝L�t<��	$�
:Χ���ӁBs4`-�,'�)�H�a彲�f,:o�
�J�À'V��rK9���0Y�2k���H^X�㟘�j�'bS]r��o��B�i;WR2�X�&P����!�YlVK'�,���37�T{��9R�I��h�D�:�4��D�g����Z�4%��S���e�`�IԷ�JoGOE {F�R��ͤ"�'��<���H[I�Z�b�/�����8���=�;FI8&9�q�'���M�irN[{�3��\=J K4�����p<�֩)��Q�t��;G����u*�Њ�aε��.8�̂�{��j�h��^� ��!"�'����% ������16��������h�&�x����\q J���cd��lVRt�������E-��(3V�qW��M��\ֶ1�|�?�6�ݻ�N��Wj�]a�g'��R@��Ũ݁�y���ꋯ^س��I���
�,���}���	�]���^ϒs��BG`g���X�|z� �'�ԇ����RW!����/���k�-�Q�"�F/����ŭ�h�ͩٱ _ ���-0����ߛ?cF�ʒ�Yc�i���Y�]�������<��؎�I��nFPpa���eF�kmЬ�)�_�_<;��(�C6��-k����//>ĳx�<��[��JlL��e;���|>������#>J����S�5��@,�A�v��9ǔ���Y����]_oق�md��z��Z ��!ʅ��!n6;R���@�����y��p�4s���m���}�^��؋��O����=���tHw��`J��N��Y2���S�� -�m@5Cv�M���s式��0k5��JqS,D�p���*���=��0��I��������يf�j�S`��O����fD�SVYI]��θ��88�Uh��G�]�={ml7�C�}�/Q�>��&?���p"�M�k�L��!J2�������V��	n����B:�:��4 �@��)���騨��q�K &�"
��@]���L�X��C`G���\E9{C12�pG�@$|�,�)[�s�eѧ&����Z'�0EP�ӣ_�+�'�3ƗL6_���4։ȯ�2�_�}���@ͳ�
���}��:W;���:ߋ����s���u�os�@�QD¦�\_��+/����
[��?43gc�¾_D��ѱ\���'7l��^���͑��Y}|�k��Qςt7%;1�g��H�JIx��cA��6
pL������������5��\A��XC�ɸb�Gǈ����:qϙy��U���CԜ�`�G9m���Ƈ��F�� ��Fq���?�!�	����>�kU4"��}��R�D�,�c�@�~��O�N��A�g#E�3�R��|�o<�['e%C�Z�t�2����'"/�����ONd�P	V ��>(���;fv`��Vak������&�|�uQ_01�K�)�n�2Z��em����--���1`�h� <~��T��>�Y�&������}VF5@��ٟ���yP��� W�g�@�r�ޚ�ef&��uD�8?��
��ܳq �7�LƮ� ^��ʪܯ����#)�4� 8�ʱ#÷r#���|�t�� jэ����%�di�r�b�D40>2��fʑ@���[�#|��{�ol. +�!7�NQ�L�������k{��$7�1Y��Ǝ(1'*
v(��X������YT�0����N�b�ǆ�X�؀^�5Q��W�R͚��>���+]�� ���g�`~�<��P�6[��!��&g?3������?/��?�v�Np�<�/tq���|�x2�A�Lsˀ-�ݹ2u�A�o�)վRW���
���1z�E�9�=�iWQLz��h�[=�[�~�T#��*���,�q�Y�5�뤆>+ּ�w���@]�}99�r��b<��E�p/U���Ә� L���������W_��/�z��F��}��9��;ޭ��{}{E�%�k��o�������O�\1j�CcV��$����8�?��}��?��޲�N6�?������T�E-�R ��Eʵboڗk},?����D��DU`�U�`�ۭ�6���=�0w��߻g���q��c���z�N?��� :�It�?�3n��'f����Vz3	M^�<K �줋|D0)�-��6�Za�M٠h/ߢ�*��������U������i���1+ssrJ&]o53�,��]����N,�`&Z{v�P��N����f�?b�zur� dB�K�NF�4�v�J��#d6��A�T �O�i�(N��Q�s� � @����)Y�����D��8*3I<AVV������)�U��fe[M",���~�$W�5�1P'�֬H��I�ş�_�{Q��L�T�Ϩ�a���a�Zf�ںvv	_\ئ橧���QȜ���G�TKay��;��^��6AVtO6SI}>��ET`� @��uIh�7J��	�,�g;{���+Fg " C��/��W/��m����@�UK> �j�1ב�j�E$�ȧ�],�}��D�-��ف jg�$ZW�!���Ѿ�T�u�m�|Mԇ'����8U�C���G*��{���B��FM��?�Uq�`w��繱���3<Ls��+��M'���k�W�j��A�u�ޅ<r��E�Cj~c:P7�y�ԛ��JX�� �Z���xZ���=���`AO�=��rH�xq��n�{};+�M#H1���4���MA�YQxr,�xFXe�Pl���̳;�.�A���8z�@�C��i����yO�#l�4ۈ���c�xؒ.8�s]S�n��;�2h�eͯ� eW:����J����9UIm4�r���vh��1R������w6x���ڞ� u����ª��6NR�V҇��H@���8g�B ���^�g�aJgw17f�:e/�U2�ڷ�����B��_��|����灬9��gS9����Ӱ#�Q�G��Q�!R�1k�T�d��,�_3V���m���]����9�;�kI`��|Nf�s�`�'����:I{��H=�JQΏ��B�+�;�3ׄ�PiHtgXD=!��`x�5Խ��m�b�ۙ#�?>�Ѽ3G�3���ψr�f��{q�j�/��Pn�S�{�Q���v�;��_㻿��~�_گ~�]������3�}���ݻ��@g��S� 7;����>�Q�{��o��o��~��O<��ǽ�P�]��w�����^�v�e-˿����/��{����l2�.�o�m~����] w[ U��h�K.?d�ȗ�z�w�����=��������^��gdh�?�U���˽���-l�����'�M���������e'� ����ڑ�H���ys����6�C��:ͣSی���*wN����j/7?��/�Cg}*u�f�T�]���K��%ʑ'�Y��Q&ĕO��T�����*5�&�̠�AW�Z���fQ��8ܗ{eTIG��
懄����s�%_��m��Ġ8w�����,��)�;;ݰ��� ��-����S� 2������Qbhe�Q��k� � M�������A��ԝ��)�Q�9M�F��xw}��"cg��61�"�c
6y��%���s|���\��w��a|Z��0��؀�YpGUs*GLo��M�y�YQi���n��!��F��}�z�7����W�+{��}�ŗ��/�.F�Ʈ�B��k=%�7�ow�F��duѰ|v�1�5�vfq�2�M�fw��Q���7*!yG�ttn0Pׂ�Աpo������b��C�#+]�1a�����e���	��ϣ���Tg���s[x�qG^�'|v�>�X�I�ca��ļ�prC�+�\��jRzXݲ� �]�À�L����7�.`��r��Y�p�Ej��2`t�<�7=I��,L��U-���{8)��XӪ�G.zd��Z�Թ8����,9��3�\i��z��o'U�k�����*�
-�*�$F�x�����T)�S�=8X��́�?�Qr7�s�z�!��� ��j��F�=dv]�=Ib�0|땢�נ���y���_ߍlr�������K������B��On ca�G��+�hd�Y͑���ꧠ���W��@�� a1�GNͼ�kС�J8�5�Tmu�%�o��Z�t�?u�4%J����F�N�g��޳���������xo	��9��U'7�ES�b]�)->��e�iy�K��s�/�.����p���M�|��ɰ�Z�4J�q�٣��|�Rؠ\��嘳�q�su����r��Mu{��e�.1M �������ŏW�g� ��9�B�|���Ξ���_\U�L��՛* ��渳۳�Q�/^�����������׿��}��]���#���D���� 7�H!���n\w��۵�|uk�X������2臛�X��B}fW�����H���s{�%�+p�]�E�"���\;4�g#�$��U��\��Ȼ/v��� �{,`��y�"�їױ���Q�t(�Q���K)�rS�8��F�������������������R���k��&L��);���y��=�r��GY� Y��im���h��� �?ꭦ�U�~���.N�:2)n�gS���ѹӄm���p�}/g�enn��2|
���KqZ��0E�g}�9ᬓ���w4'�h�\M2�Λ^����bJ��Z�W�f��^�J@��C@fAȢ�U �O~}���t���ū�#pI�o�gW�t6��oP�4qSx�^��r�z���7�7���dͮ�ΞP��%CzN̞1�}��u��GA� j'׫�k�*C��~Jr&[��U&` Csu���p���+f�Y�3����-�)iP$�:H�S�b��2��8���4����WT�����+��)�Jl��������
����Y�;lK����QO)���5Ѵ`�^�jT�DH�5���,�*�8y��q��I0�S��tjhy�긅ڞ�sa�$vNg�[�7L���5eYD�yݍ�z(s�)SoDt����d�~Ԗ���s`|R0��:�g����l�.�Y��EH�V���4[��5U`���i��gg�{��i��Z/��ȳ�!N>�y�ܼ���;WGj��'�k�KP�Lb��>�5��e���Q����ñ�}�D��5 �T��Sn$���)�1���<BS>��Nߥ�r����pP�p�ٖ��>�"J�.�yZƋ6%���:G�,�� #;�k.0Z��~��Č�Y��NPio�g�������kܠ��� ��}���`k��ZPԚ*�
c�NQ�����~x��޿��B�l�|⦁G��#5YdÖ�:�3�j���,.���\ȶ��g�?��g-nZ��h�gw�?�k�P:��?Ǯk�'�῀*yiO�O�?6,��O_c�Q��������9�-f�_���MRaƧ�R��\r@)?Wl��P�q�=�j�g~:M4��.w0�D�@(���%/j�� �e|��FG�i�3ٞ]?g-,l��4��n�>6q�R�9���v,�>�(�?h?&�����9ZG�ijwn�Į����~�����_��対-�GO��=v��×/&DՖ���T���%\o�vswm��K��Z1���&����v~��M�z��<��q�:��J1���ޡlH�RO"�{,J`R�YgkԌ�;:�������y= [���5�r��.�=�);���H���Wt��{���~��-{3�6�����D��� �M҇c x��w�u~p��j�&9�)׻�l�����ԾaOH�=p*�rF�|PXu�Ꝟ9z9D�L�~��Ʌ�06��[���*�ȝ|�ȈB͐48��A�`��b����+I�b�P��aG�n3(X*A
紧���H�meڐy�=�)82�x�Jɐ�S�f*p����ˊm�0��+�h�������r��Agl�ʎ˲R�~Ԩ(�&�D�:��m �47P+�~�q,��4�����J���g���Ы�<�sW?��L7)�~��*�K�劌���Y%����a
�)u:yr$l�Q�3�������M�1��3_����,����5�����SWdH�Q��ɒ����<�k*-{��օ�۫���W�7�?��~cϟ�����n�vD���֮�B)�WD�N�¢����	��Pj�E�`���1^��wzO^�)�"��jo쫁�1*�.ì������P�R�N��{ӕt�sr�\*H����72\� .�Q���0�-�Z���O��4/�������y��"���XJU��~�?�4�/1�5�G�)G8��>�����E{��q	$�},9�i�x�����z�����ҩ�?tiQ�Z�.a����"����;��z�t������g�9��٩�M�N�&�Q�-��~1b�+#���i���`�g�+���9V�`Y���$��\��K:r,<�$�5hl�x鿋�K<��#�7���i�x �;��=�i�ӎ���UW�:<����aO۹�?�a�=?�?��2ٛ7o�O��޾}W�w�ė7jv
�?))^��&���Q�>�,������j���q����S�.`_u�SĵDHⳀV4���Y8�m�
����cA�3@�p�ϩwɝ�O������}���������{a��g��.Բ�";�c��˄H��v$8�)Ue3��PrJ��u� R��b�n�{��M�ly���n��2X�c����ŏr���8��E9�3��#{��/Zb�=i����+u�}nv������}����:۫��ށB׳F�Y`�+�ٜ�`(��=������1��A��=��7��I��,?U~�}�t��SpAd�M����=(4C��%:��v���R��t�7���eXSs*ߣ��>G/�� ��ڲ�vMfњ���m�^1<�j�������h?��}m��6>�o�\�IGfi�Ԍ��	��,��}*�(�n�}� ��L��	Dv�أ��\;gG�'ʮv�(��:��A��U�;�e ���My��5� f�Y��8���N��E*݂f�{
�\���B�MU��w<��mpL��Z3�x����tT0�tz<'����,���&�۵�X;�kY�}^�Q�p��@g$�
�]�deC�
�7q���1����ut`V ��+?&�G���+�LI���.:�=o�u�]T�&
~�#+g	��s��z�a�^qK?|z�K�]m�|��ө�!�6�� �	�Oj���=@�=�T��e�6�])�^�����n�u���P[���aoU�⠆���хZ���o鬱�?�����X}����)-6��������ذo��'Fz
Tl�CE�)_8Xw�W�W��ۿ���~�`m����a�ō,��ꛎ��p���t�f���o�B��$���XN5��4�KN>�ը/wdh�N�:3AÈ�j���k����m�iB<� ������חltpI�F�=n���+�kI�l������j&�r�燎	�R�Y���Q�1y�FY��÷؜�㐵��rR/N�ccOmX�_�T���6mbM�|<�� ;U�>��e�����:�E�ʂ��;��S�T�+=��\�>��9؎�Wjns�#��$�э=�ץ>���ȝ�g���;`�J^��N;��&E��?��#��s�yW9ҳXF���P���r�3L���7��������^+�56@���A���P$ן���t�Ĉ$688���7�cqT˱^� ?�xAA+������#�*�v��3}��쒅xIn�9>�K'�Ί��ESu����g�P-�g��
����9�^yu�Î�*��g�k�Tt@�5J|Z_��{;�s�����z�3�^������ų�s���y ����������
	������������Q�
|Ꞝ�}������_�},`Wʱ�{V:n,�*h&�|�[��:�r@� ^΁��599�8��)-$� � ��m~L�b��I��U�����Rr���<� ��2�5�^C�����ݿ?С�}��3��Jc{S��:�<<��	$uk�^[,Q8�ϓ�"{0q@�CHhg��A-��iO{����nP6�~FX��V����p��C�2�T�l=��� n��A�_Pqs�Z���F��7g����ܔ�}��W��~�K�����˿���֮�;܎S���?6�3l�g
� <@�2X3m튼�Dyv���w�^l]��;�dP����H%GS4#E6lʢvC��I�=d�fG�uN�D�#�R���wf�G#��\Y�8kKs3k�� �V�"�8�〦�Z<����"�E��2� ��U��S�����pĳ���y؟)�0n7W[{p@9��R����Px0C&���ve�(�v�8�DߪG�m���� �#�����P;Lv�tK�T)�0�N�y�݊A��U���A���� ���nE?h��$�&��µC��a��ź�\��	J娭����5_�8�_��bq���D`<#dn���9�e�.���n-�_=�dy륰�U���$w�,�����>-_f�o'7�)О&d�o�BD����'&z���EY���_�Ͽ��������|CІѠ����={I̳jEع|�fʽ��Y)�P�g4��������_�Db犍����M�.���)VGƛA��M�+��M&��v�y�0\��ю4lݜr���6�n���Z�8����`��3�nN�S�^��n��Kea��Ũ}�s$Qs�4*��E�ڋ�:_��,>N��}M��d�6�m���/"�u48K�U��4�y*-�ϔ�tA�	,�֨YHrD�� �u�!֟�EZN������&	�L��c��x~`:׺���C�	jy\�3�͟u�WW����N��3ߝ<u����>�����.k��%�V餂|�ug�H h;M
_<#S�t�������桘�t �����ll֐`��5���r�'�߿�����8.�x#Bd�A�@v�.�u�|tA�l�p����r�������ީs�c ���gq���� �ۉ�O?�ݟ~-6s���tN��
e�s.�~=9�]8�^�.�ڌH�����.��1-�*��k`����?���3Q[��%�<�W}�n6��D�lCP��u�s@�B7��e�Zߪ�6"-����<�ӟ�
�U�-�� ~�/������R��c�`c��[\���&ߗbOM��Z;���E���6���ph���ɥ��*[���4hn������WϋSv�u�����<<�������f����Ŏ�H˄s��t$w�\=+�d'�8�e����4G�	�����{>�G�=P;��#d؋�:�e� �ph]swsk����#�r��DӃ�vd�G~�W����Y��[
xlx�1�Gg�ף�EqJo!ұ�f�e���C�� Ϡ������,�FM�q��#З�;�$�qm2���@��;�5bD��(�[ b�Ty����K#�ۡ�)����Dg/2�T�Y`�Z"�m'�Ҕ=f?V�Kd�Ge,��HM��{i/�Xqo���A�{Z�f�Z=�����#p�(��s�q@�H�cyN(�Y��ݲgЗF3�|�f�r�Ӿ��NB(ndPCX��=������^��`
mo:��k�K�IM��L0��L|�i;��M�(��OaL�|���uhtܫ����T�ϵ�}�k}���ҹR/�27����T0���}JN�n���[��h^��27uG�t�i�m�Y��#��>g9�9k����u��)�J��ZFÈ��3R�X����!� ���9�e���8��Pb��t�;6��b���vg_������������b��M��� -����7�����R��x<�{N�s�Q���y�:�QN=o����	��B�Y�i�dB	Y(�Q���V���]e>Q�;;�Ȯ���������a�+`�z�І���}�o۴j�ӬJ�6�am�Ù��T�X�Ԫ��[��f}E\�R�΢��������f�ߗ�u�\?��8ܽ���z�D#��1�������6g��϶��~�S�����8H^LN�`���XK=����:VE4rsZd��p�>�y�>sPV��>d�S8cU���@���[���B���W�ר��f2{��:�4'����
jDa�*���8~���={�L@n�����9.��FC�l��˖�x�Xcp,Nϡ8�FM�ɲ�L0
�!~�32x�����gc{�q����Q��ֿ�f��`O���b��湯˚.����v��[#�]o���-i$!0�sYKH�PמG�j����h����jT��[�%�r̺��n�'�����sI�<��4��~P����uK:h:K���Y�A�(��x���v5���|U�dq=�︖Jwco�e���HjN��j�Z����}0΋�;�郱��q��Vy���cq��]��U��I#�M�}q-Ѥ=�~���o]���
~![��G[��un����Q͕=wV�~�Z�1{��M��%F�5�J{�G���Q�Y|>%R����%���ΝZ�p��{�m�Z������u7sq.@�����oP����Dq�Es2���h?>������Ï�?|i����b>��U�������{�����l���޽?��;��6R�+ ���D I���%d�T�2�	�ծ8��t(!��H;�/l#�ԟ(X���<1k����^�xn/_�����IǹDͬ�Z�4G�5\û�T|�����m�V;�vd ���<��no��w�}]���n��\��~~,�sπ���\`�1�jE�;��GS�'�zdf<���`-���^+#NQ\w$��i����=��X�k��y}�q�<x�\��N�z�i�`���!�M&q��r��Je*�c�F����!��&�&�A�]kx��bl�%F��,��af�cv��lV���wa�n��Q��N�Ε�.�{qJ̞���@�ޘY������V����lT�5�&;P����d�2�q6ܓ� �ʞ V�:�a�L[�:֫��T�]���^��؞d��֫�w��,�A�5i��(�+�+2���=	e�s�ư�?�K�5j�X���p���ZB+��EC�.(׉�������W��&C�;����=]?��@�r����E�}�V����0������#g����l��pĊt������~e���~��R2t5�ب�Pn�I��r���3%Lon`<Vu��ҿ�أb�1Ϭ�b��N���{fdms��p�	�S{�G���
�����Gqe�fkNC�e�#`(���@α��[V�fC���b��8rs����K�o-py���z����l���]��-�[s�d-��dm�}��+s��m-�^\^`S�s-��Ź�����6��k�P&PW�y�ہ�;}�!�!Q�E�X�i�� E�g��F�ђ*��On��<׸u��ǦD=F�͡o��:y��K�~�B��K*�EP��+�1聧�$9�Q���T�`ԑ�C=���%G���E-D�T��"s?������W���_�����ߗc<����FO�ٗ �VRy�\f{Z�g[Ly3){��8�F�)dv�Y�C]��^%CXM�!+"S3�g�=���gܨd��L���8V��|�}� �oW���boE��P.��s`��K���E����J|d�+������
� �����j-Ր�XƇ*H�li	j�iqV}oiw��a���}Y]~|�b`89�0k�.��倉^A��P1�(/Us�.��� jE�ͮʧᴸ@����{�L�ʜ'�������t�������ü�9{���3L�ď4Q�(��{�{�nm�F�E�g��pMX�p�@1;H膣�T#�M���������`?�~m������?�������b����06�
 c��N?�IPO�^V��E��rNԦX�᝚*[}p�S뚍Ag]�aOe��a �[�P џ~��^ ��T��qO��kF�
dT������x(~U\�rG}Ty�+63^������{ُ�������/M����_���ڷ95d�Q�=e�}a'D�2w�5���GN�HT��\��hs�%>=s���r�X(��!��p>4���v�T:��䊌S��vP�]�]�\��M��Ϲ���|ʤH�q����_����ho�3 \�wX�	$�]��͝7�U�h�=�>��ḁ�7L��F�I&;B��I�!*qﶶO
��@^�5�~`�NlX�L����xG}��j�S(4C�y���*�zw�'Քk�3�L7k��Y�� �5`�@�y@���.0\�=ԛ-3[�����@��p���b�M7�y�V)�19K�:�m�0�=b:E�@�X5�s|������ЎeI�=2K@]�4�I��pf�{���bgώ����|�j��f��5�x����n���ͱ,]�Os"����h�Y�υ�	�8�#�~Hm���ݷ��/�����/X��/~��ѡ�!�����x�vwd�k����o��V|3N�5��Y���CD�2,�}�g�{�r�i�JQ#S܉�|;AY�0Ɔ�NPKD��7�'Z�R驃��[�n��0���v�ӯ�d��Ks�~O��=�<��������B!Y����,��p',���p9y�������Ǐ��x���'�|0���W{D��N`r`4��`��+N�)����x�%�g�qy&��Rc��2��)I5|थ��R�~i��:�1hs�k�(~���z�Nhaf�<�S(ޒ��s�ڣz� ����������2��C��AE�G*@͌T�vGQ#���U �lE�T_��#��݈��Z/4ݞ_*+Ң��,%<.قld�@K� ��"��8�ǲiI�L��Z��BK�5z�����n��^X��߻�'@{F������;�;�S�}��2��'w���J���9x�3���U�{����=ٲ7=��d�2-�5�^�-J7Tm��������gœ�]z�̂r6����� q��d5Gɝ���}ft�"�P���0�[D�v�w���~:��oR�r���|�9k�ȓ�t�z~�9f\�`{�̬-����(�?�7�M����b9��?>�iFV��KvǙ���XU���-��G�u���F<��Wvyq%��S�0G�;귿�����������i��������:u=�v�u�u~�G�F��|GPl�
W��F�����ݩa�}�2�� �V.��ޣ�!�oo����}�|mϯ.iS��nmW�����-P��V[��p�|���Hl迡�t9(����T�{vuU�������*��/^�t�V�AﲖME��A�qR�N�nZ�s�C�������BM��蔭$�� �j�1l:�1�pVu���0��6J�ŎT�_#p�Q����>��'��0.�;x,��f� J((a����"ˊZ��!Ӄ��g`	��������AcO�=	�l�'K�i��;���Aj��g�Qs7����Z��zO�R��MJlHR�u� 3,�Y���5Pwp�<�=��� k����ؔ��g�mt�g�A6����x��7U��\�P��
ۋ��Z�t٪P��ߐ�
���s;��YnXS�;x>�<�`M���i?p_>w�j7�3��~d�T�(R�2\Cv}���16�ΪY<�D9��$,��bGL\,d�޼~S97G��1J����������7��?��{����~x��YJ�n�Ӽ8�d�,BΓԔ���.��Nj���s��F�0Kb:�1#F�u���u�9	���9A�n`mWw�����R�9�ZR�x6����}��(�� Y�]vsf��'�Ki�p�\�x-���gw�yk��N|�t���qz8�5��s>��ù�zz��7]"E�o��������+%?������g@����΍lh��+�2��=^�g��գïK��[<ww^_>���v��>�-����?�xn��GO*p��{d���� ����D'*K������asv����CAh����A���n�k5�d��,'��ރ�s�ۓz'!��ƙ�"/��R��,֪���i�*�����A�ޅ6,��ʉS��j�z�]�-c�Ͻ�m=���ٞR<�ԭ� ܥ=�p�O��s\s"��b%/t��d��Pmer�`��4��v��Y65�S�,�%��O2ehJ�u��M�� �͒��c'��e�lyϣ@�= U���A-/�5��	��@a�χV�%@�>�yj��ȭd��}�� Z~GEr����ᱽ_�j��-N=0 E�+p0�&��	�[Z��wms$@)A^�.�h$�gp�t�ՁLއ�Ƞ9�ϔ�5A�'��H�D��N�����1|���}�ͷ������7o����z�3���[���������O�������S��
R. :F֓��f�Ci/����W��sR�:fV�DRR@�g).����D��сiPt|3Ϲ�&f�o*���既2�7#)���E���8�gk���îY�o�P������>~��Od��X��KG�,�s��vsAJ 5�0���D\kfq�s�m
�ݮ�<d�+��<�z�眠E 8׳2E��=���aU���3+��(MݙY=�,ԣ�keoH+^�;xb@x���CĂ`ƜBVǉL��@���A�Y�z� �~vG�m�sƦ��f;G�_Gϖ�CA�,�u�:k�ɚ��:�Ƒ�T 0�oJ��٪�[���t:6�N
~0��c���	�%D}�י]D����S���j3����Ǣ�������轵��^;�y��  �+f��`�J��LV� �!8���j<��r��?��]���\ySh*
 �w:ߤ�Y�ۇ��jT����{���/�,;�m��u���}:8ӹe�b�I.&0�&8��]�d)x���� �{W��W����[���~o����l���o짟>r� P�x��޼���|i/_��/��Ҿ���a�r�(�̔>�oCç�*���z����eI4"�~�	{�U�l��o��� 	}���"���rD꺿�9P��-��z���9�֜w���#�� t��Q@��QV\�r :���u٪�8��k=ɀ����������l�����J����OˉO��<�Π��X��Ǎ%M97`C�Y�)��H�1'�s�䶾����+�ZG��ܤ�D72\�P�1�Z��q�w�C�GT��;9�O�_7b�Y�k0?1#k���� 	�ՠ���Q�f�ExἠG�|���0����vR&�XlV[Q��6�{l�T�q������S-����v{w�:[mE�IɃB����x@���5:�����,x��Q��h��Ï�|iT�_Ԩa��i�%/��E��|�K9��3����lHv�Hm�C����,�Pd�-I~�1�-���b!�����9@D���j�1�E7�9�Q���|���"�����]���"�*~_�w"A=�;�l��y�7�"X1�bv�� �s*�)�l<�t��j�{̒	gm�
���&Ϡ�܌g�: T��!_9h�+��;����`��NS�`�I
 �I?~�c�9<���r_[���a%�ϥ4��c>���^_����G�'#S������B;�qkЄ_�_��/�����W���|��A�u�����������?3h����U���;�o�#� )��`sh�y�X���1^����8�j�	bX����Sh������G�=b|�Fo
/���?3"����?2�fW@<�z�3Ȼ۽�և�O�w�P>�Ķ���,�lǙ k.����3q�z�̱E���j���p/%����H?�);�}J}���8x�G���VRP��U�]%�<H�O C��|PdA��wJ�f��ޡ�H�G3��� |��~���w��Q�~�	�����d���J��X�������`����{�g�V���� �:Nꛉ9�f�E��꽠W��1�^��͜)�~d�I�_�rj�+ PC`���z��O�ㆾ`���̮>lʴq���źt?��S(K{p.�|nh5��d�b��"j��N�#��4�֐@���;��`�$[J��:�� zu��_W�qR�YEO�h��cA+�/��+"�m3es���B�9M��5Vt�z��m��Ee��E����9�!��������?��~U����Q��n7�4D�/_�X��W��w�1����+{�}|�HcQ�\�%@Į#�4v8�'�k�	�����E[�(���5i�p6s_�-p�Y���EO��7�8i������O�u�����O��SЋ�����W�"���8����8��G[�O���{y�N�� �dOx�#uH�ߣv�7���.� Yy�Oƣ�u�.������K��<	XL�`!�ߦR^��r��ζ-����O�i��i�{��C���Ȝ�CZlK���
�)K�"�uB9}�.�P�lŴp>���8k�ϪI@���ng��}�<��1��TX>��L�{�)�O�˵�*�L8��"������o~k����?Vg���k��,d^��=�ڲ�Lj�l�����X��:�1���J�C��c��h �[4*4��`��Y�R��CY,mZ��&��-xB`SwѾ0�o�}���b��G9q}̆8T`=�\�>?(��'��x��ɜ�a�n�Ӊ"Ty�ނ�v�Ǯ�ӡ�E��ھX��Ѳ�Tˌ�!�6*n�d͚��"��R�Y��bL"���f�81Ҳ;��ذ�V�=�< ��W�x�G���.�c��]Wv�in}�Hz �N��Ә_���\bH|�z�PO��jq�S{�����^� i�$���B6��zp�8��!�qcW�^�_~]}�o�����1ϊ���d���������o�S�+��3�*r
GÕך�9m��kI�	�.?aT����ʤ����X��=/�y�3Z�����@'��C6�@W C(d��B�wPAEd�/I b�:gp��N�d?���j����]����|��+�n�N�XJ��lY�L<�	�W�@�&�)����h�i�f?&�Ĩ[F���I��P�jtv{44�ܮ8��:F�á�dA'K^p0��'eU4Ι�OR�Z����{��"�k�Ǳ3�S��������.�DVs��"��X��-^�ٕh�B2�թy��(#4�ܲ>���wbT5��A�j�[A���L���xh�,���HB� � 3e^l�c"��cqtkv�����*�g�G���d�@S؁�q��-S8�7�cFr=.���I���-��/�A#���GL��s��� Y�k����7���ϡ8��B�@�����L2z� �v;��������P�����������?���������?�EQ�y%ŗzc�7��T8Q�ϯ�!��n�1�P�VPm�N>=�D�Ơ��F�fY�"�}7�J���U|���q4���-���z�4/��K�{�9ui���/'�X������=UL޿���㖗��<=�i��)7�!V� vj�G(@����dO���7寓���r�����=6�jAQK��i��`�w�|v@�s�y��k�H>K��������G���9�m޵�D��cĕtC�z�e�D���G������;�c3@a�q��b*�9�@X�xWB�5d~A8hƉ�y�k�ڬٓ�k�D�c�m���g�������'��ǟ�ڰU}_'Mp"k=i, R5�X�I8��\B�;�����a0
r���]��-C_}���u�G68�v�OLq��i�|�n$l$P%g��E'���`��&��B��y��Z��Y�\\���ؐ�����F<�����@V�������y`�_vm�J[�f��=q-���`Ѭ�;h���*�v��X�:���{��{�l`|�M�+����g�/����NM8+p0�,�c'@;�Ջ��F
/���G��9�)�4H�1�җ�,�9>��o�Jn�ʀh���o��ਨ4�,��2�
���ƽ�2v}sm�޿���߲_3��S���8�+[��m�=�	��֢ k�c�[�T���.�[��O�^��'ù��)tys�_��o�ψ&	0�5W��Co�d	���'�pP����D
��O���o��^�z�f���������{eG��YdPrV�R�!%���򍚸�(8��YdZb.�-�z)��'�9vB�/E�R�=T��(�V��JI�q�+�̍ �%�/�$qsV)�B8W�}mZ���Ƴ�s�yH�{&�͠��Mj��J�l�u�} )�}��mAt��a�Z�~ä�Y���������ŶDĀ*w9�M��\���e	�9С/շ�"�d�x{#������)�s[�C�^dGs؂��9�@/�߿X��`m���\3���	,{�� @翡Ĳ��Bا�����YS�K_���s�m�'�٣P�,����Р�G�϶�f�J�!�х��{����?������_������Gn*RT��ё&Ɏd�X\9��n��sN��C�'��z\�����}�pb�w�6��؊��d��,j�l��ɚL�����-������>�� ���Na�_C���s�C��'~A̅��ʏ�����R���gѣLV�^K� ]ԼwƊ5�������,�,?F�� mh�o�&C�G�+�/��Z�R�՝O�,����F��e-� ��[�!/.���'k���p�:�U�LݤIᣚ�&�^J�����8����sXJ7srs�����
���g�Cl�$�A	ޕKDg�hE�Y��3#�(�m��ٲ�=%�,�#�H>S��������B��� |��g�LO�$���ѵ�O�����,��S6-s��/��z�Ρ�O���5;��Px�ާ�A�s�^��j_#]i/^�k��xM��u8�(r�Z��+���{lN	!�24��T�����s�~~�Nt&(��0�-�=A��u-�v1Y=�+KУ]P��5�BC��c�j�H�ݣYS�
{%���
�g�lJ<���'�O *��|:�߃�ce��ꖾ~�"~����Y�q��=�d'�$|,��o`�m�yI��ى"Ų2ǁ��sL؈*ջ�L�����Wo���w������ގ�vu��=3�3ORqی�<��7�Sf�x�
i��zIY��+d�9�<<r�&��)hM]���Ą+��d-�1��@l�-&1��c�x���IA$=� �suEa>������,������'����A��_�\�4���ן� �p��}���@�~X��D��n�'�u���rH��z�Kƽ�`	ssw�����e<01�����o�S�̒�R{���B�6�m)7fe�6����E[��Ū��=���Z� �T��1WP���k:8�"�Adyx����q�A������&�p�h:�����}+ '�-�>�p���(3�L-����0K0*�&E%ĕ����pr{����6�"A1nx>mx�Z[���۩�4����7���m����;uIƱ�Į�� u���*�s�J]Wu��'��Wk;�s]����o+�����׿��~z�	�����ꌨ�i������y�,�DD)rwHhx��㉀[�����H̶�f���2�Z�������2��n�\jW4yc�;�j��g�#t��R<��b�h�6]���>� Z n��8�}Qyy
f��E�Sj�$-���\s\g�B�ܹ5g�<|q,� 
�7���҃q/''YC8�= 螪,j��N��gW�����|wϓ��{%�Y���A�1��r���&@0^�ya��_������y��dI�A��6��>��k>.�jC� �Q���r�E���Yp��Z�Y�.��h���m�)��^gT�d)-AZv,��2WX��0>�l�4����r���mP�rYs��i2�c8�YR،b�$uNo&�4�Y�^�c(�6mNhR�S���@�.�0�G���O��T<{��L������8FDʅG�#=�%��:��x�rR�q����VV@��v�ۼ�O���,Ns.��jΚ~��o����'M[	-06�7`���'���<� �1�4�Z���ee��Q�Zi��i�{�N%�-"#|�Y�Ĝ��Ԕ���թxf��� ?��n�Oʿ�.��p^�DԤ��^�g�TS�{�c3{Ѓ@�����V�eX�U<C��6*�AB�;�A�R�5�F�\���O���?ڧ�C�Ad^V^��؛�,��b�~2���Y������=c�vv,ƽ�i��\tҳ��Oj�Z�
NO.O����]��+KnQ6u�L���=К��Z�Bs
�2�Ϟ?c���>]ӯ�؄�"��C ��� ���6�����[[$*AO���M^�;���B7�Y|s9:(1����Գm=
`!S��aD�(�\�c����=���1[��I��F�	�?z7�p�=�H�}��WH7��4��S�;�Z��>[�~��u���>����= ��9�a_9��XIY�� �T֢,>c�~)��)���qmw +�A�~EYhh�T�F:.2Yc�*ٞ��1���`�x�kqľ���!�� ˴�QIr��V-(�ZJ�%}������6	���c�S�<gO��λU�؁�R�)l�a�>WV͙z����#����k�ư�v�,#��6S�|ń#�����W��W_٫ׯ��[�
�pt�?2"�c�_�z-5���+usd��c �P��Oʤ�|cLRw�y�}�Js\��@��^����-3�oƗz���f����$/�tjNk�P�P?(�4��{�O�����Sa�b/��� ������Z�t����|5/a��`���n,��	 �hrl�m������	����ZKB�+����C�z�{%3�~���Ł��4�~x�ݽ<k���Th8E]F��I+˓���,��;�5*�%�{b޸��s<�Lj������sI��Y�a;��5o�Kl&���wzoF�ˤ���/*g��r�33���b�Q�I<6�;��,�u~�f���FR�2��u�"\T�}��fmԖ��w��!-Ur�!�aA��ܞ�Ơȁ�C�4�g�[4�a����5 #��X��1Gc�j,�k����z�X������S$�DK�����ԃ���b���9��m�$SY� ��ù]o#�<A<��e���50���[`�T��N������ ��������@̇��35�����ˮ��6�(�Ŝ!����$0���L�T�i���^�Ee}���5{T<sJf|Mu5��B�E�#�B�r_?\Ʈ���(�A��÷��Y|���f�x�F�m�-��`gf�9_i�V��Ӱq)v�|�!L0+�w#�뺂��~�����~uEQ-�t@�Sdu >�E�xP�S]��ʈ�v�ȴڬA5Z|FGe��F�g�>�@HЇ�G���v��$x���6@�+� 3l<�\F�it�M�b��Z'X��(�H����*Ⱥ��vV*�Z��ن����j'�������F��zk��҂J��,�2��;y�]Q�դ��0���Vi�6O�</sX����`�]�1��#OG�}�)�P\2>��A˃@��M�la{��xf�|�*A!���6n-��Q ?��G��4{	��I���l�dld��j_Kc�$j�r�Y�*�u��4(��^lVZ�&y�/�:ͳ�Q�Īu� �1ӄy��@����� %aSi{Fe*���8���x	�|�=-�Ɣ��#���"�M�ɟ��K�:���4��̜�h�ٯQ�`�ܘ,�l�=������/��ӥ�ߵ�x����eۣz�9t��<�����:�5/���Ď�PD�.��꙽��;��o����6��Z0/6�Y������_ط�a���{x�����V��Ym���cS�Ml��(��J�#M�b�uX5�����0�gc�ގu��[���~f�1Le��Y��!Db,"��%�0����5/Ԏ�9�ȃ޵����v�]G�Q�}8��e���� WQ��'�O��5���+�'M!Qn��6�"���;���,��֜:�u���x���.��3�i��������52^iu��Ꮱ�U82�z�]v�2Gx�w�o?:�#�Ə��D��|i�g?t���{�A�@��1Kη�{�-|�Ҁ�2ߚ����?|t�y[��wdO���6	���=հ{ks�����2j]�լ��E�3���Zڸ���b�4�*�P�I�`w�s�����p�7�7��n��jc���C���NѺ����ػ���͍��}��K9�@��ʮ�%{�|�DuG�]]\��j��6�x��#��gWԢ�ϭ���7k�[9�Rd>s��n9T�~~1b՚�;�xZ�Ue�w�K&j��Q��ƥ^/���OG��d��/i�j��=�TLd���=	[�͊�b���׆c� ͩ��LMQ -qnO���e|�Ã&�gt|�X
-)s�䙒b�ƕ
�o�j�y�"R[�a��5�&� �n�o�n��9��ug��a�ˤ5k�2'�Lē'5��z��U/A	Q������<h�9�u�������s
.���jT?J�S��6�m@��Y���n3�E33�,��Y��o�O�ѹ�j��P@�s��;��X+�*�͞16��Η�U]�h���"�a��-Fr���[���:�Ú�gk8C������uC����z�&zҼ}vu~YA����ӧ:Ǫf���zuG�r�\@��.l����衔�/�09H�$��|�����>�N��Ug՗y�:�g/�U=������{�T���6���Z�d��XC�u��܇ݾ:�����?W'Ab�t�~K46�~O�Tm��g�_¾ʚ��=�6���}��	>�=�cI�?�v���!���*��{�·�+�	gљ�$9��f��//���3;ߘ]l�s��s�!�^l��D�Q�@�Pi������:��c4D=;�׹*���z��jo.���&8�ޖ��E�!`�N�\9�KUv<��͹�_�؇���m��@*�P��P�ͷ�XR�<c��i{ɹ	��q'e��z}�����L�W��2�.\�z��,���Ʉc���LBؤ���|A&�쌵ih�E���;jA�F����z�%[�����·�J�v�S�u�N;��a����8]x u�bpd��`t@����^���-׋�y0>��>�u=��'�;��#��z]�X���y��[f!���P��N�1x}�mb#dX�O�?�k�Ӿ\>N�����:���^�+k��x�����PJt}g��Wl�=y��F�F5L�9��9�����X<���@�W�%��հ&3`{&!�#���-�#��E��ﭠ��7+~#1�eĎ.�<9a�1u���>B���#����6�&
A�,� �V��z/^<����L��R'��/��ۿ��N�;���G{��-(�*���ƾ��+;�)]l./�����- �
�U��Ŕe�I�n�4O�"�����m�e���hd�h2��;�'��嵧$!4�f�Թ}B���tQY9�ÒMq�.�>����O7�8e��š�V3Ϣ�W����c��-�G�_��XP�J(�D\�=�V��O��,�?��"��\���~����Ex<�/- ��Ч�{�Ǔt������䑥Țv����4�h�5_�o�1�d�u9���|j$%OMʘ�f-Ӛ|>��K����%{���y�蟇���"z��&���#�t�Ge� ֫hX�h�9p\��R�°��~�;E�@^'���V!"��C9-"^�|ɚo���N��E!���
�`���ƚ{/db��k�Ȓ ���PL@�8(�4��B&�T��^9�1���� ��	jIH����ZK[���	T����]� ��q-��ޓ��l��8��!@XJ-+7�D7�;T�@�P&�|��lT��^-j���&s�M�n�5�ò�|k���/��zj�?�gz��2>c�N?��k�O��$�&�s�bs?�ڶ�3�F��9�XwB9��R���p)�@�Lr۔1�<)1�|q<�m=���9A�1}�Y�\�X��� �5D�.@7'�v�%�n
�;.�e�E�ϙ��S����u]C{4�c�D�\Q��9�?�[�{�{��F�Ua�QׁqKu|����D �)5��娝:�,�o��3�\�|�¾x����G���ޖ~qE�[},�B�8�ݑ{�ٶ��/��rEJ�BQ5���L��``�U�����x����VN�M\qm�ф8F����[G�$:�瞊��ǶNTb-��&�v���=; ^sn���W��˫K��ߗ��;�X�T���D?���mNۂ���ǵ~ k��	�:���W�AW %`�s���\?C�£Zu��WQ��BM��zy]�3t��s�_������gy�)����5s��x����ڷ�!��w�@�1��j�Ϋ��IY/� ������ђ�v�͚����=�Ic��&)?���K۟��qQ��j�u�X[k��A� �dW�\q��	��1�a�������0+��}
�{[Ac����*Z�����^{��7����n��v %j��k���Ω�1�\ l�E�s�]����h���y��c2���Tn����v�DA����5�<WWϘD?843��|\������R(-*���ѧ�Ȗ7+_�~��]�Ȕ��es�[S���s�%5�(=�I��xY�R�b)�Y�&����B�L�1�����g:_�����;�����lD�����#���n(D�#�I�I[;v>�R�[��H�%R�z�JI8���k��,w�#�#Y�G>��翴�'y�m�˃�4���g�V��w
��Ɂ��%�i�
g"J�t�S*��yS�����:�^�B��!��X�nEt!^Ծ��4?O���ε\��ٹ\����^V�ܣ����X	����I�O50ߕ��ƫ%��Љ�9����nK|$����&<�� \�@�zZ=x��";�\��k7��N/��.�6K�c-����'���2g��N�m�5�;�$�"��=?��C�Q��l�yP�~V�3ի�-�����^Tg���7��c}���D.���2-��XȻf!1Z7L��uҋ�����ʕ��m���&����G��% 4�����7Q��B�n�s:#l7k������u����:�9��faX�Ȫ�d`�I|�� ��F�?N�6��dZ�퇃�#���횛3k�`A�bl�Y�1F�N�'?�d�!=Z���u4�O�"� J�Q��ݓ#S�A¢�A�@g�6w�?լ ø��C6+Mr�P�2N+�5bK.\@Z+3��9������+<-��Џ�������!�5�$U4��(�p�<�^�<X8bp4�3v�5�C٬����Qv*���^�T�;;��#��?
l�8�Ԓ�κYy]���p��[  <��(#�1��G  A�]���.�9{�0C�~m�=G���K����}i5J�_{�����HY��֘��N����{ `M�_]����/쯾��*0��*߇w������S=h�u�볫ޓ�|��}�Ӱm�!( ¡��:IPp���v��̴�V�k�^�Q��H�$��h�l��]������.1�	�?��\{]����ٳ՗{a���?f�q����#���9)U����'���=� ێ6�}9[#�U�BZ�'�n����/��~�y��Ce@ڛz�[ �-�֬]��?�k
��<{.3յ1p���(�[&n�a_�yroH*�g& ��B�م��5�	�E�&%�5�Q���D�.�m$�|�^��w�g[=��^L� *$����\��ڻ�G�(ʚ@���Y��G��ge�+,�Y�C̵���Pǖ챣�؇1P��޹���{B�h���Q�&�t>a�Y�p?�����<�9p�c�,i�ؚ@5W���=cѪ YY��]r�v���9�*�[���m;k��5{��O�bnL\/��&�ET�����Il�dw���B�^m�F�b�9���=Kb#��e.I�+
w�4��wL7�ݪ�r���7~a��?������?����Pӷ\��޾c�@�if,����D&�w�P��ܜ��Z�p��b���ڨ��V���
'5����Qk�����q=vZ���K�#k��G>A��[�u�x�J�Y�q� .��F����V����p�&��+�=r�mq�,NG�-W�	�T��H��d���UD���, &����!	��v>?�T:��ey���#��/`�T��<�T��HLj���,�	�Z�I�^��\"��_sԞ� T��Ɯ-.��l�� ��UJ:y=���4c�L;�����k�[�͌�g���ѻ�K��s�U\�z(W����F��w��_өB:"X{v���n�a�pqyŦ�ϟ?�#q<������jI�_��	 ����9&W߉:I|�F�z|f %b��D�,j=��82��TR���`�Nq�Z-e5��>y���������������/CУ;f<�uE��A%�(A��QA_�!%�{�8�Z�I*6k���T3h=�ϒl{y ؃jcݠf���p�Q�!.����oKx����t�9N��v�e��_��sh
G9�iul�� �EXV�Lg,�T������	:.�x�Z��<��������gs$��E�)�l�� dp*]�c�S��>GP��{��Q^	��GN�.��V���w��5@�@�R�ke?����͸X[���\s���j;�ď���,J�y"　��q:DQ��>@�D[K�;F�Aɼ������5���� �9�=i�,�zS*5ޣ�����D�ĺ@����s���|m���g����`�����~�/�����h���
$c=��@�8����ǚι� y�>~�ۛ��|�l����R�AwM��m�7�ɔ��oH�h���3۲9K���>��'��������5����7�_�T��YUO��!肌��V�1gmi�QKmh>
	����,��Cf�8(P�{C�j��S^���i��OR<� �1!/�?��֨+�H����E�Ѽș��}�Nަd���lRb�C ]+*dy�j7��E싦���s 8l�?��:ϴ!�y<�7�ذ�(%H�H)�-f�$�������OI�I�G0A��:2W��x�ss��LH~ͼn��������c}���{d
����V�u�efG�6�D��q�I�E0c���� ��W�?���}�r{�xuà��迕\��x�G{=擈�A]�Q�:y��7�p(�Z�E8��>;Ӂ�B�c%c8�ą?v{{d�	��T4�s������}�ݷv�����=0 8���翷�����_}�}�����^�6��gG���QT�^��aH�&�w՗!����7+ �
�_V�:��_Z���R����m�9�@?�<��_UuD�]�JW|��O.�NŮvn/z���5�ѢެE�<`3��r��'�!/��F��W��*č����\�S��F��6�t�Qm���	��a-]��{�1�f�]�P��`q^�#���=�J�y�8�{ŦԠ��s�,�an�U��h)��NP\��	G/ΑBMj��\�Ŋ{.m�e�<8�Nֻ�] a��gݺ��_�j��8U}����`�o=�&�-��ԳA�,ȷSY���+�5��P77wvs����\��#S�mu 6��zY���}�j�h��Ъ	�(S���<����30t$�	�` a�Vc+�@Dw%��P1
�r��8-2�&�Q8l A����M��͚6SS��Oj���V�����O	��~)]��hm=U�B]PH���H9
���6p�ov� +���t<���
���g&���RH�8�m���e2K�<h�$u�O�V��N~K'/4��/�����R���$�y�Y � {"�;�ߠ���Nk�'�b���g~��QٞҔ�J��י�Z29:�*�������u)�-Ŗ�}ų��\�so�L����(Ij4M\鋀��܋�m�Bʰ�����Y��]�kΓ��*�P�}TmS��q�Eɗ+�:fsG�e�W���ñڄ;�T}�r�zqQ���I�����k3ϋ��Y�I~mu̱f&�����.��׹XU�������5��믞��+��^%���W���#�MZ�|̽��(�P�o�-�W��o��,U@7�a��?h��|'
�#�9'm����)ث�\Ȇ��Y9���ʶ+ YoR�@y�;X�n���0��EF&Mk;�
6��6�-�bE��8�l2rh�g�;���\P�a���␶b��"��I�P]&~����\=Ru98Ǽ�]� Hh58�wE�����u�&���`]0��Un�u��x���{��ql_��6���3�4n���ͣ���Α�p�D���83�����U�ײ�CƑ}���i��W��lE�W��zi7K:�GNbV��)�6��IP��a�B��ͮWb~(��j�v�6K@I�6���q�v� �� %����`�=o�l��,�e��D���+d�x��e�m��Yl����9��K[�
��OYUe�,�X��MQ�4�I�N��q`���2�XTH�S����o�P���;{��
����\�XlV�� H@ zb�}`@�����ӵ�w��F�.�- d^zo4�sq���4G]�����}=E:�I>�R�j�9 6�����#�=��ͿHޤD��p���H='�J��������{f�D���H����I��H�.slt^��S�&Bs��Dy�NC 2)<�����Ʈ"�0۝�с�"�2j ����vq���ٖ�d����SO9e��"�P�vB*]���~	j��J��kz����gO�s����<�o��i|C��q�[����-���@ֿ`���1ksgp*T�=�,�OАҼ6����?���ȃ:��$\�P6���a�\�l���݂����qp�*�WY��Q|q�=B��3��eѲD*Vt�g�6u7�����0�(��9-n�fz�G)PI��vS0 �R�f6���9��K��A�-�@�a��c�Ό��t��g��.��z.���no~��W��A}6:����f\���D7�ٝ�\``�D��˪�	���ѝ���L��� ���}�$@����}"���䓚�c����㲏�^��9�$���)������B
  A@�GR����:7��Mp-���֦`���ƭ�Mr���(ͽ�=��1��uG�4O�:���f��%\���~f�A�s�:'�um����Asb�����Gd}��c����_��傿�X��u����/�O��W���!��f��&W�(>��x�B|�=�v{��\TFОF��R/L @����y��DsUg��K֖@ ��2��z�lo�i���/��ky�����z�=N��6^����6Neq>�?�̃�Ky��w�nu*e>S����Rfoi�!�1����?A��W�[�^�Ad�d�̏^�w�]=��΢�:`��:���gw��n�����\s��`��9S]o�Y�����.PCc��'|a� ���<Q�e8��W�>��n//��y�e�^*�(�AV�J�&Js�Ll!�i�� �Xdk�W�GT
�Dv62)	5`o�z^dn��I7���1Q���#�%�/lhqѷ�+X�k`Y�i�ڇ�� [7x�1�+�܅ݐwe��A�=�v=��k�	͐�q���Vvqy�t>W����K�b���Tv�á�Q����G֞�r�h�3��^��A4�]�o�<�Îk��5I�Eqja
�z�?�0ٓ%��A��:��e���B �l����ACq����;��?��]�W�U��rw�� v㆗d�e��]
'+��'(:Y�\�s4�.��AJT�T�k�x=K[T�:9T��A���O�IϮ^�7_g��zΉwq��ΠZ��ɽ�&ߜ��(ѠK�2�A���{g�G�-"���PX�!Sd:'T����F���Gh�}&X�t�-X���6�ٖ���v]N�t�SyH��5ĳ�BwCʓq���.P��P��R�l���	�䘪x?��)U�o(�1{��Q���dA֙g��J��K={��Fa����ԭ��,�Ћ���E��|���i���cH֕��k�������˻�Og&-Ș���5ʉ�+'��](4ŧF���h40˥u���u������'q�������Va�Y���[����C�Ɲ�ZA�h���ݩz��BV=+г�z6V8�y��M��������>|�d/^�u�sn����y����]�������i��X�0{��e@�A�+�beN.<@綈.7����j=z�(+ږTc�<:��1q�e�O�M��j���!���g�P�����V�$�xo� �nKN���ɛ8S��3^F�
�A7�5,��2F���ܹ,9X�9U��{�C�,W 1�5�UA�l٩��LL����2z-���2���h
+�} �x�%�־�1:�B1���2�A�j,U�_��۸Rp�5p\	�v_��A�j�9x �7�3���� ��?�P�����Uw`�!ZКPoq ���۞�����HQt����4TF�������Z� ��-Z^�M�`������D�4�A2�*��6�/�&�߸I8�ǃ��ຎ����H�it������ P�t��Ƽ�j��@3C&
u>�/��="��ٕ��}�Y�F�M�u�B�����. ��pKg�������h����484�}�ϱ�}��Q��%�̌ �j�:!?$�7��<�زq��<�a�>����φ:��Dg���E�3S�uP,����0�Є��t�.�#�3�ڃ�"�2�T7R��PAO��t6����]�%��+�c��ٳ*�j98 �p�]�.d�kz�������H�=�����Pr�ۻ��9$^/����g���� �*L9�
��k���v�|T�*�ss,��-��L� M4��5�P��y��;�̌,��B�����PbN��,�!^3[��
)���]�@�5�P�<�H'�l��JcX\\]����(�<������J�:�q%@ृ1,�^�l;�}n�<�h������OW�nQY@˃}���{j����)���r��8�(��;yv�J���׸������Pt����I��0�#)�r���S=�zg�O�Ĝ`��{k��;���4��<��s`O��nh.���-�Fq�Q����Q� #��U6�FC1��4��
.��R��=K�&�0~j�'�ǁ�1�f/������g����k��FQ�\w���her�
���Yx�a@����;����m��ȂuNd:�u�|��J;�#���5�lڥ&^�F��X֜��'[��Cd� F�����(�~�VA�� E��� � ��Roˋ���9�g�.��E��2:![?2g��,��}�����)Ti�(�M}}W8O�=k�*f�S<L����J{~�u�Nݨ�~�~�K�j�g�kr�܁p��_���R��z��ļ�e/���U|�Kw��BO�������v��o����C ��ͭ^/���u�������#S2w��j����x-O��G6��~�q����D�܏?��O���ngW�#��w�l�Όiv[^���FuR������䥯���h8�G��)6pD���7Lz@�Y;ￃ��L�=�t�F��f��7���7�y����F�{s�HN7
�R�J�Ϻ�č�$k�I�1��y�K�[G� �ad�κ��4.����0���y#������;��O�v" �e�&_�����w�XG���?��˃���m��|N���B}���~MCG�HB���z��jYI?*�t�� 4Q���fG��&��gH	pp������e��qj��z��2x��[pU9х�5�� �t��3�2F�����.��!�a�L���~/����!8��B����E8H���>w���&�Qf �;�#*�\�m`;#�-�d�9y�W��˫��z��޼yC��3
\����P���W��H ���������_�c��O{o�>�d?��#�������?ٿ��_}�P^�g��z����\�}�=2���:�吚����=[�k:�n��g8v=�˗/쫯����w���]D����rz%��<����೚{C��H�+ �p�?W����'���!`�CCY�����~f�-���b*%9��>���j�&<c��L�
���=�6��jG��Pa�`o��׍��� XӔ}�Lj-���)��l3��#8�m&�l�[H��ȔP����+�_P+���q���+�D1� ���z��9w��@@s�f�p�p~V�{˞�CE%K�	���L�<��x$"�Y�Z}����Q2c�{��(���Ȧ���!�=�A�s���
�Ni�XG�dZ���I-L������ګ����tT��������NaT$������ر����j{�-�]-�jN�&i�c�PfP	Q�$I�Z9�ۢ�E����JQW%���$�֔����Kl,�}���2Vo �L	;�Gΐ��Q�tV��AdS����H�4�iP�zj``H����[D�l�&�P`�r���Ԛ/'�8,q��N�C��;P�|/|�O�f��㯡kf��pBh-͖�,�h}�T?sc�Q9Y�cktI��/�u��'��#�3_]׏�-~y^[ ���a�׈��u;��	��s��Y�}�I�E�6�b%�cI��b��y��{�`3m�-�K)�3�}�����r �ҁ�%np�g%[��*>	H�4]���2�y9h� �q�Wr��h���D�g�1m�&�8�h}'s�>?��) _i ���=�lqr��#�`\Oλ�|�-�1�5ϾN^'���fN#͑ɵ�{P���_\����}�e��I�������?����7�����|�Y�}�}u��l3϶&o�����Kr�]��b��6�h��F��ڭ��G�e�ɲYc��da4 �+'6���;�!����(�w�L͇��e��h053��=yt��|8����g����ע�+�|� �����
�2;0�� /j��/���V�VN � �z��W01b�Aּ�M"x�[GgH�Q����K[�Km)� ���yq:1�orZ��TO�쁂����J�h �:,�G��F8=<Vkt}�7�f��dM�E<�T6�/�B��T�N=���#�z�����emκX{�a M�5be*�\�L��Բ]��qd&#�$���q�'�� �)�5�q��cF)o��[���-����gg���{]A��/�P� V�uX�����{
V0X�4'�?�y�~>_�ym���{�����������ꟶզ��b|�Q��z�����tN'��˻g3�=���Q,�;Q8���D����cR�hq�//٣�"�+`��_�¾�@k�/�Ï��O��޾�P�{� +lb8�)̿�Uο$]����O Y��iC��8�=U�g�x���,d�10��ٕ����2%��y�A|+�d1؅� L�P� �g��w�[�&�=�S�� �v2铢�V�v�|�'e�	A
�d��MGѬ!Æ����>8����-�j��΢#�F!
A��l)@����W߸���Ce�r����2�g�hSy���25L.��H%Ff
��6U�;�9N=c��g���UTe�?L˾�l��R��L�o�ɢ9:��:W|��3d����uBNgɱWh�-Q�U�˟b�@�#G=�A�ui?���Y�{Gڰ�Zcg���	��n�hT�mFyِ��]�EG#���y��zӇY��=gp4�=f>PF u�;������^�Fu!����ɥ,'��B�
��J�X��w�����"��t�m���㎟>R��_�F����f'�vֿ��{�&i	\ؽ���^��p��Z��Xx�j�
��|2M�	��/�&5����@'f���{�f9��b��-1O��q���������iM��&�b�(�R�IrB��? �f��&��B��"�:~�Ә���N����&�_�[��N�&�豆�ȭt�/���*��n�8�3PK �6�b�R8;:�`�������9��]�P_N��y-�&RZ�F`����4���@&
[�25�܂yZ�ܨd)�ZL�zp*����=4om�č������~��h�*���zn�tpG=�F3i��@�q����ǆ�k�:��G����L��ƀ�CE�>v����!����ڶ>)��2��MC�1#�]�^��$2/�une�N���KP��D�(>��5/q���m�C�L��"� p�+�b��F���r�O�e~:���3y�yg�#�g�<�ְ9�B��b7��P5l�j �C�bu>�9q����ȴ\�l$��ٳ~�tO��þ�����m�!�u�����E(�YL!i���I�f��f��:��I>���R�10�"V`mF9�s��J�ə-�k��%9��I�m�$.�W�O��1 @���l��=�f8�ޛB�F�x;  ��IDAT�ƚ��>$ZWϞً�/��rC�
�1hq Y?�}K�B/�kV?<�L l�����_��u��l����g;��x���~����w��/��o�~d�o^٫ׯ����;��+�yO`R��`�|O����W��m)�����:����Ƴ
�|����/Y���^�~g�2���3�4Q�@�S�q�:o�� ^�ha6�I�2+!��z�a��T^��D�*��+*���7� ���Ea�!1�s`�8j�P��ʣd/��2э� �����s{�ei-�_�b�h���Y�ew��Xd��p�O3WIA�� ?�skT�����8j��G�g�P�3~��5�8{�Vo�Т�ʐH)<g"� �j	�V�E-�����M^�<(Q���`����km��@�C*��W�r�r ��13�C2g_��ڸ�E�ۃ�q�	��.`'<+��L��T�)U^�C�0
=I ��(������Qv�܉l�`��\�:���RPS���=8ewу��ޥ��-Q�Pe��{=8ELq����Lw6Tr!>=:^�h�E�Ȉ��Z��͎�}S~�|_Ս�Յ>U��1{m��u�i�<�����]ȧ��C��gEc�g�rxƨ�É���l�����&T�5�E����Dq��Y�Úp�i%6%w�cqk�n��`	�����Y�=�F������sL�9͋0��yc6[S;9��	D��dMv]���n���@���E4c�'�� S�M}l�LƊ1�h0��׾��V�QR�9mE��S�L6k!E���EI:_�ThHc@���w��rU����H�	q���4��fE*BY�2���i��*ct�דKB�T�>����.M>\���
G�����MKo%a 7����KD�%���{s�h��[�� �V������嫴{X��1�6�Si�|߼�!D�ߘĜ�ᜇ��`��1kFVk�)��K�Pyl�w�!�3�h"�.�#�-���8� �C�D	�c6$�~L(^�j���/.����{�칽x~�^8���d?��w?}o���Zޡ��V.��r~%��j�N�`lNY��f/�MĆ¿�k�I>�Yu�\-���s�A�x*X�H�gg� h{��U��Y��a4s���l�f����5P�e��iNm혬�
6���w�^J}���rx^�m(G?-�����Y{�k+�B��o�b������W���(r��B���y�Q,s@Gh4��ʲn�(	�䵟ܝ<�+2��{�]��RV���t�\��:�*8���R�<�D�a�Z8HI�����أZ���q��-��СBvu v�����qe���cfvk(��`��[K�̀
)@��`�a�KwFV'��&��Ȁ�W�I�����tV�5�IĘp ��C�jB�5y�ʃmr@���.�0%f>���6k%���}��(��GQx4�;ڊ���:�s[�	�'��Ǖ���������HҖ��N*K�}r�k�ݟ���l���d��pi�./Y����K��o�-��~Q��W��&׈���͵}����V`�����O�?������#���1���;_A�a&H؀:u��>����]��w���6��	�T��廧p���-��4�i������׶�(juuLvP�p�|�Ӹyf�V�nށr[�cbF
�v}��K��	�N��&v�ۮ� J�Wt!�\������Z1�Z*�-!����]���;<�a��L+ob<{��ʥ�3�禂�l���=�0�V�u-������7vq���E�$�q�g��"c�?\��ӲC�f�TX��H�LԹb4�.C���h��/l�r��J�f"�h��0Mw�w&�x�4��[!!(:*�]Q�����Gfޝ\�Cc�0H��t&�J�>�� �)��Am�i�jb�V}��{��;ǲ$pr'�����X��{B橎�|+_���L�������Ǿ�s��q)9��Y���}x�~���NC���A-�@O�[;�O���:���ol�I�oS< �x$j�����ED^ݲ;-���IB�Rmz�E�{(��R��ӞQ�w﫱x���s�ЃN��{&�:A�A�'D3�J_شg�Y0e^�]⍫0���;l���F4:I�ז�
����j�,���ɉ�gx��NT�҃q��8�K��Z8��9(B2�z[�A8(�~IYo a�����T���^~�;d Yo��e���� �ᘽn����(�qݤ?�Q���HW�Q��ۓ�ԃG�mx�4u`��!8n�q8/0r�����$SVZ�S>��~"�E*N��dr�b�K�I} z��������|��l����x}��u9��ce��Ws>��xo\����מ����:���}��k���ϕ���p�����P���^Ohp��9"p��;�"Ә�q��4,�:"f1��v%Z@D�es���%�ë1�`�Z5��G�bwow�7��
l��f���ǯ�3���"���Y"s:�� s
Fv�8�HPq#]?�o�����$��)}Y�#{d]Qv�;���@�ԁ��#N��D	����s�?�ze�)�t���͕��Sv*��j�y��D�|�QЯ*t��|0u:'���<�z1����Ig^d'�0W��qh�B�����y`����Y��+���+Ks�T�l]r�i�Z��4�|K>Fa�$5`�i�<�q6eLE��nLc�%m����I|A
�\�6�5��)�x��3nN.h��w��#�G�}��D0�&�y<��͎�����N㠺#�:��%}���;��ϔFQR(y+ڔ�N�2���(�L��Uʔq@�}��%ʷl ,	h���s�5�F�ww7��?��>��C�k?ػw���~"��}�.�ի��F�T�Î��U�AP�c_�z~Ԇ}��Wv�ݍ���O��_��zxQeqo!�U ���ĵ@f�m\���#����M�ewp,����D�7�l^�ij�y�8��r\�j�`��F>��s���<ˤ_�ƥ^C�W3U)QK5�A��!����U�V*���v�� 8���Y������vql��+�|W��ݞ��7(劣m+ ��x��=��?gO�5�̠1�Ǆ0��Oע�VP
�sy	��g���U��8kfQʤ�v̡���������g����M�)4�ۗ����x�+��3ź��<�~�
]�)��H�����no�I'�"�`�vIa�:i9'خ�Ɖ�*x���/�Y�պգ�~��T�k9]]<����4|�Y�`�V�˿�*w�٬lq&S8.�}��u��@\��<o����n`��n�H1�e� P�5vYǚ
�Y���G�z�cK,W��d?�����F����hǺRl�M�Xd��t՜��{����զ���ܸm��RZ�/$~�&������	�+
�U����g�����@_�x!��d.�x  ��N6�7_����LR�9���7S���s��������Q���R+�7� �N���O�����z�Hj#�aٲ ��q�}��o�����`ij��&(��z1
x�"�*w,
��uMU�	t��)�,mV4	�\.��pWR"(-r�H�RK4B-#����K�*���l�{�5�N�)z/z����*�z��6�Y�j8��)
NF<{���Yo�W��-�P(|>�qN��ï��[K�?:�1}�bUqd���!�*��~pM����#_՝�����M'�1�x�?�ၓ���U�k�0o���ߢ_θ�Q+w�{��l��♦�6�t}��y�-�ҥtb����+���'T1�^�Σ�i�e����ɓ[r���
���on�yh�j� .�կ �� ӷO�I��
��Z�|������i/>�����K$�J�#Q ~�&�d��U��l��N]S��AM
�&zO؏ x��P���ws�"�>�f�e��E륽=�@'"(��1�G���Ή�xAv�0D�n�r�p떔�sN��S��{���:�in���sH�" vi��u�a2P��t�Q_�/K���A�Eԫ�#H�q��U6�8̘x;�`�"���֋���Qk{��ɹ����"Y���{��IimR�
�j팽�F��T�mQ�5i���@/j�*�51#�Eq�+����r3����F�o�3�����#v&����>_����wvt���1�-�92x|�2Ա��֭8v�Go^�5���C���nk>����U�u/�٠Q��6b�A�� G?|���Ѯ���j�`����#�&2h�$��Z���v��P�E���x>?�/��¾x�{�����r8 ��}<�=��8��oo��\��Tv�RI�<�:ms����{Sm6�
�bf�(厘��.�]�r�o 'Կ����١��?�?����"��^��o���~m_T�{eH4��s��]d�������w>��?����������ط�|ao^�g� ���U������ßS�Z�\��7_�����_��S��LUN�j��V ���@��%�_<#�<`�����w���
�޿���'9�H6�;�\��#%�]��n�E���dO�F?T�����m�1'Tk	��t�
d�b��}�m �P1d��R���{�nj��;�'	S�OuOT�h���F˂A`���u�f����v��ye%���>�2 (�?��
�p�H� {����}o�� ��_�Qt��$�&���T4�?U�]� �͛�����&y-�c�����jJ��N��e�B�첻qL��0�(lKG:���3�?�냾�~�����?�u�z���	4����w���?���N�~�(�Z���Ms������E�B���������7ؒ�JA�\���`��v�:�"R���'���>���ҝ�a���R\�6,E��<�u��	�B���c�g�l�a�!�B��q�D����s�$#�;�� ��j�
d�!G�Ɔ����R�ca��(6	��5#N�1U�Ns>�|w�q�h[�#݆Ԁ#Dҟ�]��>r���o����w"*��ei��=	����8#"�'uH&�ݚ�>F2���E��wS��s{�e�҃�>�@��T��Z�u|����v��إ@�v�H���GF�����m������ulC�CrP��ȋ���"� 탊P��/_V������l ��q�7𮲤�U��MA��
�#���(�.�=��̠���A�4�p+�������h&�M7s5x�"�6�<�.��!��{6�r�2T�MҚJ�Wekχ�;��|�z��`��AQ��^�3h!�����328sY-렵=Xlv
0���<p��&����YIawu�{��"�,�Y ��H��${F���P���G�A+ ��Hp�e�OHR����4��)������x{�.I��J�"T��Ҫ��=�����!w�E��J:�ݞ��ܣ��<��oc&:+##����`��Ņ�!��cGNC/,��s
s��*AI�����;�bQ���/5��pv����!(V��l�{ҍJ��=K�f1��5;�-��dR^?��	k��S`e��}7�1j!h�G�w UP���6*�@/04�fK��N ֌�Z]��.�����ѡ�úJ�[A�m��
y���U��OZ��ݭ\�}���@&�}�l-T��3F�YOǣ*r]��(���	(���j!��ZW���N�6[���6Z&pp?_���:9�[_�U^s�h��g�F��ExJ�ڡ�M�^%���㕬6	p���@2A��q%=�L�EK�3��.��J�z�`8�K�� �n(�AY����J �@�{�D^�x"g'�;�A[�l�fЌ�(�~�8��Gr������}������������#�MN��GO���7���Ky��B����4(�K�C��w����ʻ�ٸ�Ϟ��7o��W/���yr�1X?�����Z~~{�|�"�ir�O���7��7��gS�ܨMn7�_<, �%M�����ϣ�hجbz�R.��\�� 
��&	�a΃|����Kf� k����B�}D��E���}�Z
�:��(�[U����c. H������SPo�s�1����%�$G��PUڼ�R�i�AD����� q��~��\�\�ej�t�1�t�s�9>?֠D�H�|6 ��VT:���:<>b�p���|�@�|�f�oo�.��I�=:�'O�Yg���X$���j�=�<,j7�w�&'�-�����Ê0��:��1�>t�7,���������,���^~��or�. ��Ǉ��C9K�q���#A��/�1�I���X\Ͻ0g�6�R��+�{l��f9:�wE����Z	�mV��͇9�9�� ����;�Ne�A�-\�Q��\1�F١ �&٭��j�KSSBq�#Amz6���,�@lɻE�'p8U͉ �������F�Gu���7ٚ"�E2�Fǧ4�'�4��L2�����u-w�&�(�J�q*G��I6�du��o�bgY��݄c�ؘg�4kf���X���)��W��N<�l�hxǇxb J|>�W���A��Al���y�H�7��d��5#������~\�������LW2�9�<��ٝ��T�j�p� a��`(waC@j2V�	t����d�$�P�I�:���R�`�V2��Cr70�0��%Uj�8;��#��9�����a{Y���*jmH�B�ʕ���V4Ny_�cGN�W3�e�[G�E���c4���I캃�-������y��|E]T���G�5���9z��wZ����k���O;{*T��������K��t���V��遝����`����������h�xR0Q�,���N}�Vp!����;�7j��JWQ1!"ٮ�x��4��i�im�5��&�f_��IY
2+�Y�v(�ɹ��!NՉE�|�d���u��_��6�V��S:��9`x�ue$�����d�}��@�� OeZ��[�f�[)6�WJۋa�L�hl�� ���}���妹�mu_�  �: ��f����dCg�)�A�n�^��l�I7����x<��E�;Z.�>��A:��O���cfL�y�}�-(���jAg�Kγ�/�o�Y����[�,��a�@�R���u�=�T���*ݟM��A�B�k��1c,��[��R��	�����cI�6����1!�:9��`n���HV��C�T�~��V�r��ZɄc[GO��":S;^����ũ����F��?���}!g'�A8}�0fpڧ��d��`%�;U5y��J�/�ɋ���U�9;�H��Ir���L����.�<|���'��F	D�'��&x�z��y��4��J�E/���ۻSy�x"�g�\~�H��I�@�ky��<��iވh�z����}H��^��ɑ �֪�Κ��\���"��缧�Z�W���n�����?<0��J=���if*�J�s�T!,dvـ�ь5��F�XO����$,dސX��ł 2��쁲�u����hd,3mb��G��G�� �:�O��Ҹ܉'<�<u�&=0��Mf�9��!H�w{�-��h!+��� ���� y��D����f��a��j� �:Ix�� ��vG���s+�r��'�^iPtc���m��T�	%2	��Wi�:�z��Ŀ��?��_>�I�@c����!�zΆy��i�f�q��cI#�]��˴������`)�2� Yav��f�����c9��kN���kB�7X{�u
�}o��*��9��bΒל�yݙR��,
�v�'
!�8� ;,V�w��57�zz����h`�>����Ui��d�{7l��]IMl�ؖ7A�5Y/���q<!���u���5��icւQ�J��h�E׏a�[q}rl 4Qx��f+(7���RGJmI���=�ls��^��/ۻ���#� ��^C�+��ԃ����L�Y2?�������y��;<���z�;���S��.N���_.cg�V��
�,�cYPfy�l��w�"r�໶b��f}���TVk�3�M4����Yc��{�ʤt��m�7���gtl��A��V�|~�V�i���(�u��k�����֙)����Ll���b�`w����������j�<)�ȇvz��I�r���S�^Q�@������6���q-VGf7�j\�{o�$Z�4;�����,����y6�TA�`�B�!覯Yw��p9�Y�-;�w�3I.QM��22~m�h�>��8֤)��l��X����]F7�xf�^�\h�sG%,��#m���ֶC0ᐨ�{�@�t?���8V�Υ�U�iUL��1�Ϣ�qu��z5��6Q�:��d�4�4��*h�k<�����l�t>h�G���Hq�#4dWh E�R�T`D+���q���wZcQP�F㒢a�ֱ�z�U)I�u��&�-a9O"����|i�M�`����� �f1
��:������~ivGAyk�Q�@�Z�i�'��L�.���q�@�zf�cD�k�$2��a/��/Қ � � �S�*�b�t?f)ʝҏ�M��6 U��f_m�ڵ�$���g��$�_j@U�Hh�e��U�i�����C�e#5AB/d!55\O�8��2�`�r����4�^={"��?/���N���YQ����7�gc=�J������*|�0^&�{����޼"p����1KskZ�p�
S��L�	4�z�H6����Gǧ�$kT���R��[9����q����Nӱ�rtr.g�i|*�}�j�T�T��[M�4�i�m����]k�
�@�4~x�͓�N.��]a���}�'���	38��f�F���ڣ��>ye�ǂ�u���������0c�duJOU �>޿
TA���N�F$�q����X�X#'�y���k�`���� �E|'2ph
M���eN���D&Y*�T����@���AAuJ�z1��fп.�i��t,�g�����"��y�9��o��'��rO�ҕ������]���Abڑ ���M���g�&��9H�4$��@��r-�K"q4%��� |TD�g3���V(�bp�Rfs],��y�PFO{O�ݽn'��������H~n�<t��c`(��L8Ń��d�m�zy�_�Qx6\eA12Xi퐽�s�'^#7=�/85��B���Ǻq"z��]���[0����71���b�Ţ�nZ���&�Xn�P��b6�T'�^�[���y�wg� ��"&$ 9+���e�b3t�0��=�J.�hR���\(kԭL�~���H{t�Nǧ0�}�':�'�:�ʛ���D��]�y�;�[X˓=�Ci���j�I�����020�{_̾� X�O�ә�8|��8�ƾ�(�}�o�g�w��?�2��
��sC�,I'Br�N�7�RD�/��i��8��&I�HNǶb݆�_Sm�j�'f���0٫#:p.��l:���ym���N�L�'V�Մ��`��i7=�F���Z�jG���*�&1�4+��4q��v�M�{�9O]ϋt_D���I��u�ՖB�,h-�Қ��;���Y�)�]�8g��t���?��� !��ƥ2ѝB.�[Rx�m�N��yi�ZՁR];_�����s�Fm��T�E�N��
����4!�#ع��<�B��y��%*r�)���~�7*�Q��)�����.D�N��:}_�кf�t���S���YF�EP�,��A�}0%J�BV�	QI4lc"�c4�Mω����h�G�:8%%�� -����c���C/�Z�� X��|؊��v�ūX��#j;�J�.�"��UkH�Y��,E����mN�`�m�9x�fۨ��:�%�j��i�9���H�Gw��3F;���e�^��=(_�ou���$�v�P�����vJ�ʑ6�e����>Ъs�cf ��1�� .U�~Kg�`lF��)NP��J���w�X�ƪ���њ0��I������X �O�XS^;�j���(D8\,ٵr�"300�2��P*"�X��)�{��:��+?��z��ĩ�x�T�=}$�Ώ�xN84����*",+�"�٧Z��,��5��g�3���ʂn��	�e��<~tA�k}��ʓ���=�7�u !%����� 3Z[%�@7�Yh=.�5vpU�x���6�~����F���w�y pܙh�niJ���5�4���B�Vz_��WFR���"d� �eL�X\�֧�t��̔�_�<�x9;������Sw�ܫLD��� 蛎N�[N��V{�E���0V�4a��Y�����$� +X�`�Ccaf�F����5a[�p0sL0Gj�/e��z��r�6�d�s�J4$�;A������s���g��¢jX,���Oc�A%��d"���7���^�>y�&���	����#��|��?@�	�~��Q�N��cs�8?#Hh۾A&�;�����ȅ�~�:��3J�ć�8�t��G��� �����w�5;q��bԳ Y!��^f�CS�]����Q�E�k��Af���ud��n��M��8N�d;:8����a��x4K��"�=`�,(��d�,Ԩ 5R�t��f�&����e4ĠCV�Yоe%��*:AIM��;���A���'�3Ψns�����b4�U��tm	`�M��J)��c�UI+d���^�z�׆�?3��1�������������r0n�'���% �����/�A�to�y2_�6p<�����_C��a���� ��|��K*P�y0��5O*�w�|�=�\���R�b��(�D�-�!�ƛ����Fl�(���7b^]8!y��2bi緋�)ZV�(���;��+́��xyCաr"����*���0Pl�ҿ��Qmp���[l)�e��k9fĻ*-�kĝm�����iۧ��k���,��S����Fsm
;�8Hr��ET��}@���@�V8�U�;�	��x�Jq�0���
����!f���Y̱N�����G位�Ӧ�Z��n%�G,�`�mQ�U��P���2J�K��i���X!�h@��|�sэ���:�M��,���Jϖ�2�l�FSXtjށ� -A�_�����U����(��4��wG��bvĹzR��fy�7�:�ʝO>�;Jk��6X�>��Q�G���a�h�Y�і�l-h��*�,d� ��vF����
�g��a4��X�K�
�"i����gy��<{t���'TRђ�%씶�[�M�"��@����%ol�|�����(�]�T>�<�+Y-TLa��&c:3�޵J�kFn��Z�-;0��a 8WWr���|��$�9*����ڍ]��qַ�u8c[�%E�Q�lup�j�F5��ҷ��y�8�#k
�F�F��yK3�D�M��:�0ә��5f����V1�����Wlѩ���fF\Ч��}���L�&�m�4@�b������xH+{�����4��,1�[k�����k���A�S5PTF�N�9 lPjL-��D	�h��!.��O� JgsH�ϻm�s<<J~�lL���Ϳ�����#���WZ�m��}���膁�L�_5�b!`�Й�i~ao�~�s���C<~Ӱē�Td��= �!�ջ+OӤ���yM�'�B��B�s�ܷ?#�T:�j��,3��ň�͢��7(x�|�X~������K���Ed���O���r� ۴�/?]���� P8y�"���Tee�7�n��y��T:��2S�ڙ,mt�҃��O�&��qL�d�O�#�>�x���Rq�B�	9ͬ�O�VkB��b���S3XmY�h9]����U��,XL��pv g'�r
	��F���=��i���R3�8���,�eg#n��E�0NF�T�1��րQ0��z�P�7�e��Ԝ��Կ�öL�����$��~�\�f�::ĭכ%�Vq�x&!��N��m0�Z�gR���#J�spX��n����,��̑J��m��8s�E�Y�7p31G�_C��>Z^��ks��ײ��Eo8���ʟ��g���X�2���q �km`��bP�m�����7k�t䝁������hT��hC�H� �Y-��I1bA�s��sp�L�9��@��ze�0�AV�����~�:��UeXlr	�C�Sˡ�R�ket&5���/Ϳm#d�#RB(i�"�����h� +�Ҿ��,4����p��#�z��;;����#D��aٹ��
 \������5���e�}�3Y^��s�&#�)�"?��$�r�K�-�?ݶ���M�4���v�����C9=��۵A|k�P������m�X_1�dc.���u@��V�������E�;J�Pw����=#ś #�_f�������&�(P��`��q�[��[4v�As�h��G�NJ�Ľ�c5G �	dA�%e��V����o��5���!���1�:�ub�6�����s8x�6����9��"��c���{��
1�A/���}i;o�����23�8i-
�I�lTHA�c�!���8j��g,Q�u�I./�>{4��Yegq�-%����0�?���{sQ�l�>��dei�5*b��҂
� ��JN'�`�Œ�N�q�����1KP�uJA��Jk����C%�c3{������&G��� Z��&�B��z�#f�
���]#2P�V�@���;�ڈyo�K���6("v�;
͚�ue���uQP�u�_;���}x0���W��"�x*�����Z�[�=���3pP5Z�^i��cv��Sm��먡�	��X�ʱ9;"U�}>ߑ��yZ,X\�sMS �2LN
ƪ`��� t�5*#�H`�gm�I 2��Q�?��t��|N1��F���a�j��B� ���Y��~Ν���*����&�)`����l��X:�S!�N�>��^Z�@�y����	��d�!kĨ��,|��a%��V�$�i�2�{���c����6�  ��ļ��Q�@��!h��㖽A�L�eR�\�;U�Fz6�B�\�N[�����h�n�
&�O(C��J����Gm�0$�bϦl�}�_�p��^����Y_�g6l��o�j}M
�_��W�/q���r~vl�n�5�7P �Ι+�e8����=�E)�=�������#�2Fw�����/_�n����$����Fs��,W�Z�F��1������Mض�EѠ61�����'�{�*j�53a�-d.�lp;mr�F�X�>[S]���jݐ.�^7Tc!m��Z��!r,lc�ǐ^�`�I����ǀ���k��+ѢPJ����u��"����dF?�R���Y|5�n[>�>�5Dy���s�A�ON{�a��_�wZ�0�p��2����S��_Cq��_�W~ѯ��jQ����}��nޜY���K�R���V��t���SU���Bθ�1|u��B��ju$�ʟu�evwk-�[��u�
��R�p~:nk�KU��Z(Ͷ��S���ri�Y����4u�	��|I��B��u��+����}�I��O��wF��~}~3�Vb_�Dj�����S���g���E�!)�s�i��?K�ӵ��5EB�`�)����$p2���K+�./?Ύ4 -��p�`_"�;A�	7��<�ˍ����!��C�(R��� ��[Z(�j�V:ucCg����G@�i֊�Ҋ��e�l��7�D����5 �{C M��̕F��U�:�Y�
��2_є�(��w[#]o��^�r��H7�D�%�5�ҹ��� ��rwG�bkM^�@���q U]�y|9����������DF�Ql	-a��6��������^"c$�Z׾��l���D{<i�F��L��A���C��Ĳ��A�I�MkN�%#p2������9 T�`��ViǨQAV	Y����9�n㎰�Lwf��4ۙ5�r���Z#��8*���yq�X�A�Q]86�*�JL�~Gz|���6$�і���|�UhDF��@�B3ˠڍ������qd�Q#��j�ܢRJ3��,��j�ڒ��FWwU�۶A�J�U��ݐ��X�k:����^��o�&����=�KϞ=���f6n�
J~�z����o�ؔ�:���*��N��(�����y���l
D9p�V)� >��q���zT� �]:���%�����S�L��C�v����Ը?'�{)wk�	�}Z37��JCH[D�Ĕ����[����.oT������錉���c
Qp��"݋�f�X��	���� ��C99:���c�5���(@Z뺡2�Yr������O���tl�yT�I�ݪT�ku~3g&�	���>g��O�36d�\����g6��2�G�A��b#'��2���*��U��*���/�(\� �nZ�x��2��m�����f �P_��(���(��P�G>MB�S� [;FtB;���v�cj��4�[#�8},�}�6�u,8�5�J��ؠm�^��Iw;<d� ���0�Ga T剹�I�]��j�W�wDӛ���֢$*ҁ6̴��1�Z���pv���L�RԜ�-�yT�cX��P8Ţ�Fi�W�ܤ�I�57%t!_* J�h���;.Z;��JJ������41�͂�#2ZPX��~l�i��B�CUŊ�I������`gi�P=M�XIZKLCo)h�j�&9R�0�-��MK�_^X��zU�,�Q�+Y[)bdFj�X&��e��A3_�����A�fyx���g-���g\Hَi�ѻ"�a<�,�e%Bg��-�ýѨ뻨�!|��>���h����r�6�#m�=����!��0H�.��'�ڍ��O���F��5Os�ȏ#6~���s,���}����Z40����Y�%d�י"6^lB��РFF��l��x+Zͦ$Gb��z�2.�i�n�Zn`i����P��`۔�0��V��>���i��c9N��і|�6<{��Y���ܺf2Pl5���'X-��M�[@hFҺ�,;�Q��� >�O���P���n6V���E��)V&fS��F�ץv�k�@C�:���2������aT:���]��
�`�Y.q���y]8;�7`A�����r�F����<�J���5�,�v�S�8<�)�E���4�[Y�������I�bk �Z��~"ܾ����z�p�iʆ�▋_��.��3h֛�2�n���K|2s�Q�������	6�mM^� 3�"`#hK�w��#_��R1��n����<SĨ���
:�ɦ�
֩s��fCI	�H7n3@����-���VZ�UjE�#h�6��׷M���cx�3PZW�A�2(�&gq�� ۆ��Rڟ� i��$d0��[d�9���8%�?��xʄW�%쬙Y ��̯Ws������k�-Q����LN"��SԎ_$��4��N�(9l8od1?^���\��K�# GdA��5	U�3�P�vY����Eor��Ncb ���`�``Tz&VCG?�aM����~к0��?������XB zT㘈��:(c4��i`����&�#�$Grv����9ە��Kof2_) E���7�����5ޑ��]�Ӵ.৤c%_b�^+�06	TBX7���4��pl�=�|�W:'Rlӽ�p{+���<y~&��Cy�h&��6*����Ϸk����L��u�SL�0��iF''����������n��rzv.߾�	 N���*�S��[m��I��|�����LQ6 �h��'����g���$�;��:���E��k���^���lܗ1У�3&pm�!�x}uEq��W�	0-hN�N(���'�:z4�@��2]�?��Ol{�;M��1|p����4��y��q:~�ϥ�� �X�Z淟����&�߿�݀�ۛ�0��� �BiA|����P�Df�/a'Qό�
����e�6�gVk�ʤ\w�>Z���:���b�L`l��e�e��/�	Z,�i����)Nrt���	`M�ؚ��6_5�dBE�~~���,�$�{����w,�*|���������^���	�NҞ��4 t�}�9��-����Ϧd�,z���� &k�E��R�V	}BY�a^�<]eK�A�=Z�_��4(~��9S��l�� ���	���N4�
0rjt�@�wڟ~�g�_�]����� @������H��9���׽�D�Ɍ����|�v�qd��kC�&�����2ݏ-3W����x�;��#ǈ�B���耊8(�%�*�	�6�����ݐjS\�v:=N�3����	#�0�E1:kp:Z�n!bB�G�*_'	WPJ+�I�F�b\6>���qK%��N��K�"�(8Zl9Ʌ�t���7�5B�E�h��^[��c�Wv7Z>��C��^�;�{����2�Wy>2D����T���>Kj/ۿ-�*��}���w����p���]_do��_k9L3u�/�b�~����Ȁ	&��yf���72"���2�Zcg��J%T��@�0Q�����$@p��󅜢� U�&4��A��f[m|��31�2��$N�t1���J2�S,,�v�0��<L%/�.�͊���1��5�eW��6���Ձ��bfX$v�vY�Z/?���}�JQ���Jm3�n�a8��Q=q�>g��6��mB����� ��琊Y�L�۩�,�k\}먶ə�mYc���N{9Ū� �T���E����gn3PjSi6�d��d�j�A���Ӥ�F��V�
p���6އ}r�m���\nd�LRY�4tڃEkִy
�+�U�v���iJ�a谴&�b8�F<xH�m3��T��hw����\��'L�G=UF�+�ucHkX|�R�&f��\�s��'v���*�ت�U:�c}�^M�
�t&8��n �:��.�~�&b&,�Ϟ'���Ky�|��G2;��o�U��+։�	�X31�eԺ�~]#���
vi���9�z;���d���E��Q�γ#
P^���t޻�Ke���ݖW4��1����Nhܷփ[]�%.\�����pJQa�4�!�\+��=-�\��j� 8j�P�����QJnI~�@#M�t��`���[���Y���k��O?������)%ͧS��ӟ.?˟�����x�~/X���(��7PZN ���u'�	�ӽ�% q!�	8��哜�$�s+�6y��g Mw����׎q��"�>O�#�+ d��$���s?���oTM�":O�����x�'�g����VlH������k�I�lXG�d5i-~�����Y޿{� �B4c<�x"؀L$�!Q��dv4�q�#$:L(ǃ���ŝ\}zϹ��˩��c:���i��H�][;R��>�3��C7W�˲��������c�Z����T��!k��֚D�x�}@V�6�c�LPi^�|�$HRz��#e9��Y���z�@�r�`��TWpj�	ܦ18H�i��Xggg�(�9��4�����g�Wc'�a�P�A��/�7u����m��[��)c����ɕa�n\���]���f��E�w��)�R1p�Dr�M��@�L�&�X��0<4PҶK-�ꤰ@P��_����/| �=�>�o���ڷ�|������@��%8���T-�&u��VVC�@4~ EOȷC�]�v�g7z���i/sk�@����
j����]�ȠacC���J�L!��^%g ��$}g�4;6`��rSi���V���(�< H+��-��Ky�Բ�R�8�:�FR�Ԣ�J�	lr�5'�F�a%z#�k�V�bE��@Kͨ�Cfu$�T̝9�C��� ��>�#�)������{z���r����p��d�~���!�����������K������tRWZ�x�\玑�f\���n�ܘ�0ص�1��Y���p��E������^a��/9���ƾ6*�2߽��A���[�w��.o��S�3xQic�˼�l_�Z�`��=Ź2��/�f�9խ��pP�uW�ch�$��D8�8�	Q�D�>q��\�4C�:XsҹNJ틣�6�-��Wu�A�+�X�P�f���dT��L���1d����)7T�pcY�&�]@�i,�y2�h��
����;�l�X��H���6`��wgT����ȢTg`��$��^RJsގ����8'U�v#�0�e�md�)АP�H��"�\m:�N�]�&;y& f#edu+J?�p�ٝN\��J�{���YZ�e6�2�ZT�Z,<<���Vo�����o<����m׭{�R�.M����VC�=��	�Q�
K�2��)�{*��a��*�rk'S����ް���8��>~����tt�>��$�Ը˫O�e!��s���z��-A�:�x+ @�6t���Yd��m���w�A�(8�8Wԉ"{�^j��'z�^?�k>�w��6T��0�}����{b�N#��]'B�Y�ʬ�׏�Mbt��|�\�n�NL9��r,6*m4��B�>�MŐ��?o����A>|�$��������"j�'��_�_��Or{��z"�{�)C��7�h��|>�.���A~���ȉ*�L�z��u.WkZЌ3���(Kڟ!�9c��������U�=�	Jd{�0�1=����;���t�w������6�Ez��-P���v���Ž|��b�a�&|��g�( ����dG����;b�'T��g	 �M(��m�緤�~�J�jca��k[������马ނ��@��G]�L8]o�5যj���w�h4�F.���镶K������ky����B���D�f��Auަ��$�Sk�H᎚(�V�/P{���UjrG���|�l���Od�z,�d����t�� �q��"n=��?g?:��r�;:E%{b���㿛䀣`nC.�~�V�	��t���QD���v��p�tt�lt�M�Qw�Y,i�0"&�m��0D3���r0��v\�?�9���{���1 �=�2�;�����6��`nI���ne,��z ���ez+�[#Z�ϛuj?�R�^@;�j�i�.��ɐ��;�0c]"�3K�C#�@2P�V��B����8�@���G�����8
`Hǫ��U<��b�v�\em��2ʛ8p�����C�����EXFue-H��;5�/�̻��:A�`� @t;Q1��fd��_�@jS�#��_!o��Q����/j�b�_g���ݠn2�2��~��F����]C�;�! ���8��_<2�⩅����z�kBr��h�4;����x1�^��/G�ՙeƤ�z���\�]�Թ~ E䊑���{1:J��j���Iz���_�"�z&��=rs�!r���w
�	�hٝ��`�Z�����@�^(��U D�����#h{�F������g����:*l�|��ǌ1@� îN�ۨ�B���hBux0!��l�xZ�� Y,���"��#�Ƣ�q����ϲ�pD��^kbǇ��<��pN��B^�b6�t�D�M|c�&���Z,XK�|��X��S%?PI��a�?��0
�ם�Qu�LX�V-�G�ds㴢X r�����x.	�;����a��a� GLv��zێ"	�UeVNk
mr��:�_���.��(BbuY��yt�T�C�"�����`�``���V�:�y禇�z	��ֲ�>k_*o?͹��ɖd��D�M����f{�2e�*g�X�y��^����vN�(P� �"ἡv5h�
�"�r�W �h̊�Æ+|�A�1���:�]�$f�*.l)R)�7@s���1w+�Տj0�w|WŚ��	�Du^݆Z�Bg�
�[�8������:��d��~��d���F�2~B�׶5*?�3�����)]=U3Y��TF�iP ��[*���}�)���ׂΫ���v%�1�f��SR�j���E�������U�?-�i�->��**��Q���&���.}�ͱ����G��`\T
'�˼I��H�h��_ɧ�[�OB��N�����Ǻ���1S_U����T\i)��
TZ)2��(��XD�X���6bIq�ר�L6�!�5I6*�Pʄ����=Vn�~��1`Ϸ�3Ɍ�vk}� (�·=o�\����i�cg����ю�S�=��L8��7X����D� "��p`�̬���e1�����7��f��k5 �k {��cߠ�Zg�Ƞ���-mc��b������[�Z�V�3��Ԗ���6;y��e�7��u��t��3HsSE(J6,�k4+��S�<�dwlrW�P�p4*��M��hu�ĺ-X�W��δ$'O+��`՝5^��
�z���>��]�3k�m�ip�'k�M��}p���4����}pI�A�m0:���"MpM�@�*���y��J���F���
Y��q��'�"�x�P���X��3Y�h4w���v����;� ]0m��N�[7U	c����Ԙ#s�s�.
�g�zJ�6�o������/XĊ�A&�g��z�*a��2�!B��G�zB��'�2jEۮi�)�g�o(�E��P�tK�R/
YX���s���@�׎ͻ/������U�����j	f��?�`�%ټd���H��~:e���>���/�U>���L�Dx2 �!-��4F�)��F�Foa�Bz��H�~W�;��B���\#{�!8�x?8�?����������e�C���P$y�QN�^��(X�]ok�Y���l��l�������@�[���\����ޜ`g��y9�B:ȯ�R����t�ڗnbi�����ŗ��'�5(<G��ON"դm�I���y��,=����	ս b�h�V���� RY�(��'��L�p��J��Z���ц
Q F Ǔ�cn�O?��o^��x<g,�rÇ0SeE��H*�D��FY�ͧ�e~�^HKЁ���FVh�ADA�l����f�9@w\�dbsOߍ@U��� (]�*��C:�{����|��M��Kr�Y��J�lakү"U�Ƥ>R�-h5֗]��4C�J��Xs5t���Z�����Ev�*���"M��p�x�Aoqt~�p5d\86N��b�����6j;;���536��8ŮQǞ�m�_�uZ�ʩ�1~��T��{rAg\���Y��V.S�Ҙ��i�,.W%��I�v�$
Pb F���Z;٫����Ԅc8�p�1� ym�=%�{�h`9�^�*w����]WZ&O�N��uP�KI@�l�$
���5��i�K+)xb`����JH!m����:Q�����!���x�ǁ]G53]�x���� ��~���0C��]c�N�h�6PJ>�6�b�ht�yޘR��%�.�ad�!ʶ�Z���"{����y��������F��N�u�cH��9CѠ߽31�uc��0LJ_�r`�E�gb˃�7�dQ��'�>ٿ5o��ժH�� =lQ].����@	��R���Сe���_�)���.(t��Њ*�U쓦��c�s�p�j֩(�i��X�G��p�j�=��c�[�΍��z�{d��]��T��/hU��m���Z0[�"Ы-Vu=��	p�o�5t������:�7ݻ�$�S��(���]G�ZW4b����Ǌb��>}ͥY�t;��N�W�"��pQa0T��eA�� �cq��bU��	0�	QIvv��jejjr�1�~H�{C�����?��!x�V�D����D��7Y�������H�H_������L����^�]e���_f�T���.r&K�,Jkr����=ք�B##UX*��@E���"��x��.�a�=4���&]��\U;B; ����L�ir�N�X[�M`! Y��292'r|r��$B�������>$�e�r�T׊9®�_0���R�*$���e�Z��ȏ��/�Y�+J5� �^�38�Q�F(Y��(�6A���u������E��y0Qc̳�?){K���9���̂�?oYઌ�����
�Ç:�p��l�׺ƈ��.�Y��24���F�O�9�n�J��=-��K��h:�1�\}t�G��Ǐ�'��̐����Dj�Z���3���t��zv�Шv���Uqj��aѺ��H�^d
��R�o��ʛɪ0K����[��pq�W,(���IQq
�S	�q�hf���V�<�̞�*U�#M�o\Gp,*
a��v%[8T;!��� ��x��C9?9�W/�����:�#(aU��-��V��7�9A �J� >9p�:�G)�ƽ]n�𞠆���[y��<}�B�={*O�=��tftLjH���$ODr?{0�`r����y�Z��"���+������m�wcl��D���u&���,M���O���L6��j���%]�!�9?�)��cRV��v{����\߭�a�rԺ*��l>��%`�@hj�Q�OP�f�"�3LA�bf!t-���N��Vɹ;*;��]���*<��(�:��aE��6��MՕz`��+�S�G��J�q	"�}�S��Z����G*�1�?�Ƹ���5]��m0^|��Z��U�{)���cu� �����Q�A�7���FUt&������P��'�u���Un���� x��_�D��j4��X�ȳ .ТM�U��L��Vm1��ma�L�ej��Q�*Z��ې���t�`23���^=�D�g8��s��W��A�z=�:�	�p`� �[ ������h������� O?�	 ��5̉1|���%�G��g�zO�����	(�4��Xk�lCX��o�5f�ڶ�Ǖ�`�`a�6]g�ST$�pI����nbA��|$\g���HA(�2)p���(��G2Bk�x,���Ԑ�N��F�-G��L�>��X)��L8I���:�lNX���>�+�˟���Cn>_%;��ثw����4<�R=���RaS����"?�9��VF��a�����v&��}��#t��nj	͢5���(L���2Jr˞�*�n� �j�M�CQ��5$�`ɸ_�R�>���Jk0�=�z?%�H�FӋ��ʯd{�a��)�d:��^+���0��ۏȏ�fG�@���*�ER@�iS��?йAŉ��C��	�;���JO�@�d����,���}Sst���
_C��3���||���gV�˦�wq�H�S=�fP�5�	.�l=�"�z`��1|rd�Z��Oe�[�.�i^�7VG�g�9AMe�A3:���2r昣����V��&o8LWr��Q�� 56���˻wW�6=?~���&�� y�j�uZ��4�l��_,t�H�9��n��s���%s��e^�-U�_�ʋ2�J�
�v���w�ϴxV ���f�\qp(�݃2�N���z�E�������X3nϯ�[9G��T����׏aͧ����� =�4<���E�T�f
Џ��D�d���L#\]\<b&��v���L�v}�U3OA��Q�Q�F�?�r�K��Bћ�*����?���x#�a㤅1�}�Qچu���'����Zo,����u�ZCѹn�i�Y�Z3G��5�1��
g;�>��UhK�**�*H8 �o&�NA�0c���|�(�-�����B)Jh��kٮ��@u���flXT�T�OmTd��C�s���y��[y��[y��{9Kvh��UW̠PR�����n������&�UV*�-���]��ݵ��	|�%�u/K���1X� @=Nc��M�V#��B�����ʱqK������=�8�A�}X��ѽ|�z���cm�Ȇl�T|�fV�it�*so8�,⶞C����;��J��X=	��XkF�m��dQtJ��{e͚�ld�$�t s�J��L���@��tڛH3&�6�w]�]c=�h�kĢR��]�� �`�@�``�6���H�j��u�ڥ��p������2����	�Bk:��ܸ���!��G��kY|��(u���|vpH�q �5�M(
�Z�5���ɩ�_Q�32�JN� �(͵0Ik�
}0��>������`�N[4\�Z�Y��-WO�\C`��U 6-P��5A[Q�4s��l��ep�Y�FY���=�Q�E6v�+�4���w�}��Z���� ߥ�gg��Ĵ�xB�Ay�Q�~H�@+�]d� �m?(~0f�4ځ���"��v(-�MP�����3�:z1^P[�|�U/��Q�:-�{��BwA!�dS�A��&b!�0>` ���i,a����5��1�z�bT�5��5��dCi����#����-_'@I_�����/��7��?�k������[�.t�ѵ�Y;��v�.
������y�!R�3�H������5�oo��gq߼��Q[�N~Y���{�����w�3?�7;�ē��Y��a(�á��;���Q�D�:𵤯U����/��G~��4�2P�Q��Z�*���?�(��>H�aB�q�J-��.��}ڸ��?�/?���lnwϢC8G����o�������̂MqT�q� Q�Y�̠���߀~c����K�7|5h�?�3���U���X���}R7Tqa��r�Zl2�"%.�����4W��=(5���G�iT�0��Y+Ů�,~�6�.drwA{)t�T3��#U���]�	 �dM�,��hJ���O�����q�v��ԬC�#Z��Q,��Z-l�m�M;�v�Ekt�UC�7�,B�C^��A�#d��p��!|:@VD���v��j�O���X�9#�3�2��Zp�:0�S��� {�s�! ϳh����Z
�l-�HB����0���g����� ��#�!��W�xvE�B�2�f�@kVXf�̒����N"��++;\�^9�P4�i!���i��ݴ[rϙ�5'������jA�F��j�qf�ڮ�G���j=?o��=��Z���Ͳ�s�]Y�є@,���	
V��.XƪS{ ����-W��f�%DM-��&���+�8B^�XO���5�(��'��Ӻ?�Ӄ�LF��:;9���T�)��2���N�SQ�'2�=Ԏn�Kޯ���\�Tȶ�0�1��ߙ��=�g�_ɷ�� �^���EHJ����;�z*����Vz
��^��O���񟡒 9r���9�r|(����nd���~tE��8o��!�(�`z4UF�$Y�v����|���!��1F%�$h_ԧ!3��0�G����Nhq�l��"&��Q)kKጒ��l�RU&#�b5�����K�SK�8�zN����W�u�uk"M�d[azAʨ�G<�m�
���@�u�q��H�d,���)��߫��z��
l�l���$]��{��VIy(���s��,�8N��l�j�#�Z���%�|��b�}��b���unV�gb�����`a���)1�;��ˇ��BX����Š�@S�����}�'���ya�̥2�x�~_��[���Z��׆Y;�Vi����&ݷ!�<� t[�,dS�NN����A�͵wm�a)H�g�Lj����*���Qt�9.��>�W��ʷ߾�Ǐ��*� �����g��A�cA�ɤ�@1�ߨ��6[j��}�x���1j?4iOV�]��`"�* �2Ȧ�A�� +���6�=�%k�pM�P��H(X;����R;	�;����E�%0+�U:�a{	<to�z���N ���l4�J�ҁMݵ��'Ѕ��ސ�;����֟����Q~��G�a� )S@���.��j����0�.ь�,"k�H�Ek�+�X2A�
cʅЯ�kgk��B
�
;�s�A��*�}M�G�0FkI�����A8$�
����A8���_p�;��v;SGU�-�1R�r����I_\?p |iz�}}������6Odgn���q�MGL��7\����`j�t�����Ç�����"?]����iG4!���w߾�
P!Hv�B��$�xR�r�C<�g||(�Ƣ�&{��_���]6�n����i��۵�,�+�SR�r��QL�r��y�$B��K���|��P܂y��8�56ݑ�P�_�I��a��Ea�M�h6t�&�`^���Ez�O��x�K��F,h�X+��b��Ί	7�Ҳ�̊�:|Q�}��&�,
�`�ǔ5-:Y��0�ꤧ!����F&�rAĶA$�3o����t@�g��F��w��d���b�I_8_��df�~�O����b�n�m1X�Q���y����׾����Q��i�M�z�5,NG��3@Y\�2^E��)��5l��5F�y�"�5��͔�Zx]�[�ahG�Q~w�)LL ka��v�9nûi�?�8�p��7��;�xTɱd�t�;��8��6-Z6�@l��yk���\$��\HKsVt���{Ym��o1�J�ʋg����󉜝ɤ
,,/�gkw��$wr�I�n.e����?J�E������;BB<��:��Y�7;���������/�ȓ�/�L�(�$�壒��"R���XѮ�'�`���ɨ8x�V69r�Ar�K�2��A�u��L���F���9�xNB�/���N�N�ڂ�m}�� �7���=;��Ё�TTh��5�t2_���pj���[:�*'��!���R�4:�9@�Q�:�G��m-���W���T���mЛ�9h:[�5��"Nbr���aB&�5��B}_9��0���-��*pC�f� Ȕ�{FG�-�̕l���5�d%p���*�����Ev��,�������^Ώ���ϭ��/d�j4���D 1��7�-k:��I 0�R��~�*Ӂ=��k�0�b�9>>N��r���	��h���-*�m��B0ə�?نe�2�I��]��ߙ4�f���g�JY2@�Hq[���˪d3���H�_U�C��i�%-�X�J��j�Gt�qI�z�9V�������_��+��qkI%���(�>����[i��b�'il��v��74�N�5M��#KA�'�,d���{eu>��Jd�*��P,��.�-	����g�.P�[�?[�Cb@@�@(a����:*��^<��v�����Q��18�� �<e핢��v��,��-�haR���QZ�| L�҇�N>�]q���?���ȟ��o�S�>&`�+k>M[]�6"� 5�F�S�`��2-��@vN�I XZ;��`�D�i��( ����q�X状yo��[V��\���~.�/A[T2Ը�&Xw?c�!�Κ�h<�ZcGA��	�hF�ʑn[�~M��tsg�M$?Y�Έ��u��{��FGPv@�݂�#��J���?}r��Q�f�Q����gy��=���?~D'�+n�H���$���UH(��.cN��x�*;8��8��GR�������3 �k�<�K�@�/�(42z�P�eMp� k��=���֓���9��PJ�ҺE)�����5�Sht�Ƿ�_���YH�5>kj~8c�J�����)i�G���"[y0K�1�b����|M��0�������,H�x��i����j!���um�����t�ٲ�sNX�J[;�6w���Nc�L	��8�pbhv����,���VD�}�g"r4j�	�h�f�O3�"�'��f�t���7��IΩ�|3p���|u𽬚80������E��.콉5������<]��ʞ�jf�B�c�� �9g���N�YT�'8�&7�=9`ǐɂ��ё�# ��m���i}f3�Ջd8A&Dệ��l�-�Uh�b����p)j�F�kԳY���&��{�jcSH�^Rn�M��?�  �]���j͗��7��L�N�P���ّ<�8��O��:O�>fFr�%�?ɖ��b�XJ�^0�5��bM�J�:R-&F�YA� ��3!��:��l)�	��N/�ￓ����7?���S��3QYR��2P�6wn�Y���h�`;�v�( �L5K[�`�	���L�/��u��<W �F�B>~/�NI*��U(���)Z�D��N�UVEB�Wh!S�z���\�4(�'e)9�� �Q%��L��	`��n��{ �->R��~/P$��um����R!b���F�)�(5��ʭ�q-�&hp_�PeJU_��j�X�u1 �͡U���<�P��j�r�Ny���B䠳�(+�3"��"O��$]`0d^�{x��sۂ�e[Ӊ����N~�����?��ꁴW��|�p)?�����>h�	#�U����>E#=_U���^�d�(ru�a�n��WZ_ ����}�v�Ec��ې��Dag�L[��lǾ����<��Gq���X��o�ބl�Y�M^�fV�&���T�#{	� �������
��6��{/^��ゥ"#�>���;��l�{y)���t�'�
MZY�ZnŨw��XY{�g�iSun!����e�!�O�=��G�� �`Y���o�s9F�)A��e��孓_��^�i.�n�m�a;d��M��O��@�JKnL��L1�Y�#��T�m��$���GѳVF��7@	·w�hi�ˇ��!�_���˟��T�D��N���Z�v��62Xl}�r2#�p����LP�"��UU��Ni$<���y�����X0�H�DY-�=����P��	+{o��'�/���,T;����Qq��	i��(�`�$��S �%L����k˾��;.�t��F��G_��0�J�gʒ{����h�{
K�q��<���)�37���������UYGrz2K�k+?�}+�ӟ���rww'�(&i��Gl��vr~*��|a
b*�j'mT޾�dh4�V� X9�	��Aj(�Yꍴ�{�XEC��a�E��D�0��㳄���M�D\��W�ËeP�M�V��d��y���i�_�ns�����:ƣ^S�P5�E��������A*;r�uD���(� #8�bsFZ���׎+*AG�(k��@�<i�s���N��#E"}d�H�wy/Er�������*a��p¿����$��Q-����4�-��x��O��ZF)u�a���lC���r]��T�j��t<��V� 42e��G�j"��u�QA��h؀��\l�u�EYO��Z��k�r�&M)|gј������|Z�dY�5�xO6�<�!b
�U/8��ۅ{����T'�N� �Z��w�!���a{��͎�?������.����p��Gk+�S�m�%�4_�5U����i�ک]�@]f��L2VX� �`�n�@��"�]��5��3�h��x&繜�ȭRuI=9RlD3h�eF����z���_cU��l#��f����!̑J�����5-C����a��G�jv�0nZc=Ś�� i�
2F�k�XB|TEn$A�r�ݳfvT�R^�M+h��{��g��JDΎ��7���߿���<��g���AХ,����Ý��H}�5F�"�t��;��t$F����^��-�꒶�Iv~�i�*h�'�����?��?ɫo~���s*�-�Kޗ������ߗm�.ʁ�6�u]�����t�øl�!�^F�YDSb9�V��P�i-w ^���j��_#�er�@튁s5f;6���z�5̵��Ls5N��Nc�L�%я�8�4.���jk!.�^7�4skٝ%p5����t���M��ɑب��s���y�#H`' ��8t��/���:�3Pg��'��ڎ�
�5�q��fhM��lI�yQ8�FM�y��WF��ȯ�u��V��xĞ��>z�x;��m�"-�!Qߣ``�5�U�d�
���͟�6yf݇��:�\��`��9�V>�rF����^޿��^�I��o��SJ�E�����a� �4ُ��t�#�+g�"��G�j@ǔV�Q�'��R |N�&���l�l<�9 �!ˬJ�!�Ss�	W�s�Vx�Y�1J l,��>��6,n�F�~"�ߤq�Cq�IZ���J�m�8���<�M:��ۅ|���OW�䤎�NKPj�4��+�]0��h�� D���/f��6�ÀC�V��]c�&��Mҹ�Ҿ����1@[K�H�e����6��dsf�i@��Ny��)z�u�d���J�AǺ}�FĈj���5RM���W����>�'T?���~s~q*�_��;i�P*��-A��?����?ɇ�i��c��,���A�t���PԈ�8\҂�5"2��*�X[�`^�Eg�d���j��a��!ݷR�m���Ϡ'��r~+��,��RV��	p�(���7����>9Ns�ne�>MG5ʂ {���$�7ų`�Ɖ���=��{2k�B��Y)J���1.4�5�0���B�Ae���K�4�Æݱo���WBK�[��;e{���F�GR<������;��1'�^>�i>�ֲ]&w���t�"�� ku���������W��2G#k�d:!Nϖ������\�G�X�t�������.u��C�������?HĿ�y_��r�΅�8{t!�޼�7�|#�1�㷦|��"aJw
�=ͩH��_>�{8�a���c𫿇�7痈�}�ޤ�ϐ�����1��#���=��D$���1
D�:��;��ҟZ����+4�Xj��":#�h�-Z��ĆM�Ա�AdE�,��Z��%�	�ˢ�����oѬ0RDU�<\zV(�?�������p��fD��)UA2�� jA���3��o��IǶZ�рT:��R�2Q�2	C*�1�C�E贁'b�mH璀��i�%�W3��X�S����	y��a�Q��(�!G�@0Չ���}��?�[-�q�o�"�a���t�i�.�[Ϫ������h��\���'��U�d��@���΃I1�0CK��d�7��(\�Y?��,�� P@QP<џu8c֊�f�U.��担�q�)b��!X}�Sa��k0���\�F��vou��#\�y��Z�Zg��R�t�����X#e1:�X�9�y��P�P[M����m��X�yr�/���G��y��Ϟ>��O���`L�Ӈ��mW�����c��YC�z�W-�/س�O�.���C��`��C�{��d3&�����ʫ���w�� O�>g���V7TJ��V�{�ldJ�:��3�v�����Vf�;s.Z:u�@�0Ƴ�.Ο��ݍ��8��d��Hf��b�ϊ٨�Z�C��)x�<c��m`/���
-E8tT~�c(Ҁ�zg�h?����[�]l�n�!�p���磔%͖T���� ���	6?
Fߕ��'�#�G:��i�F�8�,K	�5�C�j�X��h�W��S�-��
�ISݷP0A�u�i1�Nqk��tu�r�A~T@�y�h�h����1#���M�����������  `mO&%?� N�@�%$�a����LJ"!˧29�PIn���e�s"��zZ8�d�A��~��ǰmY�5�/T,�D� ��X.r��`�Q�d��b����t���*���E�[��&Pu)�o�q�߾{/���e�\�<�R�nXGf���&�����B*ַ����C��-�PŎ���|����LιR�G���Rf�ϯ��n����Ff�˩J�#�� ���	�@�'QwV��ـ`���H~��w�O���?��<z|.ը4�FNO��Yu��
&� ���d��O)Բ޲�A�����B<���(P	�偸���:���N�5��A_���5�P��͓wmg>��5!��l�mS?&�%�}-7�?�}�*����rg{�Zש(��c^�7�v#.T���.�0(�������DcZ,�#� ��n�E�����`�i^�������|�!�;8�xJ�L�{Vr5#�P��5t��jBћ��`&�3�|2Piǩ����t��}��G#D��s�w�<��lS�@L�"6��$.&5knV:��f���'�������?Lݪ߾{'?|"]�0�B6���@���;��?�����[9J��@}��W=�R��[3�!���6t2�y�����>�`"���L뫇�G�~dWǋ��\ؼm�5W�>#���,�j���[�V��juX����Em�R�zԌ���S��@�Ql�Gu�V:-���bC��v�ӳ�y���)�Ly���5����l��e2 pf�J��@�����iYj�(�ƫ�=F�c��vE�m�F�mP,�X�I�8q��a?8�1��>#T-��Kc^�%�q`7�Jr�h:ڦDf���<� xp�?�8���?��X�)K�ۜ�y��W��A�$�8O�۩5��Q��<��Go�~�1�x�LY�����fR�!��*��&T���q¬�nIр���ͮ�������z�@y°��k���J��#�<�\���|��>W��wQr�R���QTr��ZA���IJ�)���<��6N|�*��ٽ.�6/Ο @���T��e���ɨ5R�~��+�g|)(RYf"9��
�f�_�޴9�#I5��< $n�P'YE��=��#+����dewg���n^u�F���U��#����2@"32����LMM-t������'����3���s9;>d�-6���F�!k�,��!
��� U����l�u���ZH���(���!�P�7y_8��Ϟ�/���_����3AM%�U�=��n}Ҍ����S
*P8
���RHm�e���T�㍩om�ȼ҆����u$��c�j@�臼�-�ג�#�/34��#Ԙ�V�l6�>��Y�v`C'80�������>�I͋�L�h�CE����(8r���뻅��/�� ����Y�D��V *� =�C'V���GTe���G���a$�s/��r(]6Y��AVm�|�y�^E��t��(�D�ٯ|^#%R@&��n�dD�	]�����f糩�3�p���� �����A�m��┝��k�W��~<0����.mH�P� �EF�QG��8T6uZ�>i�p7��שc��ޞ#0��,�A}�����h�麋Ed�i����ֶ} �u����ւv�̪Y
��"�;ŏ/�/���Hَ�y�N��{��/G�֭fE;���9�f���7��A�b:x=�*K4���b��m��|���a���tG����dY�
`omfj٬�E��aǬWb�KA���	V�����A鉰����l�N���S��?�����;���0��@p���QU}��)�{�@2�����Q>� >�FF2���[��
uV����M�ƣ�4��ep�6ʀhd��Wk����|ˀ���=(�ݼ�����[�"����^���!��1���J���T���Jsfose���������&�w���@��w�#�|�C���@���>�*�T&�v��C_��P�I5`^��'�ul���c`��Ӗ�6����XԹ1�\��������O�R������A�Z��Xl��;���	OÒ7�9�G�*�������__��N��n�º��Huov(GG�r��|���9����]���mM&�ZC[vN�*���a�"IA�S��s��K[���,c3�x��u)�1iT�L��
5�<?�`���(�K���U︻�E�.��5�<P�~C�uQ�;3J����S����LQ^�PxB	����?��([��7,-$��-��T�Y���;UJ�
(J6���*59˛�4�q~$���p�Z��A���ƫm4��ҕ]�f30�jn��[�\E�L�Y� ����Luݠ�YgG</<:(;�6���D�y5&�[ƿrTb+�	F#�\<���6/3��7�灖>�2f��0�s'��4�?�?���WP��o�dC����KF��qxH7���s�8�-���jD��x����	Q�v��+�F��k6�V����,Ⱥ���������VB���0��\t��Q׻f��H[TtU�p�OW�Z'V��i'1��~)0�͉u/ҫ���C9�e��"�֊z��i����*��x�6Am+��}%-�*G�)��z��B�<~$O/�d'=�y����o����XЕ���8q}x�GjQ*~�m��R�����AI�>��n�/�xH��'/(t���K99{��}UO��\b�tƔ���[�s�S-���9P���Yp۾I�iۏ��,���<V̐�������~�8J��b�^���0�ކ�ފ��kɂ���Ek.Ĳ)�� z��	B�c�'P�����4�m�Ytv��Ѽ9�3��Kh% JRt�@N%�;��8~J�&�U���-h��q� ��~RT�2P�E��f�@r�Bm��D��1 Z��%S�8����4��L��"�gb�Sq]Fe�rYr�{^��z�Z8�2C��2�1F4�T��Uᅅ��e�TpAA����t�K�`��*�Φ�e�Ͷ��O���EN��)1�[���X���Ա�>��\-�m\"� ����	�����(�)��auS
�Ϲ�L�C�� 1 ��v"(��kKP}�	2'd�0�Ttܰ�&��z
a�t�o (�X�m� �0HK���z�����yv����**QB����m�^��0bfyD���]mH�m<b��XhK��J�
����g��o^ȿ������y�T�S-�J1�u���9b�A��r�y���Yu!wy��ڕ��<Zd_j�E�i0�������+6^���>���V*�ïZ�m���(!'a Muf_ xHjkQ�VQ�bC�G� ��^��{�·�ZIt��u_W��FIuG�DJre�}�?��Zb�?��|ŹfU����U�����;��v����h[�B��w�]H�7[�_ݑ)V�⬙xгcD�5}d�M��⠨��|z]N���0%���x��m�O�˰W�c�P����p2�T�?����r�䮯n���)\:�T�ʋ��N���Grqq!''�����>���c"Cw��|��JV�G@Jz��b��9�j�)�0�M5Y��4蓱M�����!�#���k76��\oB���XP�!����XX�%��MԆ*�ŵ]�������M�ʨ�����A,$�g�!�p������)`R��N�t.+=Q�Akŷ���h�o���m6�{;c�-��P�B���.;�y�jW7�0��Mu<�JZ�*�hV5;�G��Y���ѷ�y�h6��@T(PZCK�l���r@��"��̷d� �ڨ��fM5{�sjp?�p�2J|#b�TK��P��.t=��-����xV.��T�@�� �E�S��u�\w����nW[��O�k0���sV'�7%;"��t7�W���[��Ւ�#���~|����b�9˺�F�6c�͇A��w�@@3�O�éz���֠�u�q-:�/�]��(�x�J���+p���E���)�z��M�l2����T�1���:nĬf��e�!��Ge}T����XU� H	�������'�œs9=��������CV����C^ח*�9ZCvkw�ʲRLT��lR�����0�O��!�[�8{��/���9�:8��0�	��w!�� ��kc]O�:�uӃ$.��x�8�eGM&�R}��ĕR��\���{������8�7�/e}����-k$o�p���e>�F�Yvn����������!�O=�]�z�&;#��ԕ�h7�t�1�sEn&�tt��"��kl��B��W��(�!�5�����`cQ�-'4�M��+}^���Au��e?&P˓)�����h��l{�`��uZ֚=�`A�bZ�:������u!j0/b��J����'�a�l�
V�������3���*�:!SD{uMdgw��!�0�i4�RS��ޔQM��b��Aa��)�I���׼?p�ݏqa�}�v�o�Ew�PZ��G��ivԬk��P������Q� 5����{�����=�Ή�w���\��9	�,�l�	���*,�&Rt����Rp٩7��˟������ɓ��<��N"���u�������YD�����0+�S�����@s���P~�����˷���^�_<����-Ǖl����6��GG%�֤�ɾi����F��ϴ1u�&�a�Z>^߳_|6�j� ��n�a7�fHQ�S��.{�a����l�R]ۤ�ژy&y�䎾���9�꾯"�U'�k̞p���Xy��E��jP��l3��&I�i?8h5��<�^�p(����GH�k{�v���f���ڱ��]=���z�+�$2 �o�����h��z�+Y���0o�Z���?`�u3��Ɨ{?�I(�^��%Teł0��lYD��i�����V@��2�4A�ZM0�j#?~,/_��g9Ț��Q�g����v'<&��G�y�N�d���0���˭ �w��_�1R=��m*��H*Y�P�@�=k�)[�a�z�ơA�w�hBe���4PV�Oa���O�lo&'ǧr~~�P�/�lmH�HF�3^��d�tZD�+�8����qu� nn��~LX��(�&��aC��������ˠ��
Ơ�L�/��<�!�D�x/�ҶL�^�ր�_)dȠ)z��c��L�E���P�mub��9fp�k-D�,�RTd��f�\J.AzG=l�����^�[�2��炜�J�3�zp��`o��I��!ۧ�}�[���ch8��[�W�>J�O#Xv�������@�E�1�A�Y��/�mXC��*�$t۽;T��ʞ2�p�)#�,dӳq||� �����v��K����ߐ�UBwAд�=�Tؾ�.%+���*:�=~x��րD�����T�Y�.�Ń���Q�kk4?��TT!�"x�vv��p&�����P��NǗO��x=pVن�����������,�#l��f9�b�?� j��	�Ŷ��h橦,x��b�LR2��z�����'/(rqr�$?��5�c	���f*K�&ƾf�dU������`k��#�%�('_WN��ql�ܹո!@�	��>�/��y�n�m���:ͳ	��	Tq���[Cf�L�B��3L�hbh��@�~,�c��j��4۰�$���vs�:�?��~���E�����γӹj�h}�D�kUtFI5���d���
'�EY�*�5j�Cd�5��2�}��,b$��
^P� 0eH�<�:�X�ΥR���(�"�t�����C�M��{~�:s��F{������ֻԥ\��W�ɪ)�~�؃�����D��<����N�]��������`߼���v鞁�^޷I-�Ծa�E�ڂuf�ރ�%P�nn�$���=w��F��� `F�^�X��RFPm6+Y]#k����V�����ۻ�l������pͲ7@��2lM��Z�W��C5�Ji�[�pJ��ё����g����a��;y,� ���*%{��Ʋ��^O�;I_߫׏�wd|��f��9����,�^=οk���ȱ�5#���}<��g�u����U>~6���#�]�v�ًg���������w?��o>���N��A{��n�[Z,b�5F��k��H1�����}�P �eƬ���}dC2&U*���&��oE��pZ��g��轧l/4J{,�`hyHo{��c��W}půh�r%R����}��SK��2�T��?�`M�5�S�8�z3�~e���C�v\Q-}T[�Ej*������L�e�&�u�6��#���T�.0k^WK�/�u�5Q@�(U@�5�q��'�����o|xt �{�%1Q�~�:���g��JkuFu]T7��!3F!4�����M�k ���W�ï`NU'ik���O��^��ő��vg��x�uX�e��)�1r�Z�dh�X�6�0�)�$/�}�_\�i�#9:����x	)����eѮH!B���餡-Go�U���Yvo�,;�@o�x�����k[Һ��>�pw��WlV�Jv��C>F��l���K�oƉ����莩���u�ŭ�e����("��Fn�*�&�cn��W��p�<>	>�Փ�9b<�.�9�X�*��������R;�0V~2�虫�g����_�/}���`ϛ���@C����@�؜!���Q��A������pP)^�l����c�}|�/�k�4Ô
b�V�lYx�:�R�QT���t�+z]����;�>Bz�itVܕj]�tl���ǳH�q�^�Q!�#V������#[9�	��5\��s�������xrr��]=�g����`*�}ί(�:���;]h�e3�E	HJ�E��hm(�	w~�����ѴQGnxp�зd��/g'����39>},��'�j���Z96Eu�h�8URU�Z��Ox=/_��ӕ�f3������D?� 0Ȁq������r���^���ↁl��>�K! ��S�\�6��W�[n8��r5\c0!f4�@
^k��5��F��^3��N#w] �]ݒ�z)�L�ܜ�s�t !���93�M�T��תfCP���G�(�]t�r[�ꨓ�}"1T�i��a�5�����"�U���7v��N�7�[�\����
.�m�F�-9���U��������}/@0Ej�����`i��PsR=�49d�!����}�+�0�۳�]
��Di� ��Stj��C�q�>NȘMoor�|���Aޣ�h2���N����1�f�, x�ʭ���`ᅛN[��L����Y˨�f�=|��%�
�L:8Oo��X\���)Û�+���!p\��N	6�1��v�d�����W���sL��)��̫�P\>=;��/���W/�_t�~\0����H��_��Ї��oY�ϛ���a��5K�9 �O������"y�݄������_ :;;�Y�u%��Xd�-D�e��0u��L��S�f�E�LJ邍52���U�}��|t�JAT-RPC[�h#�J�0�ِ�SClN;�_-]k�-��T6��<��b���}�z@�k��0H���k��1�#��vPS��� ��&
s��@�;�~���7}a$��-��!���(A�;/�|�x2��i��ly`j<�rޠn��}g�0����+2�Uq�5�v�w�(VGG',<���3���%J��mH���(3�>0�	��M(��\'>�s��{Li��4y���Q�Qq����g�  �T0_0Ƞ�&�uY� ��ן�4�����`Q��C�7�ƨQ��`woJ��8�����`W�.����r	teN�����X�K�MeM)��NTi�ֻ�[��N���蔟|X.��)b��������*Nk^jSgt1�Dĳ�T��7@�ńC�S#א��h!8�}ӹ\G$UY�Z\�(�8־� 	��D�E�l,U�F3MDL��_��kg��#n,��m0s>	�S�C���\�П�'s�:V�:)�v��W���W�B(k�|�'o����jVy���Ҙ��M1].VEU��n�Rd�����5��@�5%�F�Ѣ
�!o��u���]䱃vW��}c�R�`r��G�u.S�Tz�B�k&��?���"��8��AF:�A
B_�͑`{���XΡ���Ue4 �W�c2�n��vTzl;'j��JRv
?�W/�˫/�ɗ�.�p��7�������~G6�j��>�錬�Xe'�zH^��&�s�~�Y!�X�M
ꓦ�Km��)Q���������s�8{J*^5ڳq
�X�(T�mA-�R���G}�,a� (Ҙ���P�`�@?u�1W�Pyc}�F;rx�H�/�ʇ�?���[�]��1���zv�Ҍ��Q̸$���N�~L������k�Y1���~�=�9Vt�z�Q�i~�.$�q��s�t�M7r���ۻ�<�<�RYw]iS�eI1�Q3Y�����P��	z��ZRP�"iUW4_�h��_b`A�v���1B����b�7�M� F�"z�N�S���z3���� ا��d�%ܑ5%EQc�A�$ť�\���t�췪B���iv��Is�k����
ŔD,P�g��j����}	��XM��t��4�A쏅:)�>ۭ�ÜkkmsPx�m
��!�	��(�X��u��ohS�Ze}�:��\߭R9;ͮ������з�J�1����L���x��S���f9�Ѧ�nawd�vIM�@����E��0{,;�5��ls�N���W�����Z�="�S�c�Z
�~�V~�=\�_~y��ŜA�lv�$ ������G�r�j�>��u��k�E���ގLr`�Eȼ�A�M�TI-��zq��d�j����K) #�hf(�߫���-��6�^��1� �AlX��*���n�tS�[>��UQ������*ng\�wD5?�S׸H��0��:`�v:�a��m~�k��;e9y-�'��
9h���1�ϻ��6GT8i�G�+#�Pj�d��SDw���{C4��j�Sh� -ʍDYtB(%�Rn*2 �d��
T�$����8��y�����E���q,|�M"h�:�;pT�J[�Έd��ʜ�7ٿ3��$۰��r�I�?S[3� j6%��L�b�XCI��ĩ��x�{]�t'L9���Pk g{9�B����I6�'�%ݟ�$p�̆�N���8ݵ��R�&mZ���Q0�"�+�BM����|�������L�֊6b.�6Y�%QJ�ܠ�q�	%��c��ET�T�1E4����.̾h��a!7T�df4M��\��x+�ِ�TJ>1��ȯ�ɧ��0H�!x/5ۨ(���A�O����E�:̓�\�w��\��s�.�{�=����>qRQڑ�y��p N��d��J@�%� �����i�o��bs�\�� ����KGz&�8b�lvI��yGn������:=�d��O�.�Q���~��������{s��١�3ꐑN�N�7��-5��c9���#�"k(l�_���(5XV#�}+ ����)�
����`Y�ͦ����K`=Wm�:��<:?������W�ʫg����l��cr%w�o���� ��5m��+Н����_OP�r�oq��4Z�Ջ��� �r��.�Yw����#�8���gr~|�w�`�N�QX|��Ak3v�P+��R%Kdk�;�n��v(�s:�S��K�f�h,o��w3���$��>���r;�\C��E�ԧ -b�4�$����y,_�t	874�g��Zv�9���sL�����0����a)��(nE��dG����(���A���D���N��D�bk�����o[��5����j~׼.87����4�P��o���x�r`���9m�^�mtq�b����g�ᓦ�kH1���^Q�̀F��[��hh�r�u���'Oq=]<>�ã}f] �2����4A˛l h� Ѧ��%@��k�j;v�f��(��_��)�90hX/�+�- 0��_,�+m��z%w�5S�Z�9��8dRH*k�ݷȡ�U���	����։;�x_�@�D���>��Z�tf��AeO}�W_��A�S�0`�2�g������;�Q�*�F�4�v�=
���,�z!�ԃ���￑o���\\�|�?j���+��?���{���s��^�T�F��=ր/�1���:�y��Qn���G��?��\�L����<�>����ﳝ��Һ)�J�lLhI�^&X6+��� '*sA}!�"Av�c�&Lh��
�k����<��){��m�3��x�������F�#U�u��:�
h��3F��CT�. 6�N<�꺸)��[��P޷|��SR��=s�t�9@n����At� �@�o���G���7%�Qn�d8��Uvq�>))B�`9MG�,�� VK�1`P�ӑ"Q�U�6<{�$O�/����ӧrzzN�|�2;���XhȎ��0f!�:-U��p����&�4Ca�vz�wl��4���
-�w�÷�O�����U�����q��1Z�@�3����z�/d��z��]��ą.�TY��L���NvF�g{rt�O����=�����
w(ww�h�F�uNSR�f��)��ih, Ⱥ�W�-��M\e����
�@�@0�̣�Q
a�1�-�D)�D\A��xӃ�ib�<�ǚl��.�Qt�-P�QA6mP% �QYD�)�
t�X�D0�#�!Y,��A�*QF�s�Q�n�0�O��q������]cl�*�^�J܌������>��_͏} U�im��8|�~-��c���r�J,������H�Zu6��e��_Kl�;�i^?{�A<�5�Nibk |i]@��72��i���E�A��f�����ڂ�;:C��n�%�)�?���m�%JT=)�ͭ��j�S9M�kVc�b.��K��Y�.(��b �R��VA��ŹU��ҵ�|��Dm���2X�iM��Wϳm�Z�G�.�A�k������ß���g٬��R;�Ԍw�I��Q���?r%���w^C$��|�)�6F�e�7��S�z.(�>:{��ׅT�G�"&*�`�ƙ��ᰪ���뷾�z�}��U��m)s��s�d�_ls�O�������w�� ����0;����l���N�t@]L����,�PH	��p
V��P�N:�lñ��1�Ƙ�����a=�Z1��خe��0�y�QvXSv�
��ڜq8�lI��uPvT�Z�*	�wLA�G���� �aW�uO���4+��ByH] �h" ��EY߭��A��.�wP�d��"S]��#���b��Ȇ�x�vOX�9&-Yd���||���1@Ԥ�Y��8��i7��! ���^����Dsh���w����������A��cruM�w|u��*j�+>�P�����O,m���`��s���:�QQY�����	� @V�8���Z�5�+�k��O�=�6��˗_d[}̌U
�%�9�q0Q���� h�yޏU��!�ɔ6g�Z�qzrB_-)�1�	��"��Z���?˿��?ʏ?��{�C>��9k�R[��R<a�\�b9����r�sC���Cd'�����=��|�n����'�V%��S�5�f�Q>]P��&eL� Q�^���*@M��{�BJJ�@�}���5_�q�]��94��v"�$�������eU9����M�����9�Em������ɖQ�����A�6
����̗�붾Ђ�����I{��1bV�RY\q6��V��J���Mnt�28�#ȑ ��t�:���tvJ��Ⱥ"gp~v�h�J"��
�_}�R�ǿ~%_~�,�� n�c�=��M)jSw�^64`	�V>�)hT����E��r6�Ĵ�c�����cl�ש4-�S�,�jP��_��`��T/�v��q���ܺ����7�ЙMv�����h�#@���u�̟�ir�"J�Q�@��\0 @���Y�)�иC���v�+e6m�`���I��f){@wq�@�w��p7[#��衰��hZ���)]��N�L!_�boQ��N��eB��zC�4F6r�P�ԋ2����2w�jPT?U�!B��Vc@��.���T�@�>��A��*TJ�B�q�� ;�W�_�\~�t�`�6i�/A�yH�7Q�ܰ��fs/�*q@W�m���Ф�JWJ��u(0>��z�ҳ�^�u���N�0:�v� l��-QT���V�-�VG-���*]�$K��46��#Y�QL�ԛYz=��#�U�E���6�P�^c!J�Z��
�Mi7+*�!5��KG���3DCգ}x4�r��A���c��[���ᡜ���TN�ϳl�V�x�Ay�
^�y��WJ��P�#T�:���fʈ�G�mh?%���)�jo,��Q+=��]�3��0��Z�=�qVF����2���-��9b&?���N��=c�s�@�èe֊HzvȪn)gy����3��?|%�~�J.�O�p���4���dq�Mʜ��8��T��ZК&��J��q�JU�ƶe#�Ң׵�`;��֚6]��t��}�?y*{�O��?c�p�U�"�`:Iɤ&S�+�o��.�-�b�S��_&�����l؏N$��,qWA���e{3�O����b����ۤ�����V���;�p�(�h-���U�Ro�>A�ȑ:���t� 4ё�FE�F%߫���촞����y���k�����"�{y���׌��E;���q�c�����(��m� ��ڠ�|�ePn���Y-�ltGewޯ�vvՖ@}�xW�(�R��Zl��Fv&S�*�ڛ/�&�n�G0З��DQq����-<��5��i�7ưa�Dj=�$!z��'�G'r~z������۬H����z�u��;��7��k}�m�<��bT��U^�P٭`��eY�cP�Y�|�5�'�!f9��kؗi��O�>�P%�jrh���׿�6DpP�1�#�2�l*�1`IRʶ�3�3iI$A��t ;�@_Q���p�R�#(�fwL%���]+�s ��L�a��O�/��r|xL�K
V��׷�wxwwM�iԐC�tYr�{`�\��=wr�3�><�9�`������ײ?S�χ$�������䧟�*���'�5P�T��1�*�7������+��
eL��s��� �.DR>��[���s�5�N��TF�[�>�@������Lg�d���`�um�;G
�N�����{R���6�1Ԙ��ӄ1m��H�v�m�jm�%?3�S8��;9��/Z9^R�mVMeV!��K��|T�D�ۻw�n�^�./���]h�co�ز�E���%x%��P�sS��T1�,�&�NEu�H�UdI�GF���`Tᖽ��4�@A�􃃡�=�,~)�:��J�(���r�X��x� �
<�u~1�uf��<{�T^�|)_~��<~t&�e��DTuGU�p�u�E�Ν�H��4N�����nP��J�
�_R���5���I%j��9��y�>���[lNnä�H�	v�Q������^�â����Y��T'ѣ`$C"�)!�����`�(�0B0Fcl�y���� k&G�57��+�QXj�d>�MPV:�- ^�aX**N%O�V*���@7���t ҠR��^Pdk�Q���(�h�z��h5�Rl�k�I�z���CU��@�QfPd��E2�a� ��@��~�1�����6�XXi��V���RG&`S�^��2�·��r��o���b?��$���됦[6��%%SEG6Y�d��RO�u4�K��������l`��B/��:R��)j�:��ҟ�?�T,q4��>��l���AyS�/Huݪ~4�Do]�^
7�Ն�RcCe�X��ݧ,28��v����ĽbV,���2�5 ���uE�7��hIO�`8��O?m
�+{X�|�B�����WK�� �F<w���"�!���6ۙf;���H����o�)�|�L�d���w������������$���F�6G��|߰����5k��j�*&)S�s]2q�ɓö��SJ^C��7xPeC[2������{[_�	������.q\pox-��A+�d������S�]�ʞ������.p�����yR�TՍ��� u�B�ף�/����PG�̠��BE�7�vGr����$�[fG1}��7�a���WNխ����5�d� *��b�}Wp�h��H��@�Jo#���b�nY�T{!�`��c�����M��N*A�lMq�d�S����^�`y��w�f��ѳ��.C�"������.�X��c�V���T�t�T1�	��R�?i�;=����N�S�x뼇� �{&��@BbJ��N�ތ٘N��s�̧	[Y���X���,�1�X�� ��d�֛�f��\q?we�U�vmD� q�XS&�Vt~&g�dBc�c��w�)�����]��h��J`�0Z�LH��?���&j�N�� �Y�m����h5s�h�1Zy��/j�h�
Y�X�:���U�f�"���~�|���L����F=F���V�0Z�T�R�V�����Y�X�~�A�XP�Lԋ���3�A�,_���*om�M���L�fP-�:::"���~>�Z��w��q�p��d�=v��(��[�����{f�p|�,AJRa
�~��'����k��W^{���s�Q��n�5���Pz��Y�M	���,�>@��`�ŧz7����T�j������8?;��O�P��4�Y%:�.��	���;�K"���M��g�����Vk�k'NiC��E���oާi�����#i`��&�I��)��j�J���o�{�'�
�U�t�VV����AUz0�gL��l��O�Y|{t�_�D)���l7�9� �qss��խ��j�ZCՁ2!c�i&V��5�!eOU�PC!G<X�*ڜ�4��:��*��mgA��Pݠ�	4��mkq%��[.4iKs?Ee�+r����ف����yU\���
��)��x`��P��fc��!������(�;�[���I����B2ǌ�&�����ى�;�@�*��p{Y��F'�}A=��6�`N���2/vj[��o���|�s��?��\�ա�]O�W�A%^����91e��B��D�������k9��FCϠ�))\{�,v�;�ܯEC ��Ё���m�������kw�p0��^�ofc<�(}�L�aT�8�L�Q�/�D[El("��G'�O�|����dg$���|ȁ������)\��U�QP'kT���);z�r���9�M�j�5�Y5Wg/��`-�I���uJ3k��f����tg�6�F�
�k���K#���9�����yv��9�K
l�ZY�{�������m����u�{+�O�f���uu���Z�ӆ�2�B���!���>jD���N��rsQ��(coN��*Ik��,�Xb�;㻨�`]�ì�8ݬ2 ��?���(�@@uD��ndBY��m4:��Q3�>�y��2�F�8��fe~Be��F򄴞9T�V
Q����4�{���{�	<G��`�U�Ӧ40w(�])Sp�F%p�bShO�Bh����,ԃe��yF	_P ��]�=ڣd�Gc?���݊�.�#ъS�K<;��9�)+}�a-����j#i ��P@ 
TE�lYkX�1��	�-��K�6���Ď�k:ːfW��v��xĞ�J �f�{�x�^�d{���{��z��H���ɤ��iC� 
��%ڽPaV� p��U���(���gg�����Ԭ�Z��p@MzWT!K�C47^�k��$9?9�_�?��V�o?�������?������k��0��k�����#檫�����cJ��h���Kä�֖�-�n(���yp~|`6��'��5�g,1�'yd6���\���zhYh��3%����n���rŚh^kޛ^8��|��ϡ���[C*�ʯ�W��pL�澿��7kY�� �da ba{��c���\�"8sz�alJ#I��	,*=�l6�"�UQ-��1�^o���V-�5�
�i�,B���I���mb*Ί�7�>&űqH{T.S���%x��a %ɲ}>�ೣe��q�H�E������SK�� ��7(����k�'4s�x|��rr�7���`m���J�Y�d�f��f��ŽRx�g�:6�M�����RrDR����QXb�Ԣ�*13N�tzaD�) �daS�#�7ic׺^p�v%^�.I�.�����Zg���#�Wx=+���"�Q��
�\�A�D�U)��zbk��5x�A�0>4]�J��h�oZ>7�B�l��8\A���#5�H�!���y�=�H��������0��B
�p��=h���O��M�s�d���k�.��W��tP���oG,�sڛ[�Ŭ�H_����"_A���a]��*�,�v�6�݀�b���% n#ҙ[C���f�geuClG�릭�]��]Qx-C��������n�R�ǰ�_ �Иp9{]mx`d��P}�4�h��yrq.�{�B��ۯ�œS�Ͷ`~w%���,޿��5aYv�S	����l��#m�r�WU� ֕N��6�'n��p��v�杔� ���.�kF�>n�Ё�]���έ�<�@�#�3�^��ԭ��<x���z�Pֳ�%�PZU��,��fΨ�e1�o�)`e���ܚ9Р4{jq�|R3h=m:�㿔�v)��R�({�k�=��G�Z)B�*�� mT�����ʂ����o�+�(�H��N�K�j�_�"�b7�3*�,1X���x�1͸�j���y�ѳ��u1SkY�(}	����1_���Q4�{�q4E���aW��Z(mk02ѕ�:� +�|�44X_��k�����;g'��ڤ�q.Z+��:)z}�	Y�����<B��5��h?TXh�2�hw��S��Ũ�A�1u�;zFP�X0ͤ�*�_�������5_���,V���Y-���Jm�i�͍P-���E���/)�其�|?�:���S����~���o���w98�(��J�h��r{G̠�B�|���+y��_���v���YZ���?�1��f+Q�:�/���`Jٯ���o���T���)�3�Vm�#��dK�S�},�C|��S��[�.�pdr1?��8�2�����ފ3�x @�RU_��r}s->~�	��A��˥t�E�]�;=x��0�����+�!�<L�}�l�z�A��**�Q�� ��W¶>�w�8��d�A���E*�)(AV4JOUXU�H���NB�J���(-(�wQ��u��U4[��H�h;:RWGU����hA���.2�U~ɩ?����GC�AD��0ux�u~~-(�>��`v��L�'���Za�O%Ջ�T�q�lci��M��c�X��ѩ\\�����x����c���"�K����Pq�֬�
L��o5,&��96�k��QƬ���)�eL����:X��@~V��� �������Κ�.��C�FP����#���N��F�:/���{6M��˛�;�.u|��>�&b՝�V@�d��(�^���/C�^�2J ��N�^'fpY+fx��`V���Y���z�����3�t��6�X�_w[��� ����g���O[�
zU�:�������3�M���\�&zmc�Q$ȹǘ�w,�0�j\�{ ftP��h��hb�A<֤��6�j5�+�S�W�lv�"�v�-h;S��o>��yS�+��6ж@;cf����#��Nk6:i���y��B���ˏo�<ۂvy+�~y'W����ջ<.��n8ޕ���vF �[�ƫ]R:X��� ީ�}�@��풮!o�R4���X�R�8.<�fwF[1�N���"�� �G{��̄�+�1�E��]�,�sm�� �� ;	O3U}�2D���dk��Ӹa��:Ef�p,��2	%��R ��~&�]R 4Uk���2:b�;�BTB]v�9z &$ԃ�Iק�e��&5��h�����*L���%��syvm��(��8)��z�hA�FU�އ��͹fƅ� 10pD�PU��
:� W'ӄ(̕S �]5��]�A��g��ܜ�ʐ��ذ}~��2�[�j��w���{�gX�"3p��>!?�9E�v�O�	 pA�v���2ޅ��������d�%��'�ڭk�ҽ�2����e�o�	Ϸ1�%�4v�&
<��Og�]A\�Ae���^}�­}�5�#��ʨ����|�q��w�M�q>0	�!yc2��0��=��=�oQ{Vӟ=A6��D�?~$��F~�ҟ��]���&�d��6߇���YLdp  Ӈ��v�G��(���u�u���_(�&��)�K$O�4	�^����7���2M��=BR���Z{����~�S��8��),�y*� �X�`L!����%��)���M��Mw�
� ������r�p/�?���c
Pa>�����;[�}�Ť�=�Y`5(�0����=Yu24R{uD����``LTP�7���q���?š�tS���_��a)�9qƍG%�WW��{�^�!;Q��츬�U�Qx���|�x�����2����! !�i�LL��%�.Ȕ�� �U�읿�I��e�+���GCj`�PΡs���J�6�dfl=�����5$)��OM�`��ˠ�7�h�L~�dw�d��SE����`�&+�{5�[��_L���z���q"x)��e<ųgDU�/Ƒ�Ѓ��Iݴ���AY��*#�d�7Ԑj���M���-x�9(�?7�%zSA�Fl�Xj[��TH�G�ـ�*5,�|�wg�y�]�����2{
yn�Z|m����i�� ޿���xp�6j�Y���OW��BW�\t��m�)��2���i&7~�T���v��D�W�M�)�����D̩5͎-�ˍ�	�8�%�<8+����}���/��=�R�#��-RPT6&/*�Z���X�O驤j�1��?=��� ��fc��m���[Ѐ����l�Y�U�.��3*f֦͐ndc#��6%�.6�ƶ3��-dH%6G��G���!J1�`��Т�6�/v��/.�_�})���+y�4�ky����������f���;"��2Y�6�|�����X�t���;V*�P3�`�6��lV�/�UFVgk� I�PvE�q���F0�!�4��fm�U�{���X�I�qZp��ԮU�"u*TE8�hU�Ђ�.;��(*��W�[&j Ņi�:��&
�p��=����y�(�sP��*�)�=�S���kR#s���^hp'��#:���m���Z���~�v�7��ߩ�gʚD�G&Ů�d4��5�8T�kE@��<z3�X7 T�Qp�Zb����R��Ip8ۛXܵ��I1��V㢵G�w�$�y/+o#�4g�6�ڵ�ǉ]	�ض �Y��`J_�֬���j�x��m(p/���~~����ꨡ�I��ix_�1�G*{��u�6���H���rm2��0�G���� ��"H\��U�
8��(t �����Q���i�v-��o�f_�~#�g%(�:������1��Z�N9�iC�4�m��l�kf�cr��`���Wryy#��޽鈠)S��PVq,��/��/�ɳ'����#���ruy������p��G uA��?����{�Q������{	�1�����^B<+j_6���%s
�h��u�3�<����x��Ko�m�{�AYS{�*+��ie�O�^e�8CD�����s��)(��Fc:0��8�%���l����z-<��YHQ�sq�}azФ̉h����t�
��=Xb�fB^~��߁�-�^ 
?N������ �3ק�ǃt�;�����
�d��9��t,��#����j�/~�o ]#��|-O�\�0E��>|d:�훷Lyà��\�]���.;B�GT�;9D�}��P�T�.I�Ft�~N���;��σhNe�
Gy>�P���0��G}\��J����<Њ}&�7M�ȥ��2�$�q!ݎ�Z�HVZR�*��M����Ni�z zw��L�O�j�Eɡ�2_Ȝ�j��t�8�YQa��a1o&݈��ǜ���3���Z9��}K�`UOe�p�״��.�V �z��-��!�GZ�a� ���>
�gM&�Iq�5|���@��퓼)�>Y�YzWU��T��X���Z��$�P��V?Q�'�V1�b�jj�_5��`�3u �&��v<E����ze���S�r[�:���<���]�Sv>�S�GG�������|<�2x���)H� u_�i�'�)�)��j3N��f��1Q4+lf���~E�4S���;"��_�X+j����}l�)j�FU�K���X�:
�+U���!Eu�1Y�;�޾@c�S���X^�-��B���%����5���}��˧�Ͽ{./�^�4����O�>?޽���[Z�[��)c�6��5��Ɋ� &��T�l��dw�Z����t$�%�b�t[��l�
�}���ʢz�����;�.`�72�����bI�y@�6"(Cn")L�gh���u��#lqR�V��e:U��h�y�KH��/���*g>�*@fW�X��5�@k���u�й��	0���(޵P��Y)H�w�ٕ�0V�B��Ck���Y�:X�:�P�MB$S��zM�'±�����b�s<��6�Lο΋��:$�j�r1�DUQ�2&�%��_�=I���iεR�C�2ڤ�Q�cÌ ~�,ԏb�P	�QS�CL�{�iM2	�Y����#��� �6�~Xn�ܮ�(�������T@���6Q[�De�}��Ii�LHU�b�:��R��sJ��Ң�Z�`�����4J�󇥼~�N���9>h�`���X��xxx"{{��7�*��%N��3�mp�������	����\����=3Y }�OVb:jٗ��8�b���|��sf���(4���i��7o�˟����������Q.��e�"X�Pk����*C[��bF`��3�����<��=�e���%~w��z��jU��t��h˿�7���y��"b���Ԃ����"���@0<�*�.k���y`�M��h�'˭�� ���9�kJȖ�^��r��|���zy��ڞBY��f�aB~;ȲA����
����O��ޛ�f^���������@O�v�M�·^Si����)Vl�����~��
#�j!�{}r�'o^��	TL����s�õg�
+<+���h�wU	��@�O�Y��F��W&����Q�2���>F��ep�r�lA%�z�%��	��BG6jC�h6�g8UI5�L�E'���.�	w�����z����7F���hJSWEݩ8�0��X0 �q�,��eݽ �WG9�Z�iX!@1��y��<wת�膵i���u�{��tTV��٪�Z3n��s�N�T�7���E4�C�kgC��8@��SAN�V^Q����k�qd�R.i���$ee~��D>{�ϣ~ѳ��PJ:m�`M��,�tpp�`�:?�RS� 'h�Y�)�F`���B�T���J	ߒ�{�d7%ま���{Y��Ab�:4�0C���
r$��U,��'���������"mM�%o��A6�nao�N��G[��ʨ����dE`Q�Mg�ɚe׵!�Q�8�u�i��U6��f9h#��rtD<��N��̈�P`-�;jh��~��|��y��\��Jn/����{���F֋;�a@�f�渉����'� ���Rg�$I�#ɍ�(����ۨ$J_�K\E�K����M��f)�5F-�^'��_e��Cd+0Q�gl3�|k�a�p�G#uv�D}O5�F�UY�y۝�Y1��Yf�D�J׻�[���!�̝.��b�mE4J��h5hU@)�F��jo�Oz���y�<d��UAЎC�2��Z��ӡ �u�m�+�Sz�'Zt c�6F�Kb�V�kY��q�34k�a�E�7�̪�G^�E�nNm�d��zq�T�wܻqM�7ɞ=����B��H؞�b.�Ń�AvKmچ�^˼Ů�U!�!p�{������~W���>�0�H�^cM���TEg��"TT���f+E����Sd��P��թ����J� �b���vVI۷P̯ڪQ�	�n�����Ǉ���\<�0�>���&=�fg�w��r�IU�5��	��@�ŵ{?9�ȳ__�2��6�T�&t��Y(cua��'���'/�?�=�,J.�� ���ݥ<~�XN�N�~���Y^g�%0l�½#覀����o��GA|���g�����?�9j�R�(�K�r�� +yǩ���O~�c�48_)����z�4C6.n
�Ok򔙄�tB�n!�Z.]b]ǹ����ZR��Tf��{g$�ϥ�����A�yKMYrq!k�m5ȚdR!�ߦ����B��@[�t�����6��hh�9y�%��We��9�����j�5���F���Z޽�`aGN�Ȟ\�4X'���`��\��ШJ�����s�,�!��L��~��EL[���__�跪O����$_��`����J�؍�e��~AJ��~�mD��8�sYkN�fT�I�S���p�pB���F�4�U��u�bd��O���p��R�2a�����M�m����ژ���.�Rwv�co�hT7��GFJ�[�(!���Z�`���h�8f��{�������௵�G��P�}����k�+:��%r��n뢆�3�}*A2[d�v������Hd`�ʜii�g`��7r4@�(�'}ts�{:uvcۙ!������5��W]��4��|TV��Oz�$����飪>�S~N��P"�-��/�s���F���=�ר*��$�5�ץTPT��x�9���{A!GtAYp��H�0�j��D�Pt��t��Sm�SWל,P筎v��~6Cl0ڂ�)m[aNV��V0�iІ��/3F�9;�|'G�`��W����G'hy-޾����jyG�.Z8��&2k�1��ͤ��h߫F��֠\�}��� GD,-��{�R@cc��Z�,��h`V����@a"���77��ǵ/�ѿ����`���2��C�u���R�am�֗�����A�T�'�<�|k��}ù��gQ��w BY?����ն'��^�iRO��z0eZ��  Sim�$�����@m�v!�&��-[���j�k�1ú��l����;�F�/P��P���% ��&��g�(ثN{|�Y�'b�k"���h>�.��;��fS����h#���l_�C^��b��fmG�?#;��`���|��@k�Jf�UJ��� G�c�v���u�@0�@���M��f<o�`%j?���Z�KE�}� ��*� �d�Eb6�bP��T�?�0�hL"IF�R���r(U��_%;l;�s�>	|(�I��Ù������#9:�ev�6}���h���o��D�O���j���<�u�7+ ��?��(��yyy-g�9`;��f�kE�;F���$�hw����-e�qz~.g�����#�)X'�����?��|��_���VEΠ�iP\�QW���:	�q���}��?/_��|�1(3�k�|�h��`���Z-�����ݲo��u��*�[�x}_c�ϜS�R�ݗ��5�h�F&t�qR(:0mv"��ִAY���w��Yk���E�O�R������.:���!C�|�1�|�l���I%��*�!K�P�AR�&R1�{s>Hkb�ϔ}7�]�����W9��xuI�M�vc�Ǌ � ��&��� �^���e޵�SzN�|�ygz���|���.�|�b�*?�ʇ#����% ���i�T�J�;o_�b��R֕8��� �d1K���3�dd��e�q�t��m��8�1^� ��LC(bΛ;���E��:d�]҄BZ0���ew���l<�2c		���l@2R� �s4�R�j���k̀���\3����%���&E���f�8�D�2��ӻl��E���ۅ��j���;i�i#�)ƲŐ�^u'��R���?�k˩��׽Bf�i���MP�;b0>�1�b#Nu�L��U��@ "�2��:W��p��&����gl����^�B�
n�ń]�Hq��![���F�����`��^|���V��$��U?Ӄ(�6�*�0c��tj3"AU������oI\Ҟ���>g�I:V%ހ\�k^쀃' I6�ύ�@3���}��҃2��:fQu�ƾ@���tn�������ؠ�&�j��P�����l0����۷�p�1_��NN��\g�5�, �Q3�Z�'��5��5.;��=�(2#-B����������\���I�&�/�mUdɏm�ã)�6+��p���=�7G����A�/�'���Ak�^��ؑ�a@��o6ىHZ���JkZ6T�ݰ�
T�`@��T�c��,9wa;�����<�#7 *�	���6�KM��K�J'0j��\�آw��R׵�r����r���@Rz���!X�gĶ�hc*w�TP�؂����z��=�3�uǄ���TD��_�cj���ϑ0�9
�5@�*w��Kt4��<�B�î��l
��f7�*y��'Kc�����{�:��˹
�C����*[Y����ze�u�at�X[����T�ZP�ŌY^�Ph���SQ		���F�S=m���m��S����u������S��g8�����m��@��N$���q�K�n�5�K*R��D��H#Y��F+��i˵�4�`b;�V;�T���6<�7o姟~���/d�?U��sF���U(�7��.�:�6
`u|�������T^��R���|�������1��f���덍O }Z���ҥ�bU%Ъ̆:�!�<�l�Tɛ6���T����EQ�S����̍���T<�ʅֆY�>H����
=x_�Ϫ�>�h�jo�SY�zgS��h-��A�<	ډ�*�*|vm!�8���Hy`�]֦����~��r����/��7ا�q���`e��G[�+1ʈ�� �b�'Q�k��=�z��'Ϟ�����r0�e�����>\���h.�o);�]C���]���T��u��e ����n�k�_+4ƍ\�x-�|AgX�i(\|Q�/jHk59���şQ��ԛ�9���4�S�����~�c��eY��F->�������y�Rz^@�()E/Xa���4�8C�a�;���A6�~���2���.�?m�'&� tq�7���B�yX��Zr"����١�d؛��f���R�i�ȟP���BT�T��cOvTJ�Ž��>�@R���4W3Q�ʇ�]E�0��ƮX#�;�0j�Ӆ�?f��D��իͽ�V�y�Bf�;T���k�� �ǲ{����� v@�Z�n ��/����RB�B%�W#��F��/us���\��������}���<�h%ڡ�y>D~lX`�&�x�(wwT�Ծ'-�~E�|]�������8�X�Y�������-���"UB�D�P|L�K/߉ڜ1T��E�.���D3�I|��*&GȔ5BIy
k�ڳ�!���.l���xf��G���t�`t��auۭ�+�����Ɵ+�R��
k�1�U4�F-#�x85���Z?��0�тp�®@��\Ds�H�1T]�\�X�c�%�5{�*S )���(�b��k˲'�3�D]�U�@k
Q��������ON���yt���v.W���������V�f�5�`D�,Ԥʒ�:�|G��|+�l5�6������l�����j�]K��I��Nw\�G�u��˞J�� �����I��a
DEQ�XJ%N�	��oQ�ʀ�O��_�*��}}��}�4 g��<v/jn��4z�;��۳�\��?@[��Ӂ�7���I�Z-�Z���\7�,6���ꕉ(l��1vJs�#�"���
Q�7�]��Bm�K�|�O`(z �^���9쑠�#[ p��@��j�����A��\/�u��e�z��o��g�����U|�B�h���ihs���i��R(��2B�V�e��x
�0t�U"����Ƃ
�΅W�h� 
���G�%8&
y`/��*`V][s�1_�����wS�Dٕ�Î,�>����~�kK4$^� �����J��"><��Tgң[UD6GM����h��� ��{x���K�̠a/��e^C�B!c*��km�0�G��i��iݍ��Y=h�`���8���֋�:�y�O��`;6*�ס%���Z��{j�geʌ�c ������,{@;F[�܅����2*��'u�wJ���Sf����,])EX���ٰ����s�Z��s�V���ѩ�� ��@�
��+�|�t���Ze�4ܟl�a-�9���ys�J���凷�e�T������W{����+T�k �R�3�?Q��7�5y��]�L���V��)r�����ӁJ�S��&B:����9��mʍ#*�5�vC����ߨ��R�8�;��Eʐ�7R�Y��D��%�R�hLEN$g�c��D�7���WX�gk�
Ui�RZU3��ң;Q#٥A���ifS:{�v�6)�L�������+����O���_�&2�Ytj �V�M��ȿj�������/^����7���R��H���>���C��ǟ���A�* �7�`��&�O�<���Z�=���6g�*u26R����c���P����fK9MC��˷��/��ɸ��ʣa��g�"J�@��%a��*-��lB��5e@��bB�M�,N�R�����`cZ��ƜT�5�r^H۰.ʅ�"F��Q�6\�l"�@V�9�������d�h)cI�:��*h\���!Q*ʑz&�sz������l�
q4S���V��3F`c!#kD� �ꆔw�ڞ�S��d>�0DK
�L���-�gxo��"�Bjs�d@��h�K�߸��G��1�S��-�,�㡀'���s�Mxﴮ�b al�VR#�LJl.���l!_e���vk�|-��`�Zֆ�� ����lnz�f�(�&�$�J}�G�1N�G�t�,&��#������F���:gRh�Zt����:}�����
�1~2rn�>��ɞ�̙S�4 gH��R��`TA%�x�����g������{������_���-���NS�Qa\7$�kx�KX7E�AEg�������*f��ܪ�W����MԈr�y�(:J��"�]�Z@sb�%��D�c� i�U_�b�h��O��o���{_�����c�o���$H*�ˋ�k��aoY�	m"?��B
e��gR�͛=3b���Z7}P/b��Ƞ�N���)��ք�t����Qe��%F	�T]ꎆ�u	qW�f���{y^tJ�4,�2=��m�����dBy=�
{X��|iJ��S��L�C6GP�!�{�eZ�]���9���5a�O�&�����r�R�V�&�	S�^��*<��� _я��z�V��v����+f#�F���Xeu&h)hV2/`|t�C�`b�M����E�?��E��;*�5�Q�����'���S���2�uH�Ba�0�gm��Uڢ"�&�+Tw�a��рm�าl`3Rڡ�Һ��C�X<��V�����#y��	���N�ү됵�짧���z�{�}�HI�#ZZB�(3A�<��w�R���c����z/���+���˼?쫸PrV��^�N�jAv�NF�V;Oq�J3������3���/e�B}�:�q\��ή'4 � +�[1cP h� ���^5H�����?�<����/w�$�R���/{s���b�x�,�+���]��}�UU�vA7�{C_ܕ��5�<Y%�<�ge�2kb�M+�����L��$D� ֚�����>�Jv\�	�E������V��N���X�7��e,l	�h��aP���f�i�J����:���~vf�<y,_��<}�7���T����8/���_�ʻw���#�0�T9`�P6�w_%���˳gO�4�FM	�0d4��=LR���i�_t�fʄ)�k�{�6p�u��/�B8t���l���(|���hCBJa"����tR�^�9CxZ��6z7 m���I۱�,È@��ݝ=��=��������$��E�Y���m�H�]�}���ޗ{���j�J�L���!���23^� 2�͑����d�4 pp0�Oo=��h���̲���S*S�JM,��r��H���`%C�p��z�����_6E�^k^�06F+�A�JF�z7C#���Z++S@��PW��ߨ��06��������p��wJ�Jg�E	�-��n�$��
�䷗�l�^�$�uM��h��a�恀�n��Y����.7Tt�c�����wJtAհ�"9�� ȕ	�������^�^���<������[�F�0���d���p�}Z�D�9���fGk˼�iB������s
���A��F�Y��u9��m;�g�OU���I?m!�f���6��F:e���i�rϴi�����LA.������U��&��)���Ճܤ�o�|�!Ԛ�y�,�e6�����U�4��:X��0n�P�y��av	���`��Ÿ�3;=d�@�	�2�U+Y���C��ބ�z��l٫�Ի�������zK��%&�~m��/w��������x���m&C�k][��	�h�������ۢ�����^rA��Z�R�7���}:�U��Ppߘ����hc|�׈�YF貅
[P�3�O�ô�u��F��!��*�������O���m8+i���]O� � 
� جa��ժ�&?T�0�]B��e��*�	J]��1х��J��1[\��	-��_���������0��{��6�_��b�}���M�6lҵ�^���`���}���0V:8׾:���C� j�*�)���ڳ�YRx�,�,�)0�Z�7]�u5�➪��l����ANHZ�~�U	���9P��	sW��������������l��Q�j�[V�j�����R̗���F�??��|�,B`�{�=C�;�
����dB�@m�&�Z��P�-�-��׾�y+����.�.}�F�&2_Lò=!D�>����h &�E��D����:����}���o9�ko:�?}��\^A�Xe�3U�0�O[�r���v%�����ښ"�W�Z.�����m͒��X�F7K��E�4`�Q<;v[�ߪ��W���Q�:Z�M�n��'�n#m3a�QfE��7#ScC�I��Н���`̔H����C�/�軵
�l�W+��.���B>�{̘����Z�[��-�-W�F�b(,2�fNOOd:Ջ='?��g���o��~x+���y���;>��߼�J �7߾���y���eP��'�p�|%wۭؿ�£+�;t7���g����ox��c���;�x� �T�� �&�prV���6;(4�*>?��qh������ ��Ʈ��� p�t��b����a[ Y����7�t����)�x�r�
�8{S�ц�&�����	䁿*){��y͠����� mc}v�ͬ��'"�
��μr��=yܱ{���!3p���2(P�����KG`��ls����c�D�M�\���V�,�s���>��s+[��Ҭ�ӿ!5�$�%�V�4X]Ov��Cĕ@p5N�<s8��Pd*���#G�+/�ć���['9��/�|��y��=O�(�Y�܀�כ���T�,�P3��U+���XƳ �?�q �{rr"_}���~�l
UNG� �U�}��fm�z���81�e�b&��Ǿ����nG��wj:kJ�8p �Q�	�
�`_uZ�B�j��*�B@����e:���V�wk|��Z�qtp�s^,�L�ړ&���5��T�a�@�&��B�����=A�>���^E�H�,�{�XR װ59|ۓYq�.�H���x4Jg�U��3d��7��:?��\�`٪�{�Wi�8{�����A�Ҟ��<�m�G0	0M�w���uhi����U�Y[�,��2R�A{��n��'6������iV���:DgoX������)�Z~Z��� ����ZA���ÏK��� �06��/Hv��kEfPlӣ��t��H���:dXiEم�FU*���)�=��_�����V�Bg2ծX�Z��.�pL�� ���M�J��tf@b���3�����g��:j#�H��<<$[�$a�{�2��-�&*$7��8�r���{�v���V ѩ�G�7�����������i�`m#1�Yl�_�*����h	/Ӂ;���)m.�U���Ypk����h��ȱC8�g�G���V.������h"�hP]խ��3�߼����y�����D)Z�e4���W5P
o�V����6�9Y��Z��b�``$+o�����Zno���"�n3�&�XB�������n��sp�H�5�ף#��C�ýقU�� ���LB��j���Ez�ƒ��V� )t(#�l�2D�ݽhתyҴ��^-��8��Ny�[��F!9����KLx>Փ����~��{Mh�
��XS�B�)m�$A]��9���}mw��U$�D�8.v�YB��Vז�oz��T�*����RV?t� ����8�A������@ ÍW!�:��S 0��l����������\^m_���I
���y}s�ޢg	��y�Bޤ���d&i�i���ĕ��[֏�[��ˉ
��' PW_�;�-t˿Y4u��_B3M�i��(�ؐ1fV���B��9���iḡ��YQ�W�A%�����5��z��9gLM�ɐj�e��r���m
���f�J�p�ʐ��G��� T��S����Y����ld�#�
Ƕ.�N��쀎ږ ��C�~k�����fzHHP.��X+�EAVC���8��H�����8Z�7t�P���7O�v뽏�� �UAIι���&���I���>�k��V]��A�����cL�h�(���5�	��!W�7�1�� ����l�� �%�K4�}k>ц{p�x_/;|��;1].lPb��oF�R�Д]C.3�A�ۦ�zC�
���4�Ξ'���*�\P�� evE���
���ܛi��2w��ټ#40�#
�u�`	l����<��[���k�P���h��ؤ}2J�2���Y
v#g��==�^����_�������E� >����&ʍ�<`}�|��ʞl#�"��dv�UjP����_����>�h�5Mp�egQ�n��2s���#@R࿺�X�&�����@��@�m۷����/EY��罻��|���_�Եk���ZT�����NA��qH���	��O�i�0;]��*�Ǵ���Ԯr�c�q5���ou��4{M__k�v����^y�� ݫ����ņ ��
V��cB��O��uׇA�X�A5��7)�߶��W��blZe
h��$�՗�XAݦ��
	$X0�r�j���=��.��H�m�P-��]�e��ؖ�?q^{	�����%b����9��oE�jK�c),ɓ�Z'�n-C��܀��։p��(�K+h�����㼳� @º �C09Mq�Ȅ��E���k6ߗE�_ϓ����g���/ .���r���r0@�ȩy�����NkU� �]2��~���ː� X�j�U���4��k\لu�@���I�h�5�qo� �L^�<c���Q�*�@�����1{h�����i�6�Rv�W�ZV��	d=P@����- �=\�ǎ\]ߧx4���C�/���|�����U
s�*f��4����|����*(ۗ�M�� ��0�N��r~q#>|���X˩�C�s��`�A�E;�b�Ĝ�C�D����k�]ͤ��R�s0��`�v?5v����Ox�+������񖅴�k��v�ǀ�ۼ�e.Ddw�ћMs`C���{	��*��Y�
Q��;6,��K�w4�S^Uf2�W���u�r#X��4�\��g'����y�/"�>JV�_x�Yb�:k%30��V���)�Y���,�#HH�կ��ϨC��Y��`��Xh���U�a��^���������߿P9EP<[�����~F��JVQ�RKe}ː���T0*��^��E�áS���u2Py��P����0[���4tm8ǤvT���yz�X�]��a�CP;���| L��ɡ�[����2A� jr����[4���G�{L��R�����K`��e���%A���0h̒SnC)!��%`�<]�J�)�%e����717���+Z��-��IS�$+�=(��A��M�
��@uO �j��ú5`u��fz��������K�$�f��eo3�bM�5�����q��P���`�~�!���5P�%�<{�1[����4��.����"�n��cӓy�6�}��)>Q��+�X@D���q�+f�1� ��`��&�95��f���{��뮰$H[tU�n+VtT�Vj(e��:*�`������T�*�j5+0�],0�{�i�����Lx<;}&o^}%�NNe<?f�5�,�KS�*��b��h8�`�S�`c@+N{�Yڳ�^�^|��?|'�/�Y�ޤ`�44�c�Bи������$�H���܊e�_T�X+��A����7*����$ �+'��{�/�jje�M)��g�52D�z洶`C~�`�|�������Q)Ю�T"�b�����ׁ��5֨�# t��0hm���������c� T�m-e
����G��{4!hR�6j��r�p���>���s�H�@G2��8f5-�;
B��rMB:z:��W6�9CtѦg�$���0зym��t�k��:pY{~5���4;�3C2=�Y�����ĝL����}(��j����]�
����sh��� ������Ǿ��"A"��H~�a%�//h�'�	�e����V��ҡ:5�F&�~���о�:�=F%��se�d��b�Ab(|�D�Y�׵��k/��қ���Ɔ(����Ÿ�j�w��ye��PZ�W@���EJc(C����jA�g�\q-0�*]���p����N�{���
�)ݚ��@Xcc�H�,\���:����cBR�~����	�.d���lq�y�KX��z��` H�ֵ�Mfr|�,ž2F���GJ�$	�0޳4d�x�����8���1e�6�bc��#�2@E`�l]��/ڣ��`��R����]��Ly"���kN��f�v���ȉ[�<�l�����v�	�ĜX�\J�.�>��=��sN������1m<�"AAV.��;�ג�"���.2�l����]Qm�0g;�  ��IDAT֬�q���gY��B��	QB�폠�+�������� @�E�)z��@��ဩz�0/�a���?�ի�����|���ΝhH�x�Fp�z��W�Ě�"�*� �|}Y1����t�7#�Z�=,���2��	�0��z�˨��(�ޱ���5N^��L������s�Fxf��	V��p�YU:�2�T@�,qS�����V*!��=��$����h��M���7���ȟ��A�L@f�.����* ¦�%8�)�Y6[�0�����/l�{�K�k"�2B�:���>�-��ł�E2��;{ܲ���+(��3 wiU�Dg	��ʻ���=*g\��Gv�n�� }G),�d�����9`�!˼��u�[�N2��,r�Zс��P�J���-*LzX�۝��S�z[&����li}��d�kf��X����=z�r�;ZE���(�Wa`��`A7�y�t�GX�r��.�H�h����CPP5{[ƣJf�����R�6a��l:��g����7	`����q`�2��{;��ŵ�����ll9�% Ҡ�j����s'��p����8o���|>�$��eA�fu�Wv$y^!O�=I�j�����v�������ԖU�U
f6�{���1Ir�kŜ,T�W���?�ס���R���t�r�g��\�@����J���	� ���8���6�P�Q��چ��H��#�J�G6��
{��X��[��F��v��Q�S/ei2���2�����PV�_E#��
?������|M����V��
e�}|
�Y����f�Y9 �p�Bڦ��
U���*ɶV��"Q��hR/��
+��87�-D����&�(�a�(���m��^r���-�%�\�U���.to���+�}�$_�TqM+�w���	�L�����J^�|-�7�i]h�@���g�����V�����Gc����R�sCl��|N���>t@5�A��I����*[1�l���N�EYB��}:�W� �EѺ��.Jოծk�Z/5�7:��9��u7U$�b������z�`w=�6j?'��r����R��,�N��Y�TM�RD�^�A�ko4�鞂5�`�,֜Av�����F&�%�~�W�C�
;�?��Cdy��>9>�ׯ^����k��MO�����Ϝ͸�lP��3sy�~��e�$D�����7���]�
x��S��Ws�Y��� .��Ο]qY�k80+��J���~أ;�-�-��}��,��QC�����mKѰcwQ:p�j�W��,�I���N\G��%���ز�-J����v~-���_��e�o.En�.��W8m&�*��F]�k�,6�Ã�P]jQ�?9�j�G# ��ff�ZY���x�G��� 7;�:�{��xj�� �{�w;�E��rY4��~��,$�Z�+�dUV�2�Zz��T�ʏ[��i����퍜_\0��7�]f,�9g�&@�oI�j�{�n��4
�	���cP�N�oUa���.��Q�k�U���#*��-xj�k~��=����@�x6<�emg:4��q8!�)�=�\aC��7�ږ����te� ���o�6�%o����W��_���9���.�1��5X`5kC@�Ȫ�Ȓ=��,��x�����:��@x���_Ԃ�
R]�h>� �&��@r�#�f�M6Ё�Y�����-��|wܻ���g@
*���{��4�m��6����I���d�6���������s(H�h3���D#��?E<Զ������%}-9幇!�dÂe�|�w��b��E0 �]'P�BU�cH�C�x:���T�Gr|8g2���H���k���W��8�*&�	i|�3��Ym�{!�h����Q
�L���a�s)��S����D.�9?|/�?�"7��L`b�>�5�2ЛS�wl��X`�gO�����������Wӡ� U�,4aa�M�=�*�kx'���<^�OU���]�wa�Qf!�� �ҵ�����+�"ڨ��u��ZU3�N�3�����#M��}B"ɃxS�|xXe9wo���{�
EU�
=�H%?bg��8�Eq�2�Ҙ�"�*bQ�+VJ�U3AR`�&���a��V�%��\��N6��o��	\�8~T $�u��(� NOA���4����Z��U;T:!�bb�Ym�}�Z1���68 �3Z%��W^�_�U�k�u���
�E���B��zݰ
�0"�v,�i߼y��h
�߽�Y>~�H��|~ /��������A����?���& -�혁:$���8���-���p�ڡ���P��T[��K�����=�o��BQx/�oYo[@�� ��mNP��S
)�c��ĝ��4��Y ��h7�-�5����c��1.m%��1���kO�I��Ym�Qy���_)ް���ّ�~��3O�����t��O��O�Q�n��|i��o��-?;�G�z�c�J����\a��h�[�G�_�<�k���0zߗ&T�E�Nh.G�j����T���K��=s��쒃�1)-�A���e�V����~C�l�S�:*��6
��$�8��>s��{S���^�S��:����N�-�|����b!��'�P�e��փB��y�<(5I.�Sz�����g�{�|"��!�*V��XX)Ua�@��T��т#x*s6��j`
ٿ;U)���P/Vz��J�">lq�d���:�r#��������5�o^����XG��99`��w� ��U�\��a���Rڒ6�nH�Z.+��,���K���������X�uo6
^
�`M0��݇	�qf�c֙m�R���,T�F��,��5�BUPe���k:s8V4ImE�T��`ǥ��U��ϫ�A�����L"(Md6[�d2O����<t�������q�	�+RY�AKP� }Oe�U5λ���������&j�3�ȵ�ȝ��Xy"���j�ٛf�9q�vIU2��E�* ��틠��
��9���n�0�G��l�U
�tfJS��{m@I�@𧊃��G�C_�D�_�z�c!�UX���=ӡݏh"9�`@�fc뢱�s��*��Ф���������a
n�YD���B%vI�`m�n��e�����d��1��j��3�3�"�����@��4q�����w�@}�%fs$G�7*e>ۣ0���$�z��u
^1K~z�,��q��8>�*b��I��je�"���3R�p 4[[�\�*�qpx*��\	��ȧ�L��4��A�>��4�4Ʋ��^^�x�>��^��l@Þ�;�N�7N{z���L���d�IELSs9����꞊U����df���=ˇ{�->��ûD�"�w7|�� im��Ҁ���=����ڒ
�rؔ�t�5��A7�U�^�*)�<�L�=�S�?S*��l@i��֨5��D¥)��I��zP�-�&d�-�#�'H_֨M�M�OQ�H(�5�?�:۔5+f��P��@���`���2��F��Q�*ad��ײ��9�T�,٬�>�4�_AE���Lz7��̊q�Oa/a�1�d�GI?	`�����9�7��>U�7#�3X"�͠��z��-��Go^Ŋz�1V�8�]���tA�v||*/^�b|�
����\YgYmVlF����m����� G��z��zpi���GKEn"�/m��-��a"�Q/���t.���}li{T��[E��~�
z�c�!��|q���CZO{2�
)t�>+p9?��=wUT��t6 �Ҩ�0�i�U���f}��7��_�*����Q�W���R����H��O�h���eO��e���t���d�Uڰ�����b�7��.�m�i?%@xŤ����ޒ�O.�s��ً%/��-aO�{�!�?�"�M�wE��{�I~�c����ˌ�(|/�N��\9��m�͐�&DB��+Pl,F��#A����o-��Zb`/��0������O�J���g��������;�%��M�����e7������^%f��8!z/��4Ry$�ʌ"�v�Pq�0��/�Q{�_V4�B��M���N(���s�`�,\�0#�A?A��sH�kE�=aE�	���~��?v����K�_{翳��}��_eX;�_2��Vy�������K)�e��>\Q�5d��` J�ʂ�fv�?�X7ɰc�ht�_�le#*ZY��P��k��ͨu��e'H٨���l�Pp�i�A�&���)[�M��V6T�%]p���4��e8
Z��e�l�XrR���}fc1�o�j��P�L0d���l�Ӭr���W0���kk͠�:v�jX^r�$��au�2v̩)=����� (߾b�.PVc c���2�.� � >�)x���/���rPa��\���q�V� r��Q�(u��tF���4�����&��ݥ�����LԂAs0EH{u�spPK��d��3ߜk(ee�i���t��|��IΟ��I(GGG��CՒ�o��l�(ݔ�F1��������%�U�?�z�� ��~ѐ��G��^�B��0���*K�	�����&8���ԬG��E��TD�BD�^8�APrP%���퍊��1g]&.���@zĉ�*l=�R=2�=Ҵ�4)�}��-*J��������=����e����ǻ���|��J�f*{똝&�4��u]�ؼ��
��聋��������c�����ʃyVWǄ�Z�,9��7r��\\�S�ll@�A���+Y%�uɵ�I#�a<��Mm��m�m1�t�ly���&4�88�	D�:��봘�S�d���|�`ŃtX��F�{�W�`����`2���2����xoC0��dW��?�bbLBޒr���1��&�{���� OnkK� 4!��׶a��*�H��13'Kq*.�n$xK�
����,:g�m6:�ͨ���v�U��`��L �����6ʪ�!@+���}1{&��]j�.� ��M�]�'���|(��cO`��(��|��� ]+��^�����/im]��	!�F��IW��`�* ��8�{�L���f���XX�*H�#. x~��h״0?H�o}� ^������ W��$�V%�?~<O@�LF'2O�6�=��{{�ɲ[
�l�$Ě®'�a��M�f$~A�/ӵ<H ��ׯ��������k��%S�'d���/���_H��6�ۖ:D��a����;����Xń���ɼMǋ���lУ���fت�%<I�I����z���б_��y�A�=���7C/h�kbw�dn��-���������E�Pn�V��D������G"	�A�ҽV��#W��w���n�@_W@����N��X(t�׻d��7��-�d�z��>舽���^>H{�n��:�>��իB�*��\�4��P�{�^� l��na�η�6EI�s���Q�2T^�>�0���L6����y6	pdo��a?%���=h���K�ǵ���bѨ�-3�6��t�΋h8�F�&yk�N}�7�ݱ���#Wiu_�mH��ap]��֣M���e1u�6���D���-EP:��qԀ!0���v���"9�v%7)�A_�����p�臊C�U�`C�EL�M�f�#���זr��ʎy
U2U&dVah�L��'�D5ۦ5<ܛucC!���I���0Zsh$��Iy�J׮�,�,�(�x�g 0̣3fէ)�@@ւ��/2���/7r�eqK�EE�h�Fl���A��*�L�P+-@+LV�p@Sٵ*}Wr*�ӟ�23	0�e����L�Vnu~��MR~�]��R�句\}:wV��6W�B��	�KdjA�SZ����Өj1\���o������ýH@k3����`̬3�*T�B�-L�BJ�I���`��5����h�Ii5j��y�Οg��\c�цX�>�A��QYq�u�a0��W�T�[��Bkj��-#��M6�ϋ�gr����. |�hv��a�}VX��7tW
EhU�kJP
P�J��*e�4Ke�� �D�%�g�!O���0�n��Y�
�e�#Q����p(��R��˫�����Kyqv��۰��e���'�d$�J:g��N��W�@��WP)J��' *]�לO�p0M�3]_T�'��� ��k�@����b'�e�A���I |
{ M���
�-�82�鉷��� m��<]�Iz�Jc���=�>���6��o8�F{.!����P%N�M�U:��}s+6�Ͳ�*���SP��T@Dձ��o?����~�ϟ~�%�X�~�A��=� $�RB9�6��V�Wi��cP��H�K��'�"������n($:������|#�'�rz�jl�\��y]�d'�
�k4{�u�y�H�ao@�c��c��e���q%��{�$�-U1�=��t̓j$K�AIv
[>�2 Iأ� �d$�����K�؀� ٛ�Q�~�H8��]J;G�!����EB
3 �k��འ�"�IX�X�ZXЯ�sJ�%CVD٦�&;0��l��%k䐸4_��[��Ƚ4���*�N�v��S�4��t}߾�A�xz,�_�fe�eQ�Gǌ� �|�#��������!�@x���S�x/��{y��[�I�s%�t��qf��S��A1�n�q��L��S����R�Ih�ЙK���9Q�U�*.T�����
�i3�8p��r�k6�kOD����� P�ɷm�'�!��~�pW�O?�����e�?��ᔬ``�2��Qؓ�=�6�p�1��
W�H�_�y���]���r:ɳ��<{V��*��bD[���������Abr�l�Hl(dq!�V�^��<��/�~C�O��1��t-���RnR�%;L�� Y��Ze��4W�g��F{#��]V���'ep�ǧQ�?�	�^����_��Iiɿ��u�#b�mZ�(��-�2|Hk�V���Y�ՆVb $Tur���:=����1�h��,�A(*cu�-�1��.a�d��||��%�\?�!xT�p��x�^roc��}��
�w$~i������0�¥������_�������?~�`I��7�,��jfJ��E�ߡ�kc��td'���l�?� �.>����q�˴����XLg�?X��ב��U&��Y
.8�G�Y��w�m/��fV��V��8#�[����(kߥ$��l�7A?�J~�e�<t����E���z��Eŵn),o ph�F��6-b��!@�U�br�-����q Sz�6g�97p�+m�GZ(�l-%��C��J��Pb%�o�܂�1�l�.S� _�0�ʎ�wX앿��m�y1�+p���cc^�������\{�q�!�k,^��g�T&	�Ι�L�2{?��7a�G��$�~��U�b��ok�Yt.�,�_�k�*�1�
�:�����a���fJPv�m�[�z��::��R�'���*��=�{�t��RZ���};:jp����&�ܴ=Ye����T:2�Bo�^��J|G�F��"��xú	`X���T����6���UG��M:�OGQXu��S�]�����aݏ5d����*9�)e��Y
�_�|��3�<VVk�OK�P��M���Nf�����>�sp�	ހ��l�0]��]��gޤ d���@�/���ad{]�ȡ���>���$�v���r�I��	�`�����'�|��]�ac���)L���lff�~M#v��7�+���W��?f����9����������(�0�ǌ9��lT���m)��aPY7���Z��t;�U�8	g� ��JE��r��o~�/)�{#�����><P�1$u�Z���g��``w����� �߱f��'	8���Ꮃ��?�����������胎��@���*�|N���V��{�����F�H�l5������S)~eA$�0zy�*�00c[ߞHf�]�:�}8�$j'�}mMm�w5�<.��Ym/�U?�UӠ����D��^I���8�-i�j7)�$���_�˿��������R���#�G��K��vA�s��&S{/��������O��V<����AmV�j��]�U��8&���)�mG�V���Rp��D�~�6z2͚"�6��xRp�ԾdO4�@`��\W���@y�K�z��Y>2b;%v��A��B�	����0!��j461a-��RY؇������%�J��<����{	D��-�艅VRa�� ������D�Ξ�x�0}�(K�y�����}NZ$ip!S��O�]ؙ�IK�8p��'U��b��{�S/�?�ζ�w���h�\����r͡���*$7���T�9��A���F��󴾗L(ʹf����<ж�R�Wɠ���*����<�K���z.^$�bw�]}���Pޯ?_���I�쫒���C��7�=VQ�|�7h��;.��+W�Ħ�A��-����}���ۿ�����g6y��PNFs�zk�ڟ/����3� �p|<��l�3����
��6� =�����w�C+[�0w./����+�e�?ǏA��:}u*Q/ �	�1g�-����{d�6�-�z�L���jY�5�z�� ��\��Cz��%���J��o��˰��(=fÀ��
X�1�V 6��A�S�?FQ�+$)���.�͈A ֆS�bm^i)�X&	`c�"��?8H |Az�`4c���TάfCuA���歩r[�"a�����X�,>d���v��p��n_�}�߬]��I��mg�.�x�mp��i^k���c�YA� 1����WJ#{բ	.�����]#R�hjtj������Kh<q��q�z�֝C�n��H^�EV8��տN�A�U���oe�� 5���r�$�Q���N	P1��(寓��d�1l�m��c���q�-`sz�R�t~Ma".��D�xx�/Y��x G�xr ϟ�����W߰���D&��0�m���F�(�},zB&�j�G�{�u�Ԋ5�᫝���3~�3+#̟�bb+�ŕ
 `���@�F���T������1��o�N؎(R�Ԛ��L`C�a�ڈI7�eɫ�4�,C�;��f�CKKL���}��m�����j@E�cT�����W �ߥ �/�˻�Lp��1�8���c�R�P����k$����ث��l4���JI[��.���b.�Gg����r���<���$�8�a���%^p_X�Ya�ɑ�.X���`*�qm�!�Cq������(��~��	�nH1L7H�u�-�>��hP�]U*G�� ��!#��*� ����!���C����HCl�%8���%_�_kY��Yb�Kӷ)�si@�Q��u���MW}����ױ1e�s�TPaca�Vb�*lJ~Q������*Ʀ���){� ��Q*��ϰ�W�&$�I}T	{�~j{_$�M��	y�{�=�T�qu|�]*�2�kR���]�>Ԧ��,A?璕���V5S��k�,��J5�d�Q闔B��s��>��?��W	���^����j�2�q����E/ȔTа�d��p m��KPR�FA;����=�8�:]�;Y/ӽ��&�S\Rʳ�C���[M�r��D.��:�#ꩨl�Fr���Y���)��'�Yx}oo�ryy���zC��m]�@����v�퓆��������ig�o�c<T��� ��0N˦g����T.���[mB_G���'U�Vj�@�!����N��t?�9;WjD��w��=�ޏ�z~=S`=nȉ�.����+�@+���_��?��_/�j��c�&���ǿ���ӌm��?��4a��Vp:���g���f��X��jpԯ�.�Ç���O?�O�h2��/T�`������}�Y�oE�A����A�M�}�/R������h�+� �/��9���@<�k��ع�;�Wp�`=�,]�i�fi㡛Ѕ�����X��Y�Ԯ%�t`��ʃ\��^S݇�vF���S�[�d)�i�9�����j�������H�bQb�����X��*�Zo�oVJ�b�*����+�dܐ����J?p�A5����X���=�3�<�`*\� �N��!j�=gw�t���ؽ��n���;{�h;�U��Eڝ����p�s�Vm+4�g�g�:b��U�ld<�؏�F#zr���f������~L��@^a� ˨]�.g�$��Rnu�E���D��)j�"(�K�5ٺ}R� '��82�=p���b ���zq th���5u��d��}��tol�(F�2�=F����HΎ���������R��ͷ�����2P-Q\��̀?��)�F���X���	o���SR�����0Ԛ��2�X���P�&�K&	���p5�\]��@r!���Y�u�:�o�`���E
�&	�u|C�{#����]LhFzs���zɷ�	]������J;j�F��s�9�k�x�V������~��\~�(�ɀ!��������t�(�T�K�5nAoӵ��3\=wP����q
 �J �w��7�c%soz��U�p��nJq�EM�y �ō���C��NfU峖�l���A:�}
]��S`��U��յ� ��Gk�/����`OA�~��WRݴ��(���U�B�'pX�lz� �+r��U�ւc͸�����B�=�nt�>:P��V�k����!VU��!A3�}�m��2+H�Q�t�	�;�CV����9�i��� Y�_�}/�B�\��=;��/_�UR�"m*���7N@�2ݏK��:���e��90��4�s
�~R	�f�JmL��1����SAi�6O��/u��'�����A �ʩX�l�(;�V{���6Ғq�zPAF|�x���` �t0�)7A��|sQ�5B��`�D��[���'y��'�|~/�aA�+�Az���D������r{��:@V �Ƌ^�)��� �ku�h�7�Ky��|��O)�=O�y��{ѕ\���mǘ�Σ����=���7�k�����l�DK(�Ʃ��~"�~ʍW�TY�e5���j��sYP���
PׄoE�|f�������e)�;d�	]����]�2'g�ة�w_�����Q�%W�������3��c��o�j�-��s����td�je��ق�f�VNK�W�M ��Zs6@k
y

�)���۰�����-'8�X������[ըzv��1���XI1�܄6�{7$#}���������C�!�-�n��f�#4S&y������,�ڂ�b,ՓF#�afM�5[i�t���2Y}�9��vZ��T"��l�AW�p�5�Q�8L�_��ɝ[�M�� ӿI��Z����]FV�oT��t��ѐ���xdC]���T�.�����!�A�����rzrJ�%m�VJ!zCpȮm76��ե>�s���x��e�������ri��p�?����n;�����閃��`���(�;Z���g� j��[KF��3�YĨ�=�-��Err��^�>��̓�rz��J�SsE�K�f�bW�$�?-�G�����=��+xU*�4�����b���Bu�6'RY��8�Xz��A_�#"C�}��;�:�6F{u��w���r�ɞ���p��@֡|������o����l��C�5o���y��S�
��i�+{
8��������`�I45GS'����F2Dб7��؀O
<�KP[�$��(���*��7�����S�c�E��dts�^� @�Z��?,O8,�9|v�
�'����@da��\�����N�{�hs0�*_b��������������w�)�X	��G������Gx=�2M��O����J5m��ȴ�G�����7��W��I`�ҵVIUE�룆��^<6���C06�X��+�6r��0+�X��	��9M 3�.�����?�5��Z�m���1T�0���B��A{-'P�j̈́=P�Rh��t��#���SD�����l��ܿ���P�u)vw�*�^j
��M��8(g\*U���Ҿ"�b��w�qFSqE5c��*DuZ۵&oZS�-=	���~�Lg��������V^�z��� *"��Yz2���y/^��w�ϺQ��׭�����������O�?�`n�8-r�j�d��������!�!v�/^39i�����%y������E�����}m�� ��Z����{2M��{D��]˕�(��RtC���BL"Qi�(�5`=�}�	0��yys/o�}����N�����4^��T��ʳ�D��Sy��9��ARIm�J�PP�GU��	g���������O��Y����߾K��صp�O��؏P�x�K�,���c�^�c�G���}Q?���Ś�ﷺ�cf�t�#'lۀ�&uߵ��J]�d����*��:W�5���>z����Ѝ�w�+�L��k����
��B�3]앟'YBI�Ȕ_;�u�Sp��JV����'nA���}p��U�`�$�CZ�ZZV�T� ����C������邃qQ�Z�6jض�d
j��h��OĂKΥ�5��I�(37[��4�����黶�k���9�����c��s%.a��-��Y?5��Q���˰Ri�RE�y[6�Q�X�
�n,f����g*����s��H�gR��j��?>�~8��3�.�J5��L�3���^T�3���ppP/�/0�.B:[�(�D�CC���Yr8/^Qn2��� ������}��P�Z=��BP{D�k�9�Ei���[S����
���;��˵��{XvV_��Ֆׇd �F!Ň�X��k�U;1@����[��k�2V=���=��돾��fRȣ��r~/'����%�5cYXC�m�v�[XJS[s�������)`��(Vr�J��@?��z���!W|,{��l�_
VF��i
��:T���Wa@�����v�ũJ~��Z������uȰJ��51� l,fAtc$���#9����p.�ΞɛW����iO�Su��j ��
?��(q��?[�ޟ����3τ+}NT�EH���j4a�	�A�����x����l��U���m�[�niY=���2��[������[9:~��h#�܃:�H���ҿ��E@[�J��������+Y��;�|:�c�lfd����F>~x+���.����\|x�
�|1eЉ�^�����
� pqoӞ��Ao���n�|��[(a���\$`�;����������J�w�&
��ws��4�b��hvN�"Ƨ�}e=(���NTM�����e����� x)𠯣�f'l!�� j��ud���D�|@{��.y�[��T� q�؃~v帶S���C��I���zT�HQ	`*�%��V���B Z�*Y�|u�jSQ��2I��S=4�Ǿ��P�8=y&_%�q�˫K�x���_
p�hS����/���� ~���C���O>�/	hm�*0���w�'넒ԥW7K��bUʈ���,I�,.T�}@l���H:'���?��H�����$�'��C4�y�:�P�e`@6@�֥�1p]�M��``�&<@�j�	(���dDv����������B{�t�v�	!��P1*􂏦��Y���O����)>]��}9~~ �H��	�&K5%���j�6n�tMn�-C.���ڥ��>\˻w���� �/�Q~yNp�Ĵ��3���v�[i�8�	k��F���濳M0���NV���z�se[����ŷ*��ű�ν}��Ei����<9[�5>�v��fg�P�t��c{�&��$��x��?��|2͠��&h�O�+'�������IVݝ�+ ��0<���WY�6}b /*-�� �Q
n���T�'J3n6���Ѽ�AdhQ�.�@.>_r�o� ��"1�[����+�i��s�]�}�f�8����s�_�N��o�c���r�:�c�z_ȑF�*r�+h IC���g�{�LY���$C!�%���Κ��aS�q�H�Q�ޓ��XƸ'	`A
V�j�.<��I�f��LVUN����~�!�`�퐒笖�֣�ѡ�u��*W��Q��}V�J�b4����Gx_�{T*+��v�@7��ӱ�YrL'	`�f1�|�QZ#�@5.�HW+��"�*�(Ϲ,�=�B3)XW��Sb�tO�v���p<y�x0]݌��� ��z�0%g�}3��8	%��8�����F��(�*K�/����ht��-��RBh��޾��E4~���q�.Lj����׿:��d���8��"^1,��X�1{%_��vC۽�Ww��_G]�u7��{$yN�$=����ņ$*�o;��2A����f�c�����\��)Y�ȼxpz��v͘�e�F���?ޟ`=;ܗӣCʴO'sV�����^�%�4��A������[/�l���
}y�ݺ����]��~ǿ'�3�d:?��������gR-�d�l��#���kr��?ո���W���!�)�wuIH���t�>�i R�N����@U�ڋYZY�S&�m)�ly}O��Њ�yZ��/k��]��Ͽ�۷����9���o�mN�{1�;��zf�>�� �k0T��41�4o��Ì'{9ړ�遜���o����z��,Nv�KO�v�D����i���_v�s�r��t߃�&� f�QG�O��p�����Iߡ���.i�F�1�j��l�A��L�m�,7��(�*x��7��P�;Q�/JJ���h�Z8�t���`X!P�u\ZϱQ��B+WRԶ���h���K�L�0f1}��������=I��$Q%���H ���Y�~��>�6���G���� �9==�������'0����P�U�YAZ��6r�~���2�R'��G��k��
�8�{*>�O��@�
F�1i�ib��.�B�ˀ�Q0Pa-��}�	��mЇ��Vz�զMǁ~�U
Γ=��=3��R���ώ�RL�S:�[
Ec`D��ݯ)���u�M�?)��@��Ճ����'��~����|����Ͽ�����\
<]� F�<:.�s����=��u^ob:�%�I���w�����|��O���gY����@��y����t�۾}�w�Ξ����׶�a����A�I&����Pş�.Ac5������u��`��q>�K�������mvz�+�O�>[*�UR|;Vl}$A�;�X �@�.H��J�����T��cw����t�_�������G�������1)���� BEV�*b�X���/TaP*č���j�����K�K�qz��D�F��R�Z+3�L��v��@B|vF��S���_aI��v�?�n����?/.[�zA�xN�巟���9�JjV(e�f#�� 5Adk�-%7C;�� �k=�M��&pU��m��Ш@���~^Ja��Z0#x�U�ʿ�X�ZЩ��>Z��$��,lL(�B2��e&y�	?%�[5����BY�p����,9(�$��ԁ ˅@ �r����͙C��ǐz/!�ZZoX`eP)������x.|�߀ hhe�(�q@,���77i;��]������=)9L�)<H��~Z���m��\�=h ]!3WE}yڻ�{�Ýɥ�E�k�[�iD��|�0�K��]������D�=[��a�
�W���sn�*�{Rt�0]����7Z���j�J ~��<�<��#�/�5��)YdѢۀ�K��1J��|�n��-���[��!�<Nu���j���ud���syyz$���p�*[at&�XػF��/�(�Z�$ǝ�{,�r�~'C�7�����/X:��b��d�^��y��/�/)�͊lP X�`A�a&;�}�V4�&��2լdu_�5�6�Y�� ˣ��2�7��z��2`΂bŽe=�:1e� $�М�`�g��� ����Ƿ������b���H�У6Q{�����>3ۇ=�*dU�ꋸ.@�N�{�0�/�^��AC���5��;�6��#�^������P@����3�aL�Mc�)�YD�R&�HA�Y�:�u����չ /�*�1�	މZIB��|R��`L*$|�U
��ݠ�aطӔ���SQu;�)��v�\��~4���`���Q�;�A�m4�'�R1��rU��sذN��m	T��Pz��W�{.Xό�͵䪹��ZnU�d�y>֛I�h�8G���zOK�Z=W� U!X�u��1m'>� �b����s�����j����^��ׂV�)��2(���m6'����:Q@����1��	t�~�VhH�@�s��A5Ik @𿨒����<���s���8=��ްZU[�&D����"� �hj󹎍I�wu���_~�?�i���fi��J�^�U��}��A�9�P��Pf�bZ��R?ܭ���A�?]ʟ��CX���?�,矯��`U�����,ԮH=���?��Ԏ�~�z���;�e�D �}�U�����ь��q��Ե�ͪsߕ�M��ɞ�+�N���9�l3Ű��b��bp3��&����M����[�OW��Ų�v�B�s��
;��\g��,4��_�`��~������D(�+/��r�ņ�ֵ5�+寵���df�i���<P}����W��%����J`��8w�v��_;��nB���'���d��JY��øN��1UG5#�'�^�_�f��8-i���X��e`
�t���&�9S�<Iߡ������4Q�EC��~Sgi�r�ԀƤ��.P�� ą����+Z��5}�5�7�;�@�i&���cۋS8V�ڡ��5|-�HZ�a��9��l��b%>��UBB�q�pO��#��Cn��� �e�,Ѽ��~6M��o��(W��WB=��	a���t�-v�����9���N�A7?�&(�� �_E�4�GU�d����7@��� ��FAQ����@U�ϭ�����w���~Myl��7�4��"�N�!ڞu��M��	F���;�i��m&E�ϋ�gV�����R�P@7}��x�B����?�SP�TO����~�M�����>�Q���sõD��R��+���!��`
F��d>$'.�����/ |rD��3}4~��/t,�f��Pz�l��U0'���}a��{X���Φ�z,�~[Za؛ͩt�M����&�K����N�O�/�)��X�ڢS3-Xh�Ry��X��g�a`.��ᖠ!�d�7�,��8��~8od���ٕe�xgcv�ӹ�0��{�g�-�_���ӧwrq�.�|�lփ�A��p���R�%���eh����
�����K�&��Pi�G�r|�R^�|#/_#�g�\�L�\E70
#S4�����|��}������h�����F��#���$3�;� �Yy/�.��5R�T�o �A�9�0��1s�`1��nRЅj���)H6�iL:<�2%@�=N�-,+��JTI�|sXy�� T���Y���9���ƀ�Is��1T�+�'��F���',q�*�
AնW\�`��b���QR�L�<���N��QHZ#F�<*f�j���X����ʀz�hɲ��:�Q �(ɚF/|D�@���쯆G�S�����Re�>��@�8X!Cx��t:{ ����#P�����  D5U+�|��\���G�v1��ysR1�����J���	��X�dC�t�c�ǈI��}��9pK���3O�b@� Y���#�H#<9>$�f2�iG �uuq#�?��w�?����/o���g&���1,�o�i{�Yܿ�3�O}��G���^����邽�U��u�~+���8ɫ�1�5�+�J�M3�8��N�������Ul66o�U&Π�VQeP�������9.u� {�b���}����.�g��3&�DM���,��G�1�_�sbF$>�q�a��m���:�<�ӌ,N�E�PU�0��7H����b��������ù|x�I�_P��6V��)������F����ZUЖ�����SF�E�@3gȢ	���ɫ�v�M�׳�bw^;��J]���,��p�@�I�f[��ָО-8d�(�?PC�LdQi�	�t �Tr��&����b�\���@g�r}nYz�o�,��9hsK�f������`A�����f�2몢4@��Z�A^r��ڄy�lЋEǳẀcAu�A�S�a���JW4�ͩM��)89�W��^9�A�3s=�����O�]f�m�����Zw�t6Y�j[mi��B��Y�`*M�aѡ�t=9��> =sy�=�a���)���c����A�`�
c;&�KT��� +��Sߺ~5�F.ca�n�hA�� z��� ,-��������OroV�vj�X���C�`k>_0�ޞ%g��PD���l6�;����줲��NȀ�]������:[��F�b�d6��E�*�b>���t�)���,z}�~P��.����gc|7�lˎ�qj\����_�׬8�g3��/��TуA��z�Oy��j�Y�*�	���<x7�!y`o`�I�Ri*����e�d=���q�l�m�識/8[y��]Ї�ւ��O��6�����J�VJ1����|��V.�>��-�`��v�w��)��fU�����}j;���Ri�M��+A��'r�⍜��J���J���O'�>ib�@��(��k��Y$��N���������������5� �A:&%��$�����M���r�oK�'?�hr����FC���	�����t������ނ���ox��#�Ɛv6������������E�wؘ�bi�u�F$�����Z�,�0)|�B4�U��� ��N+���Xl�\O"�FAG"����	vӋ�h}Y���es?�ɇϳ�S�1$���4��� �>~���ӭp�jKJ7�+����FOyUY�F��aI%�\5�Z����9�-Ibq]k�m�Hd�U������~
�:�8��Q��-�Mﻘ����4}?�
�& u�?���?���.q�+��٢0� �T�S ) �Nܦc��L I�Yeu�^��(>]��|/ٚ���ny���5�.�[�,=�`p3Ķ.ϯȺH�s����ҽ�,��/&�A-DE�Y��ݳ�����'�̼~Q�ݷ�� �Ȓ�I��������6[��X��{�����n�6�X�_��,QѼ��\3Q���*�2���4��b�ٮ~%��֎#��z��?�2�zߞ�Ľ�z�}�2����U0��Yq��JG��YGF1i�p�O�r�l��t˺���
QÓT�q�(�"�"E��Md���<,p\��`$��	�xv&����%��r�����A���&��4٢�\�(jQ������*Όb(۠��6�R���&NϤө���!g���'�qаy�epk�¼%��B&�6
룂1*d���g+��Ӵ����5���M�-,�Y��
�t��^W��6JW� !.l9�Eg�Tp0l�*E���<�t��d��e�x��Ϡ����[q:9��}
h6�8&�S8�t�[L�H�/r�eA�U[y�JR{	�%� ����" C�e*��/$���9�ͷ��NqSb�n��q����l�kr�G��K65��ɰ�\��JV����񘊴.��׼��|�5�{kCYYA/�Ii�+Ŗ 3� �עVTK����Ӆ��&�B�9_�}A��w�=i��t��@�RWzo��z��F�(���u�a=���ߠ���jF*�)��e��i?�}�ai�� #=�B��\����4}��Y�������A��vk�M�*�Qgm������AwT@�J��"֭�ڨa��R��j�r��hɾ����hi���4!bw�)OU�{{A�h���I�-Dt�[.u�o��z�j�kqh�@N7
��r�Jc��왪K�D�`@�B^�	�3*Ek4)s�4�2�~N�)���߱g#�����;iC'~z�L�@��(�vtVSi��QEkBS�$O�	�!2�ʓ_�C���$��hK��*��=O{k1�!���o���9���xC2]�����jdٮ(| �8D���Fi%u�l �gL���Ve,+7*�r}��#�������L'�U@�1ib��43ٚS��}�N�pI�yT�/�ZO���e���+��M
�ʴ���c^��c>��;n�{6��ё�u��U�,;��9S�W���d��ᡜ��ZN�^���Iڟ�x�dC��H�tCF����o�"xr��ݟ���x�7X���c�/�;U������%��k���?���?K}w'3�l�g�k�,lM�ӥ�ٸ��Y%���ߨ߆HR�6t��OI�c���4sPD�̊��-��[6K ������!z�\`Zl1\��`�l��艺1��q��X�
@�E�_��:��T}�˴��:I 2JG����f)?��N���򜉇��9�N��p�����Z�)J�A�m�9�����|q!���"����*��a7��� 8|�*��6���-�[WT(�x�Z  �ɏm=z���RO$�8��O����*EL�����ۑJ��V���R��8V:��=O>k��gs�ZF��>��o"��^�N���-��친�8��g	t�od0½����>���L�7��^�t9+ʿd��}�=b���@s�<[���A�[ �)�I��6�����t}�B@��V@�.���^f	`A��g ��;�m-��X�߈�0����Z���
݌�������sm)�Ё&b<�p@oR��&��h�0��AT1�&���i|��iD��F�w�/~
|_��	`��*g�-����z	�	MÌEA���V4l@��8�x���%6����̪�=�&N�T��@i���X�?�N�5��Bu>h��+�*�V�k۵�v�{���=�[^Ϭ�����V�gsE|�yc�`3��:+=ц�%3.��\�����0�Ji<>�P��ÃCy��%��l�=E�d��T�}�-�,�JF��^5i�ƕQv�*�����}�
�݄���~
[�v�^b���GK��,��d�եg��|N�FF �M��L��О��3�i`$���α�Ʉ�ɴ!���4
N�:�N���s/J]�\V�O����əF�$Y�X�P!HN��DVz�M�P	�2�)���^1YQ�]E��T����C��)��c�j�j��/���pZ��$Bu��䊨��̺�w�����ѽ�e���R���啛B�Xl�)6[� p��NA	ƢQ#i��>���zں5٬K!P��j��H���S��h�<����eU�����z�vβ�)��~Ŏ+��B��}���Gl�yьn��T�.Db�|��l�8�y*[θR�������o�-��Od����1f�W�3M�d�Ю���;<��c*PEŚ+z)2B��e�|hU��6ʂ ;] � ���0�{���TqB�	�j�kN�C hJ;)L� ��A����]�_�o?���^�������A[�U����H]���]Y���.Tu����+���`߅I�[ޭJ�AR	5ە��*(��)�aBJ{4�JїZ���@�dol��ϖ��oqCۂ֪߯X
�@�4���a��{Gq(���Q��ud啶�T��d6���>��'�V���Nҿ��P���x(m0>�3���� �_-u��2@�yv�_X��پlO�>���6��&G��TF�����d���M����(�6�V������ES��FE�V4��+��D��#�{������S�P�힋n���ഩ+*�%��{;A����� ������D`��
�P��d������qV���???O�O�7����[�Ι��x@�-3ܹ�hq�M-���&g����#�Ͷ$I�,1Q5�5<�\j�3��S��?��e��Ӑ�i �*���f��{EDU=2���C:����آ*"W���)���&�[%J����,ǢD��O��*[af��D�|P�R �u��~yy!�^]���F6�u�����=�>��������_�1ǘ~5�h�he��z��1Ȓ�b�z/!i�������zʶ�x�v hK�Ge��c�͟����y?��KMb�^�m�WP�dW���dT>����X*���!��I��*\�q�'7=�Mg>AM
$���-���&6��!�}J%a5����߳����d�S5D��8��^��&�n�6ۜ�76������W8У\�Uܜ�-;�!Kߖ�j�W��$�wZ�����mz�_�bΆx
��A�79�3h@��ar�?Ǽ������7��]��ľ+��o�p���W���y�9�~A	��Q���Pcr�H͎z�,���Jq	�o����뽬+�㱝�����H�a��˪b:<�TҙWb��7�;7H��F�a�̑7�q�W������f�n��v���t|VG����d�\��x�53���CE��-�;�`�)�3p�G�mP��DP�ɫ�Fm��vT��BB�X���Z@����Q��y =p����Z�����Q�MO��J:�;�U1���T0�zț����U�qɯs(��ʃ�����٥�ځU�q�`���p`����JR"���o#�"�I�h �絹�ǆ\$�g�J]0�ج"�)3�a*k��4�C��}�ˑ�n�����)L�)y�����T]�ޛ�5`�e=� X��A�0#�����p�&(���y�=���X*�3�(�S���|}�>7�9��E�vCg�DK��w�^�E��Z�g����m��.8�b�\q趈�,���PA���=��M���5Y�oy���Q*��$�`�-�b�	��0����.4�z�iȢvw�]�ȯo`&)钠MZ�fr�^0�C���$�c<��S?�v���1+M*ۑ���C�`Yk�j�`a�Hw���d�-5Û4(��M�nP�ẗ
(��E�����*�ik5 ����n^��r���u~^��2���E�jm��H��	"��﷠h������T��db/8ǋ�U����ë��t�!/�=�P���������&�T8��"���yD�|-J��,5h*��79�ю�I���E��5�d.(���f�ʨ�.B� ?�B�Bx�h�ݦ�u���۴Oe��FJ���`��y�+Uz�$eg�E)T�	��؁����m|��7�*�-��S����5&�}��v�W�+���:��!���ڋf���+6@|�k����#����H$R�pA���q#�����:�%�M��qY��.�HM�o�� �ȱ#�&>��$~}/�w�}���l̀V��r0us�Ƀ
}�.�ő֋�+�6Y��'MN���v���L������ړΩ�hE��'�m���r/�uK���J�������3V7fI�W}m���z�i�ū�W,��d(�m}�m$���h�p:L�Ʃ���%�L��hxe�P��꡹(�~P鋵,BTuo�x/�K����S�=��[I�����?3�n%����Sk�-h�����+5*���'�d#����#���� �O�����3^�@�� %AlR��1��F���o�w�~���;��ˌ�*����$�6 �P~2Cb��dsJ�&8�/`�Gj}Rj~־�nv���B�BHvQ=K�ޤ�֩|ST�Nف��p�{ c{�2r(�:1�9�B`^3�s�lV��
P�����SiE��(;(:o��2#���],A?�&��d�4�@6�D�x���P2HFmF���bA	�0R�N{"�86��E�<e��嬑��<�@���s�b�s߁�
Y�	�6�������,H��R�a����X�!z�Y8�&��w�����M�`��3��=�C�^��A	z��g�`A��{�jT��gcp�k��d���5d�:�$���J+(�]潘��ի����L)2����dʅ������?���,@k.�o_��f�<c���z���.��\PR3�z���և9_�4���<���G��^{��Du,�t}	B�Hg}�^1�7�oj��(7��%{�KͿ�(D��&��;�$�?'�|r��l�M8B�8�ʅ\^md��p��`;�����Rr�D��ߧ��:��#<���]v�9�s�Y>s y�*VƟ�D���K2�NM�oδ�S���Q2��DN�*�nfs�Xf��A�K�Ä�Co��d�Y���c������{��b��Cfw\��}�/��J� q˪���W6�Xj�-�f
��P6"*�?Xu�l��+��M*��_���dXn�!"�l�RP�6�����ˣس�+��+����8"��D�I2H|�|'C�3�8h��[4q����(.�y�7��:*�#�_3�����p]{�V)L��T[`U6g�a�w��
�����'���T�~��߱��嶣�kM,�fsL�i{�US]�U���Kʎ��㏼רJ�I�)���r`3�TA椃uq�777���h�S��:�R>5I�
��zp*�Z�p���
���DKi>��o"�
b(,�n �ױ?Z"|0��'R0�\K�!��#Y:�{���F��.��-��k�	bi`�v�X�?gʐ���Zb�A��#��hY���T��Ӟ����J���4'��F�_M�^1��xKE�\L]ϡO��FT�����8C�c�3�X���39f���E��/>�G%��]��w��^}cs/ƀ�9�Q�܀s�TWQ�*��0�DJ�W�_��}�qlNL���P��M�C�5����6U�
�,6k���@ֹ�tP��s����Yׂ����T~^Ѱ_����y5��� ����?w�d�f:_ٗO�>ɿ���?���\]ް��㘃m�� �z�z&o޼��n��|������rcl6�l\�PZF�������]��P^㬧I��_h�`}-�k/*�,�TntHm�Ԇ�W� ,����t��gj ���#�)�U�o���qK��jN�=G�cy&�}$,#Ј�Pf_��8�r���'��X���8�`��
��1���L~���$`�㻊��1��ٰ�$
�f�yn�qP�:�����ϵt̪�тp?a������N>g�����?���2�zp�A��^P�y�ힳ��{TG=� 눾�
�4c��&E�*]������	)(wͤ2�(��K��&E?c߉@������o�o�;�bZp�k� 7�!�w Վ�m��w��=���O����R�d�F1�b�ր
�;7غֽ��5�/>���bg���m	�7X�Hr���U�N_��$c�OЬ�Ri<��PMP�'��nr�n(�9�Ǉ������{R�R��h�&!�,�l4?����ɲq��)��M�W����n{�<j�/_�z٬{Y�a�r�0�H���A�f���T�� ����_�$Oh�@����-���
`��GXDϗz�ۖEr���悲�KR����R{}f[>��8��yi�E)Y�0	�l&��h�J��u�g���u����L6&l�l6��b=�qC>$zF6�X���08S��z�:�N���x����e�� &�t���-�J��g������ׇs�07���wtfӞ�f�1�
������z�k�?�Q��4�I�1��X�]�q!W�ײ���*#fc�+���&�ofk�H ��[�}=���\�����B'�ule>�z�z<$���v�4�Q+AL����`T�@=3P� ��b���_�[ƏӤ͗��� m���BQB��LT�UM����?��\������Ĥ���ф 4Q����@_��i�j�q&���w��3���+]�ҽK>ĂP�fH�!tFRl�Op"���x�i���7�s� ��牂S�^��w��`	J*EN*h�X����O��０�,d�5S
p��Dbu2`+X�`�eLbA~�1�m�C�C��I�à�nM�+c���#��=�a�3�ii4`:Yo�&j�6��̟�Õ˚ʚ�i�"u,`�y�k�h�W���ܞ�%��`PUZ�%��U�v_�_[�ă�P@��c�D7���
��wt�g�;�q^�ۮ��.��P�Z(ǡj���IM2Į�U|��YL5�,�B�Vξ���M�ǭ^���TBo����/f���#��̙��)��Pe�L��L�ȋ���}�)��W�{��`�ݳ�����8G���7�jbV�S���&:�싳y����W��h��./׬PH�����+��n1 
�Ɔ��*�E�É�����р�����i�v!i�G)�hno�l�SP�Hd�3�!�o5���H@�Bp�)�C6�b��3����:�7�[�'���=F��u�B3�H�pԡ��o��)U��F�TDU>�f���]ҡBG��`U4
[��7�$�S��e:hXŬɁќ�,�t{9�KNt"8�7n����=>�X�`��D�7�
6wX=f�����@j*�q��Ay�����#�@� B��<X����(^����b�������D�� :� (���ā��_`���S|2*e�Y0�������k�x�3U�|6l���㣊o�7&S�IJW����Py�~n��?m,Nc���{���Z�1+&�q�^'T�,Bо�c�с,(�'\��r��u��`bTD��ghL�����(����@����T�[[4 ǐ4��S�{�����Mf08���]_.)v�Dvb:P=m���e�Vړ=6&��zQ_���W�m����W�[Rq~ʫZhՂ21��k �53*�-):���2H�EU��L�A�;�z���ʤO��UrH�� N@+���	:U��7U����1���5�%z��>��*��m��C��Y~o7٨	�8��W�V���~@8�3��i��| �h�
��r���? [�����Ff�%SGL��&�J
����YN���#�"��_���f�Խ:i��>k0F�xA���V�COR����DeZʨG�j�q%��p.$�ɑ6l֩�]����C��%*�áýUm�:G�頷��}x�Tʽ�N��<�[qф�bj���.��Ĺ8!��d(�X�����)��Q������w�c��@��/�o�
���f�>�k�.d� j믿��V��$ih��)���'߫NgK9�L�AHR�E� t{$:ݳ��+SN��5x��	��6`Ť�F�6�QE���ڛ?po�Ã�*[+B2
>ǉ5��r��{(��kx1���8���AN��(�T�""b�0�%t`��lإF���n�O��<?Z��&�chX�\�!Qnb��6��D?�-�V�
�Ǣ%8��%�Rm|� �w>�^�����(0bU���Z��JnM�m�Yks����$�f�p`��eq�U^V��V�j�^5Rg�*x�'[t���^E���֓՜c9��C�(��?+r+����E���9x_��"C0�9���fd޿� �������e&�����|��N7�t:E�B�3�F�Tf�f�M��y6�Γ���d�I��S��U��%�,�\B����q.���Y��;|OX@�?����x���͆~��*��Dc�OJ�5|-(�e*I���cO0 ǳݢ��@z�
��O~By��\2��3V�d�@P�gT�t��`s�d�����̢�zv<y�0�%������ �ǘ\?X�'���JÞ��0�3�	�����3	�yll��,�`��^�&&>nwS�͎��ᙕ*���8&�'��-�30{� +���0h5k�>8uk������t3*���R�=[^Mm�FY(�f�XP$&��4X��r�#��g %���.�[2g����1�.�.;��@�_�@aT�+Y��@���.ٿ�΢ѽ$�9�yt
޳9��l�b`��L�ה�b��⦲�Bd�ʳhϮ�d:��頠x<�0i�E6���VF��$��v�簉w�mh((��O�ꉂ=ˤ:J���8�5s��
�A�V4���{�T0��Cts}AZ�Ųg5��֋����x��R<�H%%ʹq^��I����$R{�R�*vR~�a���]A�S�"	0�YPP�B������(Z��+�[���
�b���=��t��f��bH>>g���y*2��5ك
8��Ѵ<�7gd�����-iX�p�lÐ��h��T &�㊵�da�>-��J����l����,zY�Jf4��c<qvFi@��X��M��f�&��]g�$j�	�C�e�Y�����������$a�!xyYйl*��Q<g�\S2�	L�l�qO��5��b@ B��% P�ZB�<�[8�|?����C��cp5����M�!`>��ug���O��h�<�:p���h�p,�ڪ�8�Ψ�L��x����	yV�R��c��\Y,n�q$yM#؇pů��Z�1�K(��5�H ���"A!�
�(mR���)8{r�Yd�pW;<Y�_����xD}����^'���hgO�$G�-��h��/���kGL`Ȫ�B�БO�cM�jv4 6�y�_�ɛ�E�{k�����,A��y��Xi�>�#���w���L2����P�㸊Xm���(M�����]i�	�SY�/�נ�X�d�.^D�UXH�ޓ�1(�
6� ����#oin1��.�}��	v��k/�x��bj�FjOV�L.�qN�s?YDX���>�i~�m֜
���R�����#�x=�`��qdo�B�L���1����+���\,u(?m�Y�v���yD�vu^5�:3�@/���L�N����1��ϐN�h�D� R�)Nn�iy��@Y�h����(C�)øGp�����d�;N	⁞J��LNϲ;B����[nh�WYHeE��w�D	�'�Ƞ*���c~2;�>��Ƀ��T
�6��⃬��B6�r���~Xs�6bT0�N�=&��Cu�I����rx�w:�Z��N4 �i�`B�0��IQ+�]w��?"�9���r>DY2�x�4/{�P�:�5F64AȕӁZmB#4�9 ��F�O�����$�����,�90:�.�:��gYLp��H�u���,���!w�W ��L!��dp������:V�T�]����@(�B
(�k�{G���6͎�������^J�?�H��|���ᳱ^b}�ޮ�5� k�������6�gPj��?d��c��֬h�'���*�d��	^����m����j�O_Z��I�	g��2K�2���y^k�M�7�V���`�Q�[�&&xt*e�ь\�j����0ɞP�6|���`ߩ���^�Q�3[p�����>T{�TQ�-���UX���
*�I�cC�
?%g��dV���3��͗�sq�_��{�<�:.�Xr����Tu�v6���;Sze_F�!�3T0�����G���:���@�Z�[����E����`��]�ɂHV�3��j�f����ӹ�0Ȋ�@'�30rǊM��B�p��<C�-�AavU�݂��Ω9���}�<�O:6�4L�w"�����%�"=|�?9Ȇ�H��;�ro��.<�iV��4��Q=��<q^�M:*��u"}``4��$����~����z��.��S���._/QpM�s�cd��QV����*���V�q�EG�j��XjK|6�Ԅ��k�-�Bs	k���Z�ҋTyyT
+S�rׂ�=��#��R�������9'��3`J�b���&��N�%�c��q��&�xw��Q��'�-4���j���,��8�h� �[B{	�u��������P 2V����,�ăҍ�ƞ8�1B����_����s{�^��`����c�QYf5��7\-���p �Ǻ����k����֗���,A��q~���Qz��u���W���U�����/mw��$��GѤۨ�BF݌%^�"X�88�7�M���oo1���_C~tV�r1�"b!%"���؎$u_����J��ؠ�z�=��+��C�������"�c�}��iRO���w��o��G���k_�k���nZ�^��|9oҫ��E�g�ސ) �M��{�EO�;ΦA�|sq��T�V�+��]Srs�L/���Ī4�����$����2�u8_M���~E����e����?�IΙ-�G<{�Y�P�h%˃ә�m5Ki�������67�r����۞@k�;�q_�r��0Z͢qD�,��y��2���0�����if���Ώ�*����r����*�7����I�_�T�` ��
!���^7;om;���&׬3PQ;��jw�N{OC*���6�g�Ĭ���{�X� k
���#�;rN��3�Ԙc1���3!=�?9�}G�c�yh��c�wz��i:�7��<�f�x�F��W�ꟓ+cN:X\j
[��O���b�ζ��␃�#�/�tÈ�_Xō�c��G�~,�f�OM��w�����;�)U�E�䃎OR�T����u�J����7������%�"��EE�ޯ�p��l�&0bv� �mo��)"hf(4�9?5
�2�1M��`�8>n6���Lz�o�O���˫~��#U�B�z��*u�,�r���k�B%s�ؓv�	�)��]�ɒH�'Ѵx�����4����տ�����Qҋd-`2�'�i7�t�_j��H�Q�.��{���������	s��x!M,�S�<�`�h#����}�5�]� h�fZ�Y2���s��ő�ȇ��x��:�0��qG�!*����@n؍�=<�<�;�xQ��[����r�Ϗ������QU�x{�:�@p
I��[�^҆+rxiu���be�W]���<ٝb�[{��ao)�����+}�L�{�m�z����n	
h��0��0����B0���	���)}|�LAxdU�������AR�(4A�BOF7fƂ�ҋ�e�E��"I�~gլ`�g�o�ʹ*�$����|����i�]��� ������3�]cBqv軷�1��X	�	}Y����B��T����8M,��)��n�S���,M���#�ǉA5:�;�b�4�F�@��D죵�O�~M)�����8�0��)U���_;�)`�<�?���[ΟO���E�p`8�//���k>�!�s���d����b>+[�Eϋr��Z�ޢ?�>䔪����x�M|�7��{�g�OX_%�w8�
M%K?٪�5Y��5z��ڵW%��O�d�G2��X*sj��jW@���IMvF�Ok��PFn�ؓ��5���i�ఉ�۟�@i@�
u�����9�q���e��{�ݖ9��|�@Z�q�� h~���dnM6��9��p5����޼��i�u53_24vA�+p�ҹ�I�Zil�y�� �����������Wr}}��:�%(j���y#.��4��V��}�R��#R�!1��Z�rp(��?'W� �[pju�|%�{<�NM��CmA�����͎-8/W�8�C��L��Jv YT\�N6�	w�׹*@����Q9�Ԛ�!�O)�� W��с�C�f�rv��&��#�uT`��@ը4u� G������=?�������w�h����.�����|�ӧ�O�emI:�Wұ����c|B�����3��IC�� 5�=�v�a<ڰI�o"���|� *
b|:!��4e��G[*��L�����W�`s-B�j�=�#����m�:iUh,���`I��T���G�`y���������Pα� �N��4yr��2����@b��:���+*����.������$�h���^���BA6[�@�C�4��lO69�����A 8j&�I\����[���Ѳ���5���ߓ�{�[��d�j� [3���k=Q����L�2������EH��:�%�a���H���cN_y��;.'X9����@��.�u�%�F����v�� ��,.֬��H�ge�mU聀�!���������#���j$�0b,ax(Ujq�h�bU�K*�0�Y}Z)d��6� ���>����q<�	�ٰ�64)�V�/��"�;��0�]|l�}���nAV���뉽ٻ��U���=��?��=#�[��w�1�
m��r;7���倽�G���@O&Q��l�	F�q� z9��^.d�8���=|T�;㬳6��I7|�Xhj.�ѱg|d���>]�~=��6�
�P+��l8���5;����De�sA���-.�-#����/��2� ��~�����ǵ��W��A�5���}�V~���X]��s�>>|�YY	�(�ީ�`t���m��������6�:�@_j�o� {�ɚk�o��q��`!	�`�}�����Cec�@����#*Y Yo���1��M
"�g��CL��U�_����Q�O{�ag�9~٢�|�{�0�(~l�>N5ε�O*�'E�g�3��T������!'V�{K4��� @𿘔���v$�h�nǲ���B���L�}v�#6V �V(��9��WČ]Pz<�&�y�ZIv�rNZ�G�������6�&-lA��s?ٮq���z�yi��zY[?��zrn��#%��5�j�k$x���B}�U�}r ����$��Eo�7k싂�~t��:{e�F��lD/3P��\� l�[yx��]KǓ�����;�5����c?��G�\ [#�o�f�zu%�}�Z��U6�=� Nj�K�))�U�"�g��)m�����H��69&F�F��B7<D'lSX�� d�N���Le٪����N)\�mg6���+�&�=��$�R�����᠉��\t�pr�y���ZR$BF�4"x[�R:m��f�q�E�s��Y�B �-�� �D����A8�өc�3��<mQA�2 �K�Y8�K�b6S8v6�5��&d�O��u���:��H����t
T���v��%��*�e��iy�F�a����os0�5I�IA{>@�u�|�=l�T�;�(�������`g�lt~F��g��m�|m׬ �5�ӡO:��V����Z��޾hI7��|Z���&)��Ա�t����/G�s��ՠ�\iK��qo�$]��iu`���#vXBiTu`w�蘡�D��S�E^pW�;i�*�;y�N��j�^��kΉ�9+
�y.�KJeg�1 �ɒ�`��ޤ�=�8R�N��s��)c$j��7���lS�k~>�S�)T�p�s����$io�x1h�ְ�+��Tg�@��F����mD��S��c_�}|����j.?]d��ު�]�=�����J� �z�����#�s�0�[H
f�IGR%�-�,��y�(�q`���M����vw�7��[��cg,���-L�7 ���|]��WFAź��X�1�d����6+�\����U�O�l�<<n9kh��cu�a3�+�(��˵�kd��~�y�A�@s|oI�_Z�*NM��W%m�Ǥ
�*���#��k��mǎ3�Р����1��gH�?�9oU0�5���2�����o���w�D\c֥�{�l����M|�%��3�=I���ª�}�K����@˃���%O�� �+��pϑ���G�K��w'�� ���!V�8� �ͼW��G[	��6� N}��WQ��@�}>ϼy�[�{���Y�j~�~�KR7�&1ָ~�%'M(%�*��6ZG� ��e �?XR��u�wf`H5z�4v"����8*hR������8I�� �XG����߳�������ӏ*܂�F�0��Ϸ�3�&����s�su���u��+������/�?����_ɾz�d��P	�lMF[Sp��(�	=_J'	*��4��l�`���T핽DA�X��knu��*�s9N'��;����SA�æfB<m��e�v̾mJu���a/�O��}>�����}�?s�=������7^�U[�LLӑ�7�|����dQٵ�ܾ`��:t޺��A���*Y�]R������/�B���llC��r���հ��Q��Ԋ�X�&�)�J�H*~x�c�bh��3�<ҧ����s�t������3�dg�ò� ��.U?)(�9�G�B1%��]�Xؙ|��D/��0N�<��&�8�5�p�Wɩ��(Y����� *>�����rD�=R�h���|G$ﲽ�@��ĹkH�")t�k!I_�92��E��ţ�vI�lh>�ێ�m֞sB}��x����j��D����O쳡��a��2�2>�u'���'�г0�~�$�1�����,R='qqz�-T~B��eo�8�&��_�����3���k����=Yx&�fMF�:I��T�
��v�G���1o���EN{�`A�$�!]��B�,R�	�ފ�
 �#�Z� o���׫2"z�*k^!v�&=���� �PF�����)X?O�7M@�*��n�Z��=�����A������4�m�����J�E�~dĘ�V6���2�aV<�yed�<7�U,�rZ���}�U�T�X�!�q�%%�R�[��f�k�4:ZBQ{b*:��A�)��P�t��������XϢe)��jrA�Ο�.�B��`Ԃf���r[��LgV�m���@��
�&�\�M������������43="��QS��g��������k�|�y��N�4��m^׷w��p�`C�=s�J��&Tx��Sŋ�;U�7o�� �pA09�u�K84�a(xb����8���._8��,��*d��Ӊ+@���P�2N��.I��>Bs�����f}Ij~�����*4�=�V�)�@q�%MpZ��T<\�E�����*c�%g�<���=P��4|�QPZ��y-�ׯ�bs��Յ,Ke8��&2��A+�rڝ����"��1�<[�I���ٳ:�L�i�X��� ������O�8" �� Z}���$�e���ǿF�r�q�����WK~?l�`B.L]rd���Ѿ��z׌⍴h�Ռ����>�����j&�M�IL�J�}I(T,&��*�G�^�:Z�`��"���LOy������'��J1�Ty5�3��Z�H�ϩ�}q�t���T�}K&-�*�wQ�o&�ٟ90��:둴�U-Ŕ���6����ߪ�.����˼�)%���C���c���n���/��7��G�� ��no�.��â�f\=��U��m'O�97Jy���O�>:��@G-�'^{�A��S��h��n'�p;�x�a�L��/ܩu���ӏV�HT����F���.hU X<�Im.?��98`q������f�$�O���M)ߚ��j����:��^g��e���{�PY��ɭs(oK�!�I*~,��U�I�k�^P�RgI%�z�[n�C�'�V�<i׊��J }~~_/^S�3էxl�?�����'5�-UA�X��*Yv7=�ў:ę�#v:�~�XrEu��"Ds��Klb{�*�e����7�>*���Y��ĺH��+���/�sC0�N'&cQBu�p�������3���I��t���B^�����rq��7�����R���}[],R����c��>�ՅRZ(�˜��T�_d@��I�����{5qc�;jT�wc& ,iI��=7T�m(�aT/.��X�I�'x]��:UO�F*�t}�&;�ʜ�l��^sPz��$�5Q�C�W�w���+CwS��VP���P�G4��0���!�z���EF�������@�=V�����E��26DfЕ���������?|j7*d)v1hU�&�Z/��IìA�d�m�JC����
�u�#�Gj{ߘBᇻ+Z���#X9��9� &�X���9�0Ne���U8Z�Ո�@�ȓ2�@�T�_�j��G��b/���Bq�X�T:����]��5��~�
~(�=��:�8 ��c�?�*߼��~��ʦ�)/r`�5�L2z"r�������}7�8wg�f�]a�?*�gfQ��� $�yϭA%��93��lyD �}�	�d����e���q���A���QR�NF�����I��u�&ς��)���{����~��-����ߕ`�����V�W`���3��l(T���K	��������@@o��Г�Z�dsy�A�M[��ba�+�TF�Yv\lM#oa8�� ʜ�8*6g���u���dR/P���_nn���Y^��I{<��&n�����j!�n����!x��PP�P�dS����+a�1*"1�����p�U�z���5�Ae�̗�%�&�Kv�칤ڻ�L���%8\�Á�8X�>kRjg�p϶���:��~�I}�ɛh��	��B��˒8�����>Ap�����M�uO�hN���eLR��&U/��-��������׼�l?އd%���c4��G��hFq�W����E�7�:�֋L��ؙ����<nj��������RQ>����`��,G���k?�d� �����n��0�pd
>�xd�OJ1d���-RL6d�I�b��}ը.��,�(�jN��9�"+��ϣ˲�Q����W��z8n~Z%��yT�S(u��a���'�y�gz
>M�Z��&��j:���N����z_� ��B�$\9Έ��zQ��=�Iʶ s�R��V����J�.�
��	�Pbn7��$��z+��5���v�QT�fL�J�8о+Y���ٓ�ڟ�d5��s8�����e�Y6��n��vQuC�ų̈́�� �U����ࠊ_l�5*6'>�yP����Sф����������9(�+-O4T~�-n��S�6�d�ZN�������ۍ5W^͛_��Bf~��O�6�h�U���A�����o `�sd�z����&��bF�nPi.�2�Zf�u���TLp�{��M(G5��rs��@���'�}C~��Ľ�|���l�>���8��_#�Q2�,�B�f	)�����2pQz����� � �q؏z�d�?b��\R2 �F��)O��M��o6;���rp��2��;c�Ưg�vyZEK�2�K��+�=�L_iZ[0���JX�LU7M~M����F<o�ɍ�m�h=1�S<�� w�fL�Y��6t��ۅ��z��K�&x�U��9�k;�3pR( �5�s��r�6���W��m�D�����K�C*<���nG<�C�.����
�T�/5���A�Y�eH���iEC�K��dp�?_B�/t0�E��!�r5l�ۋNV�N���|�{#�*E���Oh=���:�KU(������.����ы�ٝ�ُ5���z�����n���5i�G���j_��X� 6BQn��+�{C1���>��}rP}��
��|�.R@�؈C�M��� ��t�����<)ר�Ά�s ���U0!�M��k� �����~+O��y}�>�s�Uwr8<�k�g@���m˯E�*t�|.���/�f����ۅ�M�^!���E�����������H�&�c��1��8DzcJ��\��"�)*H˪��g�佂���E�7�l�OQ��X������$gہ�w"��T�i�P����E-̢��(��h���'*Uv[�n`9�,�� ʀ�!�X��#I�O����_��_�`
`u0����5&S|~��~��c�<C<�B~��I{�N���v$�C_�xP��B9����HE#�E8C��S��R��XKg��zڧ�V�U�=V'�r����L�Dd����@͚/�&~�U������g����Ϩ�m�?c^q���U��`��S]�M�t#�i@��.@cB�%XZ����T�Sy�I,<
L D�?�S?k}���`�N+A�G��X-��O��R���TrM#�ړN��+5�����`U񉺟�V��e�}��k����y⫂��P�^�r���y������
���sF�����R�����X�`I�y����A���7�������E���SvE�b�l**T�v��W�6���h��"���ؠ��PB�{!J�u�|�t+�ӟ�b5g/2Z���<��yE�}gЯi��-���X��]͵|�^]���%�҇e�1�Ϡ`Zӈk���1��c0�Smv/Q�d���r�A]�vj��#��g��_^ds�s�s.�b�~��j]��!T&SJ���Yi^��1����ff���ʢ�l��f��Eu�Á�N�,iB��)ڿ��\���l�&�g6W�E66�#�0l���..��A+Z��fSD��P�Lfo8��
��w���D2�}���b�Rdm)���4�1���;ڭ�Ԛ�T���IM�d��,L�A�*��0+��t��D�cZ��/YV�
5�v0��*�������M㕯�m�R),���-j��A,��4b�M�~#7�/3����J�U*o��6fϋ:P4�ZT�� r��<S���X�� �C�Ԫ��ho�+�'w�e���SԤ��9��f}^��Կ�1gE�-�%H�;��ii�����$7���%��  ���b���&�d�b #4I��"��a{����	bU[�{�{V�\J�yڏ5�=U���DZ�Am�`H�C� T�<B�f��Mvi`cepuyy!�7�2x�AU�nު�{�����9:�M!��x�-�m`wp�j��� +ԥڬ�`��[�&���C�?�9�,u�˫A6�[�z~-�O��Z�@k{�����̾ �B���g��딁�[�g�@ڇ4ZA��U�j#��7�
�����
��*H\�y9>�N7K���
T����	�%0�����٘}�q@�-�yy}D����dqM�;4��>B�s, ���H8u�R�:P��c�loa`���=�������T1ԇK�j�D4���]��b�?�����fu�_��߲�����Ͽ��˛�u��J�2_PLU(������'�����<���l��m�6�j�AI��Q�֎��=���
�zG�WFe�^J�L�Q�yTN�՞��VE/������fn�b!ى��fBUY/�U)*�Q�������]���1��ӧ;��׿�/�U>�~f�Y�6�n�>A5���i����k����-g)���H*�Z"*�H ar�g��`�՚����߫MJ�*c� 0����c� �?����2=�����	�f��&
��ZN�N-�1yJ�r�.��0k.�[�\9 �/����*��3x����]-��XZS�T�:��`dߨkkd2uƱQBQ�G���&���Y5(AI��� �'��V�:S!�Ȓَ�ɝ�L�P���i����A2FCɔ#1�{e&
;(_M�P!�T຺���~x+?|�J6�/������,��L�U�����/}��k�I���ܮ]!�5�t7��!>!uOyّ���QK������V�O�"�#<;� ���F�kPY]�͆9c��?(*]�J�3ke+4S:��x��[-�{ÊI���w�������H4���P��P��HG��_B�ѕfE�H8�����Gc1�JB��LoG&�@�xa	<d`Ú�4����	�gPON��:����
�*6�XIE�0�|�I�V�`%�3HA|�9�w����jR�O�
0K�m1gΏ�~)�fFc�5��+1�E�����5��1��[q���xz%5���ؚ�L�3��=O#յ]�0�N�vQ
gݥgM�A�k0�&�]2:�OW�"J��OP'�����oP�f�P��m�B9\*�qH�L���9^��og�PU�L��쬥�Iz+;�F�6КV�l� Q��
�L�����{L�A������gy��A>����d��9JJM��ڣ7����SJ�A}q��=|$�G�ώ���B��fz��X]��W�C#�
DP���������2�@��T)\s�X��x��-/.��~/7\]e`�����X�\A�a�Su�y%�Ug�GuF7&�M�bsy�>�o��%�^y��R�f��gރ���Z�QTes��sYe �*ۚ�|-�e�� >��q����<�N���Ŏ=�P<����b�c���H�Ԓ
�����_}�/�Ɨ@�׼XV^F;�9�@��\gm����O����9� �pus���l��)R!T����:`��F��̲OETt�Q�� �j�����{7�{�ƻ�o��G��֜��{B��[�JK�����(��d�s�{���_��?�7�������?������o��H���?��������Rmຼ�����A$�{����X,�@�
Y�$�i��O�N��N�2h<1���h#f4�7�8��e�禯f���(�Eb�'��72(DV2p%��G����6�����u����Ї�����Ó|��I��KY�d���6�I�5�jb������.iV{��[Jf�x���T'��+�=Dj.�b/m�el(��z�EY��\����W��5)N�r���  Cu����06�/�T��v��=��SE9&��'��]/�;�8ʹ���҂�Z�/��?�`B*n�=�c����6���O��JJ�6kRj/�d��K���mU���Ś	�c�-[(y����Y�%�PE�z�u�$�e~��kХW�:;Y=�����Y�O�v�>�\7����.<�a�XA� [Rl ������(�;ZņX�IY��4�VR�j�O��k�o/����bA����ԑA���w���i.�?)g���{Vm$�XC/oh�H:���R� Y�a+��XI	�T��$ER�d����ہ��y�V-�j�~
J�@&Q���/�G.����@U�qLf@u�GH��t�&���+ )�d K�eJ��9S��i'y�^��/��b�F���Mz��M��a�7�փ�3��:�
R�
#2�%%��u60��XI����)�].�����J���R���o�!s[hu�ߨ/��U�(Љ�V���wN���p�U��Ԕ�)�K�������n]�g[ i�>�k�ۘ�����;���Q�u����#=�չa��	Z���=���C��ӧOr{{���iw���z�L%�^��r�<�ׁ�1�l,��p�:�W�Cl����B.�y�v:����i�������#E>}|'����"P$�1 ����{�|�����H�R�
Hl#Ղ�w��r�*%M`A��m9��9��_	U0�Zc�K��yGܪ^��7�r��;����e�u�m؜��*�k�/,����Ai8�݈��Nщu�O2�5��Y�k(~�/�*]7|]-z%��(~�qvT�-󵬖ײ�_�|���#��I��0.�u�/9+)��-i?��>������}|��k�*F=���i��#�
2@�&�LȡG�������$�7�k��X�ģ����1��m~�#f&�L�p�^6��͆ؚ,a�A�фA:�Ai'��U���S�S	�Hv�)�ʘI�]�>�y��6Ù0b��l�޽'��o�`�Wҁ�?���\pf�J~��'
��W���Ϝ����8wQ�P�Q�KS���ZI��b!yk�5 �j��O��R���|9s	fO���k����R�V��BnPڻ�5��cCfG�];�{�~8e���7ky��F�l#�uɟ����3�����C�1�s���z��G��vH�&��1�.�^%���Gk|hLRAK~N�U9٠a�a����������|Tq!�H��T�XWPs.���j�Q��Km�P�#2���Y���i-�yS=#Iy|��km���--.�V���F�q�T�ؙ�h���0���&�� UO��Ks�=|v��^(u��z�ĕ����d��,}�rC���� ��iO����1*F����k�{s��)�z�)i<5��b��$I%�O,��l>43F���\���|��#��>��<�
)�<gc:g�/w�<YS3�m��N��&�ܦ�[�<l�V_��W��׶��N���u~#e�s�1;QmJEp ��#��S��u��4O�!��@)��b�Ҝ����Zv�*���:-Y����0 ����W�����h�S*p���\��%U�p a��Ň
����`ٴ@��r9��v!��S��+W0���� xh$��t5��N4"�c>^�ϴ���*,����avI��2�'XG��)�2m"P���<6�d%@Ue>�H_��4��F�-��l����@�eɢѾ&1���Wߢ0�ѝ�����9^Uh�W��`���d)�.����fcHM��sL� �_�*�P�R�x�h��5�
���@r���^�
eU�v�dJl�PA�7��<�
U���d��>΁�=չ���U9��g��cs���a���6���{(�b�@;R�ss�e�7�~,T�U(cNp�s��>���nw��|�@�,�8���mA��u������>�֮	)-��:��p5M[;�fK��@u$hJ�g��x��$��ZpT�����|@����\��^��A�^����F��W9���o�^�Y�);z��(�5Bz]���j���`���KWy^�����H���j���{'�q��1��DK9m�@����s� �sY}Xf@=���L�k���O��5g����z�~�F��<Z�%/@y��+q��{ž��B���_�8H��N~���ޒ�f�M�`����6/�;�����\���7�Q�ϣ%_�C�0������`�,Va����@M����b���J��[_�����mWL�;����I>潌c���#+Z�����߽{����;D�s}}���L~ƾ�>TB�G���28����V죉`�X�Fdy��JA��	i`����q�@k;�4)&z]�Lj�WO{Ԫ��H�l$�י��@�,�gf���wѮ�]]*��ʀ����\p�D��oP�;�r���~ѓ�9a��c�}�:�C�[��9�H�ux�`{�$����R_��#cW˂��oA�����1����KN[� l���s���k�������6��7f�xP]}��;����E�g>�z|�Otfjp���U��l���*�"eߪ����P_)��_/d�D�'����_J�'���h��Q<���r鼏���ݨU��ϴE�Za���Ó|�}����%��U�U\�~Jip���,���1-٩ �ɻI�S��5]�d���Cu�E5N���$�|��̰A�$Á�g��as-di&��h�?��ҥJ�>��h���p~�X ���������u����M���D�0㌍a����F�}6zM�g�W���@
�5�T��)��?�q{zz����l�/I�]a>���Î�j����|0����z!���z�Vˎ�Ȟ��(�~x��P�2�$t�h���\��\�����#Yf�W�5A~�?�)���!oT1:��6�)E�3rm�nP$C����D�7扠��`�,�k�K��dph��@��P#8��kZ��ؚr��v%N}}rݦ��Tث�g�"6�UA�{���2�����5��]({�A)`砫��qS��(3}}Ǹ�L��ˠ��M���=Bl`�Ji�O���)M,a���H���6�jҿ{<�	���%�T��p��=��&�,�h����±Y��כ� ��Λ��,�^d�5����%���ϋU�^�#�r�^d{A� ��wj� .��w�Y>��+%�W���s������+�0��]9_�_"�����%V�j�٧k�Z�y��e�J�����e�cN����X]����o�u0_��!��K�:q��ҝ��:$k�w_ J9��!G�4pU����/��<fhc�󫘤����!�8H��ݕ/�QQ2X��8�5�9�zp��=�$��6����~w⌿�˽�2��w2����*��A�J�~�}�+��0��]L�:���[۟��rnٻ�3�>:eĄJ�&Sc`u{fs�A��J�5��~?���dFԄ̐4!���Ez����4a��R��q��ڵ��\	�$����_+xf~ɠUL	5�������GV�o/?��\�8r0wwK����G��p4�M�󾸺�K�����3�ݯ�ʿ��_9����wx,E� �ם��)LB�~�鸒�}��&�������9i�'�q�2ִS��I6*v4}�k�=���}��Ԑ
�
�h,}���@$.k�����p�_ҙ�$U��A� ��"F���m�o�R��D�xܫ��JR��f��dL	��8�y]%ј��F���,2�B�v)��z�يf�|�'7]�D�q9 �}�k���j����
��~ε4�7b��(�#����=�gC8x*�/�&�I��48�b"g�ّ7���R��߲W�
\�ȯq���V,���5�%z��ﰾ8�ߞ �j�����}96�9x�0�/؏H}	M��~�E�Ϲ�"�hZ5��BM&g��&�!�]d��U��#�ѥN,��7d4/ː�MD�.,��μdZ��Ue�f�9~ڿ��<YiP�xy��|՟���0�\Q�iJI:5%zd];��GFR����gñe5K��^#ƪjSɪ[�֞��w�����NN>p�fY���ƫK���\-�l;[9O���Y-h�a�T�=��>�Gn}�� 
�����A�xBv6��f�D3~sd43��|���EYK�s�3�B�P�|l Y:9;�*E�Ml�xÁO�;D�yLt��5'�*p��ט�r<�lކ�dֻCaYp8 V��d�]3�>���^�i��;^��_�S'�� �A��r��kq���F�r(�w�gj�R���~%[�E�x:��/�7۽�$gΎS*H+�2YܫTΟ�!�k4����z�
�|���u����C��,��fƤ�~Hf#{<Y`1`�Wσ0s>�(�Q=EQK�$�S�=��;�D ����=�TB=�ؼ������J��ý|� ���F��U����Ev<Hr�%}�L�ݚ��X�fJ�*5һ'jo�_oi!u&��c���@힞Y=��i3��a���E�Sz�Jo�Od}/닍��F0�W�!���y	�@��wG��SRI���9��zp
Ò�����c��D:[���Z��YJ�dv={KJ4vK�B�@�|/�4$�����g)��UAx����Y?���1vL:�tѫ�Ӿy�{y��˶�d�����w?Z'xn˒Wx�U6R�>�yػ^��lX��}�u[����I���&������&�^h��b/��s�Z�S�������d��=��<P�61c@)sZ��q5@eu�G�')���,�WH�:����{w��1��I~���/��*.�����a2�����>�O��0�p���kA4K�����b� ��b��j���T�U��U�e�h~�ޕ�,��d��jH��`r��g0�W��o2��Ą�1�\u�L�I�,�U��~Gm3`E�	fL� �fd���]a@��.�&�/W�d@�1|��R̄��O�"Ȅ��R�VRl-X�,eb�'�S�s&��;Y����P�t�|�� %	J�m�S���곝�vZ�Fo���o2x����8fۼ��c�~�P>�Z�tҙ:q�����J���֊��vș�v�ҎZJ�/)���5r��ߡ�Z��w�̔ټZdln-�І-?o�;p�Cw �0�g��p=�QNZ���h�2��7C)�ܞ^���D-��,��¢Mѽ) �B����UL��� t�TDa�ϕ�,�j�s�D��Au+��_
ZR�8*����JA3�(M�������NU��9,Y{�L�ڰ�=�*�̊�7�O�~
�d2�/�x����>�B���MC�{�Z�\������m@|o,~h��y��=VH�@�p?[���e�����Er:�Ϸw�� [�J.VT)B~vs�3c��b���5�E@��9>��ax��!�� _��g�+��f��98ڮ�ˆ�Ǔ��3���_�ͫ+���wrs�*��L�jQe�g1�Ȑߏ�ک���+/3��\=��Σ���Ơ" ��D�'6A֞�\	��sJ��'P����n�)���V\1�k6O��o.��k�<�<�Od9�hbg��ф��}z���U���`������.�I:s8��M������>n����x�w�fa�T�Ē>���oJ	8?\�:^$k��AU��W�yW��m}�-���[2S�D�	������t&S���f�I9�"7V	*N��,�8����HT���_�F�����zs�A�qv����[I����%�S2�읊�u��.�0��z��a\e<�:į7Aym�񐃂������m$$`'���@HH���r��W���t�5�&����h�&�9�v�?)|q��y�~�P�7+i����&�bi� A��̲��|Yy���C���g���}YO�0��=�,>����r������Or�ݏҡ�+=u��*tѵ�
���r�]��c��<s���|�ɂ
-���"V&c�S�o�K��bm�|��m0����=��Q��{���;I�$?�������@��L@��p5e[|��h�す�`�w~�/A��Ͼ�pm���e�jJ�\�W%_ς�SⶇǼ߶�p%�C�ῇݎ�E2�7���mT9��L����I-�Zur����&�t���qO�F'ײ�� ��rMp/��s�k�%Ϟl�i��ݤնd�M�O�߃~�h���?�>v�%tR*�����Y��=˳у{��G�����vO��XL�`vq���μ{VE�-N���;Ua�� �R�C��@�z��pi�bp�<��|b��s -*�Q�� �7�c��	q�WZ|/��U�mg�,.��v���>0QB������R|��ɰ�D��<�&��Ã��x���L.��pk٬1��U�6����g��T�=�Ns�FI�x%_�QtP:�d�@�s�0�#�e[��l)�vTG��4y �ȶ�vY��yp-�!F�̶��@��J��iLZqŸh��R��՛��*jo|@�U�(VPӔ�h�9��33@��)�ϲ�}��L�6KΡ������r�ީ���KZ�H�B'c$�J��Ē�-�¥ ^m�'��%��)�1c�\|�c~Oj��'����Ɋ�T_6.�/^�=q�>!ٕ�'F�l_����6*V�Ǆ�9���o��:T*d2��~��TT�W�3�g[����>grnL�����(����z���{�y4����2��4��$�����DR�,K�SСΠI�{�^�v���+2���W�ꉆ�X�t�s�sM%���YUያ�O�h��Oonk��)�īKfN ɒ%d��s��\շF���x�H�`=;в6i��^A���@���;���2���6���R��̭�Fi4��C6���@-\�\\9�"�k���`�F���k��ܑ�2�w�]b6��R�o0���lf�l��d<wux#�wd�j��Rmr�)�LIXx
t�0�l�� p|td��[�X՗P-#%5Vj����m����va��\����	q�SB�d��N�򳺬�J�-��unOO(�|�"DK����H�ϕ/>�~��/�q������>���g ���g\�"�:_��;eEZ�`W7�c���z>2�c�����5�ʪSQP@����+��]l,C3\=I��Yr�=�fƵ�$Z��*h��:T���f��I҄ �)^�"+�����?�@����,���k�՛�l�����h�{���J���&���"�^�=����u�u)��xO�����V��s l�x0>S�=��VA1����A~�����SSi"hHJ�����\BS�mm���k+�[_����G���\J�X��(�_��a]�w���O������ѱ�?#�z�ZSݵ�;������\�P2�g�.�m��/f��RE�x�����g05:O��N�#��p���s��T�����2�����7q�KdBf��r�d�Č�O$S�^��׏?T�.M����`��z4p���M���k׹�U����|�}��(�R���C���%�B�yt~!T���2.��&5��j~��X���D{�&����=o��0��+�Ga��x@�-�aT��5X�$��.5qNR�z��E�^�DFT�A�O;���4V���\n;%_k����3��\�TX31��s��U�Tv(����j�1����0N  �Yݲ�+Z"Ľ7�UD�S�Iw�w�k��O��۠�Ay[Z�3$�g�����S�L��.�ߨ�A��	��$�� �[Mؓ���R���0_(C(_/�?J�wr���C��k�A�xP��}eg��m�
U�1��)�#7[��N5�v��n�S\}I�|i�ڀ��<�&9��}��:c��\⎀30γ?�sb��#[��q��oz|�՟�X
)�G��U�t�_5����)yi�T��� 8}�f�iQe�0&���i��=U�bW��+���׫)2^c�A�SS���~p��e3�$�a��'Ԉ$s�"ݐ%/{�SY�R�V`�[�ݛk[�R�ŧr��h�D��Q���s!�k�f�ݔQh����\�>U�P�B�e��R�PMQ��)� h���(�]$Mpq���
�a��-�Y�d�����bN�
�֤��SY@���>�5h�����Aއ����׬b�W��D�șU�^�R��X��6���=ۑ�$Nz ��HLPH�v������D�EJ����ѨE�R�핓\:8�� @꿭���B/E��-gI�S]^/�,h�7�����~�}��"��� ˏ�y؇y�\q髁�W��rh��es��o��*�/)��JC��fh��3^;��E���N��\{��ݮd�H5�@��	�ivy��Oe��܀n���lƷ�B K�us%�͚�5p��;c�$q!!I�􁨌n���`�����eT�cW�5�b�
e�%]�\+}��S���nYu�-Ǟ���|<ˋ�*�d�;X�$�t��!��k�K&���{W��i��50��e�����??g獤�.�g�m�8Ja������������uX���EL��K��I��,�������o�~��?��~�~��P��5cE�r�Zg�Q�c&�'W+������J.�}� mP����Q�-[��<�&uΘ���!T�8Hwڸ��	.�Ӎ �	Ca��ѻ�`Pq
�-���;�����C�AI����N:D}�C�l���\����3�Hy��ަաڣe�LAUU�F�s��8����|����y{EȭP�ER=�n������k�IhP�5�4g ��:���ʓ�.gҤj�-fs��Xv��b��~su-y��x|����(�?|���&^U�Z�i�2H�ڠ�M�� H���Ov�_b%�#{�Qt�N$ڃ�?Z��$~|F�G��ķ�^@rvMU�^�3X���SZ�x�%��F�ؤ�U`sC����&s<�a�,�xN4YQ�f��jc4Q+�HȞr\p�ʠae��gmP�-��w���a���{_�LQTX���3�$����3URb|�?UA�X��(�!�@�q���V�'��9}΂k
Oj@�3\��� �?��Q��I��G}_��\��QC������<�\&��SJ�����Xc��&0�
���c�������)(�TP�����;T��b;P�#�ss�x��>E�/gc�i|H�*��礪*���z.q� ��U˿�?_�ԗ��W�R���&���@�O�?�_��CK�$9T3��I�tWO� ����?e߻�f�Y�J���LDU�<�j���]����̊��p77SSQ��ٹ9z��i7�4�1���58۰�	>$[�^ߌ
��5��Ɇ��G�I%���c��N�ߒ�JHV��E7�~�;��5C#<_�ed��U���f�✙,4��� ���.G��٢��`��hNI�7�Ѣn����s�*���C�A��./���%�bd����Z�#6�F�lBp�\��(�% j�9�����������ߏFī�\_]�	IQ|#M�u�g3?�>)m��-:�93Xl�ר��-��
� �[FL��#��񈔼�س����F�ݞ2��É��>��9D���@���"��>K�́LF0��O_K�NY��("�N]�^���`�(��?nМ*XO�
'X�qz�������O
���b7
�+��Zf��Ҏ���j)܄��b�sb����յ�E�!�x�dgߍ��:���/�"��3�'?�3 Z��KFI���� Fu��E��T�˩�^\���6*]�"�3�9r�j�ؓ����
��`�_f�l�7H�	�tk���������\Œ@�HZKM�j|�K���G�:O焍�F�5��=y-B����<����xO�.�8�y#�������+������[�z��,.	Nv�瓯n���:�4;�=�@�_{�����1«���q7<@朜���I�}��&�xzu�\^�|E���הs7zr��}|�E����N)��p �ެ2�y��:��%��&�̲/X��׽9���s���
'�h= VT�1��,�W�`�-�i���3�&6�?1�"N�n�����`�S��4�7���7�7�Y`"8��W��W�����7���Y�!-J=�����O��i,s��/p��a�m�k�ߴW�Nm;�R�!��F�u�˼'é?����h�p�߼}���吏�Π7�w���A����=6�3F�e��Ok�$�y���4XFl0GxP���ǝh2`P�m���mѾyS�f5����?ȇ9~��p�O^T�3 2�%C�_�(��OGf��@VҜ��s4,=Q�@���^��jZ{�u{���TB��Vi���$m̀[��D����G��뒶*�Xk1���'�UG����D���+�Σ!죳�}������!�+E��_��9��%@�~���W������ ��>�K�O+����b`�"� kPN�i���i�2�ӖL��c�l��T�X��P>_)���,Z*Ƣsӣ�x	�s�9!��9U)����	+�,W��_��Y�!M�zҞ��� ^G�o��`i}�������߰�6�3:�P_�Z���٥,�+F�P��S�>��F1&&D4"��&�F�i*j�4������݀�7�/���\�q��t�>�L��1ԉz�M��w�9���Wx�~����}kc;e�� d��d}3�����)h��'W��:�v��ǄH�6�H�1���Ӊ>UЃa�ltgT�S�l)ރ,�J7��A|�C��N�X!�\X��y��ח����Ռ�=Ң�),Z�2��֥�u$ )�o�?��	��yc�F6#<`�j��?,op�\��3��=� �7b�Q0���D& ����������>)u+?X>A�H�}:�-�M9`�OV����Oʱ�)Ԑ8⪫�[#���K%rX�27lȦ��9�͏$UiptY��8G�6Č���yL��R(�,ܜ�U�^蛓f���$����6��6��~2pf����勯�甁,U,<0�Lr�^����Y�S�%��2QO�4��SDߧ�%�r'ބh� H{��m��{ˈ1�C��*U��_�n��z�N�˓11f?�t�ui-�ԡ�w#��>�:K��wn��z�Q$m�T_�y�����ڑo_��7r�?j�C��ͽ��ʠkC@���W��?�y����E[��E�CӼ&�K8_��h���|1����8.��ّ���������F������|�Z,K>�`
�-��1��]�;2U3:/�����>{�U�[�5�����Y��m�l�ײ�Ju����n����O�y�c롍�SLki�ÞȀ���g�Qp����#���܆(�4�����y'K�Ox��R�3*h*vR�~���)m� �A�W}g�{#��V�h����QmH�pncoC_�������Y��l)3Г�0���m�efcA)d�,��.8����#[��AW�+���i�	�O�VϗKf8�#T��k7�����[f}4c@�K0�ϖ�@L0:z	�"����5�1zVp�x��x�R�!�`~pz�f��R����拙�ǜh� jn��?����b��!K�Hk�
1�C�����&�Nb�v�s�(V��u`��5����y��!x�$�y�f|����`%U�N3�ؗP� ��v������;ƶ��	��|Q�1A3|��ՙ�.��ޑ=޲UX �=e�;��1P,7a��ľG�z����`R��짣��.2<s�ֽ�_1���{x�9��,)�H�1Bе�l=�xJ�ɛ��qvZ<�~)�����3ڈz,��){��ϓ��9=p��ܒ��
<�4�ͨqS��	��@����ږ�~��N�fQ����s�K�.1*�Ef�R����.Ι���uP�8Y$�Nn��af�r�!Z�e�{k�Ձb�P�2�vX��Q����Hu�o��3uPd�W�Nǳ�%��8v� )�'���,V -�O��4��0\G��9jC�õUB_R�x�-f�g�AT�c6>�g��4Ȣ� (6�BW��6}�,�\�)Jl���(%��Y0����r������|Eu����KÊ�¾U�.���nyo�{<{D�w�f���w �ǐ���T��w�M�����o���r�5�!J�,t�~P~z�:����) �,1�p4e"�H�i�OM�_�N�/�t�ӯ8c0�	�/?��O�kQ��-yr-�1���2o~�A�N����q:���vk���`�0�k�42���]�5ևvD&��A#�6���9Cqa��n�!;� �LP+��J��T%H) ��.j_9|�w51��M���,�lF4B�9����6�Q�E��Z��m��P�&�ڵ��]߳5//�N2?���S����)�jm\x��v
FWKc��1����$Snk�����ɻw��O��9�~à
V�c>�7o~�ۛ�l��Ջ�巿�g��o�YΟ����LP�6XfrˉOw&}>%�N�j䆿1��������ĩ�㓭N��ƜYu}M��s5�M\�5�q52Z�9An���g|��}�*{LQMuH�;��f&`������e��"d34��R!Ԃ�*��lˎ�:Ps�"��b�kQ�Q�c���0o��ɚ��"I]��diF�3à�d�P�BԑP�O*��۬���0��'��5�U��2`|@9���`}.v�
v�f��`JB�D�C��C���ޟ��n��;ᇨ֠5ǰi�S2�{������ƲaZ'��e�N?Me���k���]Q�'2J�,�����/����4{Ɇ�������fͰ�wV� �A���[��?@��l��}&�ϲ���`�h��Y��E����ㆽ�0@Yl�C6���_���/��-nt������6�53�]��l�T��ʞ����Ȗ�s֧�����<&2��N��:ou�R��0�w~���/_�����y���l��-j]m��j�= /��G4x�NY�~u��Ky���;RQ��w@O�hkQ�ɭ�	���rZ�v��2H,v7��[z$��:~��P���AjK�ﱌ`�V=W�߈��y��V�,�g�fy�MT�c�\hA(�����K=0����Q���X����E�����g��E��h���]`,t�0���x��7Vk�!"�������Tx4>vS�-,�9h�(f=�!*4~��Aտ!��Q-�!/r�~�T�#>b�[�|]E~%b��� �4Z�l�sn�6�,�����IЭ�[��T�.7��ߔ{;L�H�^q_a�	�}�xK'j0�� �3�r��ln^m6P��`�I6�,7G�l �qȋx�&��7�x"�닂�,�=v��N������|5�j�9w:��Lv���������B�4�~"&���g$PN�5p�z<�h�hY�0h�-����,u���}L���c$5�'[�k��w�KCsi����!�G�Ny��cU��egC������H�9��d�u}I}LA��:�&xD��,�3���ذ'b�"]Dj��KB?��c��;:g�����k��3+�v���s�BJӳ��m�F�q<�?kU��C���Y?}���Q��@��AOb����M|��0h&0���7 �<wE�	����6�h:v�H�!y0Jx ���L�vr��%hs��v�qKr#�w7�yx`q=�c���1;��)n�����޺�\_'t)�[z�q���'���'y��Or��@�ԡ�a+�>}�O�?�=m./^}+���?�/�9�|��5��:�������P���ts5`R��AF����ܰ��C��G�����~	�^�����S��,=���l��L�K!�@�
�����y��k-JXZ'��8�۸ Ƞ���Zn?��O߲6�+�}c+}��}J��21J��Ƭ���Qk��`;۳���[�,��@k��ǁt8-��g�YK�����j�
��9� "��\#��)�%T�ԓ�r��L�z�T��-��Mk�&���b�b1
z��D��SĜ�Q4�yM����荈M� �3������CG�<<HԞH��G���¤xT ��~��<yMU
�^Kb�+Hd���i8�d$��8=��E�8��%UXD�Kġрy�Z|༎��עw�j!_�L��O�����F�Md|�����Y+n��7y~~P@��>g_����D^~u%���7���E��6>�"�C���7�(6� ���eK�.�}��?A��7���'7��n�o���z��q��e���>RP���<z�����������J �hX���{����y��5�d��H��?� �]]�_��噼��y�ꕜ��dM�G�H1��uJk�{�L��R�R�F,l1Z��;
��d�k�2_;4)�
�ym��d�Wt��}�*F�� �
���@�R����IZښ�U0Tʝ��sN3sU#·C|W[�_I�ZiԃJ��U� _^��FP���h�q�Q���{Fl�d�Z��=oD3UQ�8�!BD����*�|`��.�
����S��f�m1+��i��%��ݥ��Q����i�S��uk"����t�����L�|��1�?�P:Z�}�Z-D��y!t�1uJ�
�t�X�ʸ��(���4s��t�8p��84Kг
u[�)�'����i^P~�S݈����G>7�GF��W�FO�t��U�`Qaݞ6]-�>7�#xUt(��j̛��U�~��By���F�Y�������cgu)�
'@�l�����ӳl�W*�ުL�`�������,g�?6��鍖Z=�t.�P�j�}Q�����O_�ZJ<A���ou��|a�:h����2Z��P�F9�
�j0g�{0��PA(z Ĉf�K��F(���h꽥�-��uE������Y*��Hn{P
ihvM�K�+C��ޔ+w��F�����Y23gL��Y
E�£u�3���}x`1#�l\vnv�Gك"�D݁�<�Ӯ%u#�	5IJˇI�͢�n�Z����n��!��ȯ���w�`����`�r&Uά�C�'ɺ�9��6��|������r��}�STo�h�]�����A�ׂ�V�_�B~���_�����7�z�y̵w�*?�-��>��|���/_�9~���j��{@�S06B�_:Zq8���l���I{��%����I��Pc�vo�,r�~���f�\*گk�Ufg;y��G����l�w�v��XoG�:�z�,b�"�EU�H�4�����1ѹզӉ��{�!�p� �͚̐EY�Rw���r��:��:^?�Vs��8ԥ���<6�#0�U�m�hjm�Hl��O�5-�Q{7�����n�l��hK�*�5��҇��B�Ehd���Fʚ-Þ��4�i��_�ǋt>\�j�5��
j�o�M�p�Aw�����	@z�;k5���T~\��pN�����*����ݑh�PMQ_vqy���Y�$���/g��/���9�7�x���{��P���k��Ƿ��=\ʧ��<g*�6��h.��d]˫o^��5Tg�ƦJ�����ϭ���#�.ϗrq�"�B���{P��@��L��a���aK`۸���{�@�m	�Ha�h///�׿�k���xN6��Wd=��|��g�������1��I\�b���%Ye��<�yi�`�A	�[DW���kO�t�׻Q����7��u�c%�F�.H�Wс���2iſ�G�S�Ϛ� �mk�&���d�:�[�u\��5���Z�5�� ު��2Y`��t	�|��������"��,��8��g�'k�' uJU�6�c��h�{��k��-[���,�S/ܡjh��L�t2��Dٟ���4V�U�V8��_~���o�������@Vp9L��������:�>�M>������fo4����,�$�и�`�(([�$�'�D�*�/���90�&��z�=��?���J�P�;t40�%��U%1ou4�M�kE͸������ �z+H�L��q���L4�Z���E�9k��~�lV"�����N�|�A�"��9��+ʫ6�Ri��*H���P��>�GY���ѬH��<��B��~(|:8�\i�d���y�A��0ٹ����=p�'��z�1VrI��el!"z8h}R��8�s�Þ�)�1�\��.���:��d���Q�.��46,<�I�i�K��E���{����
Q��f��b�	��z���P<f Y맒�w�����kX�$�H��}�ǈG����xO�Ú�9�V~dr�kkא�<>l�����|%ϟe��:�h4�\ǁ5���駴�p�v;Y������������Oy�w��X�f��y ����x����~/����l}+qz���6��0��vu7_'㚷ҜM�����4���ƻ�����S��nں���j��͔곚s�1H9fP_\�K�t�����]���ʙ��E�FC������?}/7��g �����������̋�6����(<�Z���vMTy�H��R�{)�>d-�m�9�z�}k��GjT����41�M��y6$���-�se��&&�,,{) ԳJ��>0�����eï��q����\����P#���As��~���c�Ǥ��l�+��c��@�]}rV�^#k��b~��O	�m�&� &�����T�hcRA���ub�*x�BgHCFe��_�����V��M2P8���:Xf@��c;?��5����7/20�f�����' ��
������<�`�c�Zh�q��q�m���Ys+,2��G��?���g1�|9���2_��[;����Old�� �>���:��`�Jeǽ��
 +�fp�����󽺒�U�eE�9}���R^m{��᜸���q�(�2�im#)�G����B�K��t���(6�D
�R���=�U�S^gq�E�m\}�3+����(O�q���O�ʗ��hBy��^X:��C`Y3�E[�<^�쵿���K���i�v�pk
��k=��>1Z�:X���#.�ɛ��i�+<��3��gSЩ:>�;*�ә
���15���2��zsȇLE�ރzS����U�uz�N��)6s����Hz�<�F�?��)H��5D�&�����i�ηo<@gz嘓b�8�P%Fob���~F���tÉhfǮ��
a�`7��Lb��8���FtF6t��f�D9� Y�ȸ�m4��E�]���Y��W��7֏#o�a�f:�0��z�~O����83jƛg��|�&�>l�x�3D0�>d�j��&�
XS�C�h"=��OOg�)s������3��c#�j?LŇ��=p�U�ln�ѻ��l���\M�۵�z��7�qg�'Ч�XR�Ը�o��:���"���TJ��'2�j��:O���)�j �<{�Um2�8���һ� � �π�aZ��.�2���uټF��Y
�h���?��4#J(6�L�YPg�7;��>�#M�9l��7[�������#p��G4!���?ɫ�|���`y:_�:������ڰ�]�4�5>��4���r��묶����sݭV�;���yxP������򗿑o~�ٹ�ZZ�`i�c��am@�,�EK}���~j�Ւ�z���G����ӝ��_|_R�=��pb��*���F	@�w��f�Nxe�F�T����o^,"<����6l��o_��wod�x���V����]���qG��R���m��O�Y�f�� NL2v�JX�[;6�F��e) �$�)�{�c���Q��3VG�s˝E<�6�WFL�kјE�\��])�σ�7��d�������RyM5�@j��X%�Td V��3:�B��z���IUlK:m7��l{P�ۇ�{ڧV�,��%җ]V��R����yv*���jk�ط2h��h��_�=^�5��8P�=�8�-�y!�sv~.��_�GY�&�2�f���_r�dx̊\q�Rk������l�	(d�Y�X. �����i���W���Ōn��`Ϛ��݃�s�ɠ^v׶���^�6EQ����t
����W�4@8� �Y{�A�����Zo��[8��lB���A�hGU�N}(�'��ש��,�����1�Khs�V��>����Ģ������85I�40�k��@07�mX�����뇒y+u4R�U�Y�c@!�ڶ�s�j@��b��,
\��C&ݛ�`�݄*h/鬫MmR0�6p�t��a%х���L�7�|�L���6eA��
Zm��˩Pm�l�l����`�Y�t��K�&E��}H���XP�B�:2�ɂ��`܁��P�$)!���wc��6�{�ɬ9��:�{���k]���?�i��$��qha��'JO$���*ܰ	�;��P�we��� �d+q�����jjMͣ�6;9����:߬�*����ک�u@Y�
4�܈�.�Zj�Z�BFy�Ӆj��@�=�GfzR ���h��d',�:X�B6��Ns�/[����D�M�c�w1!M!d��nJ
)�P�W;DJ�j���f �y�ٳ�4�򦲀J��U�b!H���9���+i���+����ct0~.�3y�=7�
Ȱ C*�S��Hʉ��G�����A#VL�4�R��*Q�Կ�2/�Vc7������8[�N��Q����۪PM��R��u�S�68�%Hi-�!�HXKiTݯu}ɨ�[������pT'��u]d��<;��7tgOF�������=K�MU��ȉ��oF	�h��,2U��7���[y��k��6>[���"6} -$�sn��
��P��u��O��q0E<�wi��Y+y����������2��f�	]��G�E�wQ��˛�2;�S����>��Qg3A4:;��Z&qi4^(��2�D��x� ���ݟ�;i#��Q�������|�+:9-��-����P6��kf�S>j��&T�f�qS�����&��4LV����+��?��<������6�3�8����ȍ�Ӊ��2'E���siZ�u%����s0��#M���}�����3d3���Q�p �:*ZO�k�i���J���H�ebpjs�Hm���"�)WzT�����d�g���ո�3) �5�M����;�y�F��w٩��;�"-��w[U����5J�y��6�܁�Jz������OC=����r�1�͔�1�,����.��oe�Ȓً�o�DQ�:�,a��y�t/�32 vC���Tq��v=�D�� M4�
v�ꍂ,6�r���;��<c 6��rw8�I?F���+*�n@~��Jx�Z)ɔT��<�
�`�����X�R	+���~O��j>���{��]�=瞾�{�&C���F�[�`u"F�
C�>����������oH��Zl�m���²,�ep�IF�C���j�E�״�;UG�����,�R�l�^��J��^���,����j	*�NX��@Z>a&��t��֊�(h�����\e@wq�˶s�F4p�q}Ԯ����� r��w;̺�!�j� �}4��3�����<��v����W�6�GZ_ �����fy?�Q��/��3ك��FՇ�L
AX#��r� �F ����l�E�%��`-!�����(È��V��r��΃^��8�Ʊ���
R2R>]��e�kv��HP��ۇ�|,��rCŸ�����y���,�g#��u6��)��H�u�T
����Io�%��S�_���
�x]y��������-5op\��$B[�5Z�̫,\ICx�^��b�4Zף	��a��G-����a1�Ɍ~M��v�Q�螚�6�'��^R����M��x��:��pr���0z�_�m��Fs	��R�P�8�����uag`�R��
RGO�8&!�H�P`Ȓ��QT_6X�K-�K�# @�%_89M�?j��:8C -��z�(`��έg_���6D�=B�4�� ��Ӽ�e�2o\(;���l��)\K����0@ %Lh�Ue�n3��żh�:�� ��^Qk�H0�djuX-W(
H�e��a��됝�w�gz:ѤR�xR�H���1��&�	p�S��|i�$��i4�N$ǿ��<=�/z��BcE�
�X� �zτ�BYCJmLem���U�h�yoU~��L��vj#T7v7FT+��S0���F����t֛5i��SɌ��*{;�N ����E�g3�����3bg�dqn��4*��gM�A������s����Ǳ��eb�|4���)���
��0��w�Խ:dv�GB�N��3P:���s�� ��U�$�����<�G��衿�a<��2{2y���ŋ�ôg������uv���s��jK�\]�6���T�l8������)~a.��<���[�_}(�1�B?��g���\D*����E+n��-��9�0�i���f?__S*�4\Ѯ��k����y���ɧ�7��N>�~-��C�dN���&���ǽ���z�E `Ͳ�K���e����wL��ϋRbVFGb}O�����Y���|�mP��l��"�¡l�Q�Z>����W��6G+���*����; C�~�?ț7���^�u�,�W�u�;h���M��8aQE�<���8Nk�:�޲l>������}�HГ��wwwCz/�����k�}����Z���r��JR[�	 +*�.����,`���XX�&���xM �>�`q��'��X֜�[R��
]=� ؚ�j����l���p@�B��!��?��О�~G��.�	3>�~�A,-#x��m,[5�@����$���2 <h+�����o���H¤d�
�'g�w�:fuG�#ج�Ɖf�&S�X�����m7G�� �dATc�� �|���
��j��&���Ȩ:`�9���G���o�<ۉ6$�����J�@�_��<ڣǁ۱�*~B�>B����he���Kz�X�Mtgńs4���$V��4D҉bj����ɭ�C�gч0�nx�c�3���3��bL�r'o�a�Ũ���X�,��dr����c��
&�I�B�.SK
���R2_~��oI������va�aH)�@q �@��^n�g�@�J>iN��/�tH?;���~p-�����s��M���-�Z�!_�����C�gD�{�{��^�E)|Y���8��;�k�ҭ�h=;D�f����N�%@�cDG`Ў���Q��|�I�$h��l��$t{����^��)a1�Q�<BJ5&r3��(�Z�Lp�h�*�ZU��"�ABF��������]�t~N�մV����d�����_��S�=�����3O&�gP�L����������_�����������z�ΊR�����K-�[���`�ЗC*��#F�[��
��"�JK�l9Bx�����hI)��X����+�]=k�zG�J�OuFp:�t(�ߧΜ�&ݼh�|�5{З"�A� �T�)k{�Lp�:��v�4��6��!�&C�NHK�d�{�G�w�$�\s�(��"-4;��ܛ:�'{�픒�4k�3s�jf��N�@��t�c����ë����7ry�\�|���q��q �������.,�j�j1<�s=��s�H�9���S��9�Kw{�wD����t��d{/C�F�_��)����2��� O���N~�����ݏr���PJ���U��5���C�9�L~�!��-V��9@b<�c����v�ӱ�&�j���oh�F���Q��L?:Mj�f��ꉠCgj�̒N���V����:�e�1���IJ1L��Iޣ�8��:d^������OpN�I�/�2��Yk��
�:���̠n���6���Ӝa���:u]���VM���Z�=���o��7��¡�[]^���Uޏ�}��%�o嘴gr#���������JOg̾�Zfs�������ācd�����)�����F:LE�kA`��{ �e�v=c
6:GVe*ф�p~���j?#��2�4U�O�im�,�
����G�Wx�vt#� EG��͎
� ��CCe��v:�Z����Z�0@Ά��v*��d0|O�X��gg�TD[ H��|���kʹow;*Hb.�*���y���J���\^���6����",Q�O�d��aR�,���~���O�G�v��ۓ�8
����T�QQ�՗��WC�,UP�Ujʓ�����-���Kll���S�*�,Ś�bm�t��&ڳ��F���щ�[;�6d��S��\���ܨ�S��xh�m��EC1�|e�W~}Q��QS��%]�,�]X#Z{�Ji������T�.��*c��4|���7w���<�X��ȉX#<]Ч��Z1�T�U�Y����+H	�"������zyD=ݤ�)�c�>n��R8^�m��#���o�|wk��Z���)�
a�E�x՚2�V֠ѢI� J��kN��>�R|q���@n�e��0d�y����j�9�Y��o�q�ip{+U�L�G*�El��RXӠ���| dQ�i��٠1d`մ��y��3�f��c�dW{~���_X����q���┋݋I��y1>���gK�#������ٱ��3���_y<�ѝ�'��A�P���T]�qF)�q=�_�վ��r� � �2����;X�~�P9��#W5�2(
�1����~�0^��\�,�6H��Ǧ�f|��3K��D�o�Z*0��s�6Xj� ��^'G��L��6��}v@[(�5������b?t�<\<���aOZ�:��Ւ@�9�}7UjTP�36H`#�%�d��d�	lJ�MZ����RV��0�γs����@P�\�ɳ_ɋ�$B���4�ی�y�,����z@� �������wuݧ���{J ����oQj�����p�Zk]o22B�?���A=�{��1Њ���9����6�w���������a��\_̧�(!.�f�}4�͂�Ҫ�(�h���I��$߁���v�_R4��{~f7,�X��L�Lv]��ubNs�1Q�����<�k��׀�8PAk.X[n`�:�A*
N�T�G!%bj��P��������΀+���LV���N���.��ؔ�*�d*�B�u�uR�L�	� ZMM�����WJ��{�j�����?�(޽��|~	}z�C4BUw��㎵DTVE�BP3fa�_�V��W��]\p�S��БN���`5�(��~<�T��_��Izo�GR溮��A�HZ6�͖�~���y�{1��㘛�A޿� ޿c���l�l���ݚ�R 2Y�)���#u�/0`0�Ь�����pc2�J�����P����>���������(���� ��L �ڬz�sj5��R��>s��}�]��n)Ȅ���W_-_�'�eA!�o֠����|ͷy\���R�j�;yX?�x/^�$���r~���|� Z�C��b;^�F��W��"�2S�p���s�?נ�x�e�'��N�OX��b�j�5����V�_\.���������#��Y�T�G1=�dbn�Dx4;��D�,���V�`�q�`'ۛP�)�e�2mëtAC������"xm�J%�`��Z�fjOǮ�?!��E5�u���[�{$$��ot�ް�RQ5S{A{�X]��k%3��zo(<U�iЦ�+؍'��~���?\y�*ԧO���M�ޛ�~EwU�ӆ�j�;�R�5�n�y,����>��x�Ŗ��B�(�:��������:[G����~
@T�e� JpE�|��m�1R��u�A�� Z��9�=j�v�����{y���j�A֑���k����^#���`�l6P���U4;����RM�����`]�ۋ�D�m�L���F���)G����A���Sh��2~�y�k��ƗB*t����q���(�)@�Me�j��o;���ʔJ0A�����x5�P���ǥݑe��C�b����{D���Uࡪ{J�q��%��{PEl��ѹ;���:!kEQ���<T e��h�B�_F������kؔ2hAt�2�L���k곍�<.(&��Ze�����##��ث�o[SKYx�����{z]����	lB��Y6j��>�N��ʑ߇�.�l~Lm��v�.8s�������*]��`�u����<,m`�F�*�cSfKm�`��7g	eG���*)��/��s>j�Y��s3�f�O�eǝ�r ���2����R]^di���&m�L�� ��3&z��*���y��;y��G���l�2�����ӎS�_��Q�"�L�c��$��;qf^z�t�-oc-�Q��Ț��Ԩ	1�v�=�5�\���=`�;��E  ��IDAT
���Kט�>kİ�Q	�^{Q�~/v�F��D��'f��h�����/.W���,;�p���l�g�ryq)�٢�T�Y�od3@e��ڂ$7��� @俛8�Gq���g  
F���{�����Gy���||�>��5A֡k��ٓ�섣�ؠ(��*��#	:�7
O��p�:��_��_|�fY�S $�����d����)��Eʛk�Lg~MJ�-�O�� �
��s�k|ǻ��3��*��+@ ��6�Ǎ���;���y��$�0�~A�J�n������D���|��~�=����`���hʜk�%<������o�����!��TV�:�.�Ȃϖsy�A�*� e��<�y_�w `�|�!XC�����zG�5���s���P~ߋ���X��N>���g�����9���p� ��n2��/����R�5^]�4ϱ~Ҕ��DU ��#['��PVY mYW��x.ؑ%{��_��Nn�D�7�߅��=�����+X2GjIS*�B�Y^�w�ly$$ ��M3��ȲKl�ْxk�TZ�κ�žY�	��9�ީP����l|�y����A�|V�]�p&�u7="�zf
{^i�d���T��J��6�C
<}�^;��8�E�As��EX��*	��Q3[Sϡ/k�Q�JE��C�����S�d�g�D�ר�9�|w.Ǝu�&2�`cg�X��:�)5���6��TiF��b*a�l�v"��6L��&jkEUh��8�DjD,����G� $W'|/TP@7�S��b
�0�ٲ�GoQt�&�~7<?%o<�<��������yq���Ŗ�Y�&���x_�p�̘�#�~̖�y��A� [PJ���<;yyk ���^`5�f�߇�Wiy���B�O�������6֔���{+���*kS�� j��9R��� ��'<Q����������x��_��-6q|0T:
k�#��6�fa=Ƞ}w|���������A�%�RT��1g�j�F���mu����(3�*?̌NRǐ k>��p{�4��f]|Cϕ�8A�Ԥњ��?�E����L��M=�/E�@4���F��5Q��,�(�f�T�W��5j�{Ly�#*b[�Jm9�*�m��U������M�i�����();����Uv�`���`L�?�����P\���=��21ؕ��x�����4�
����uAO���ҏT�).�� !�y��-������8�D1�ҁ�v4�V������fr�B���G���u��<<�ʇ�-��G���S�
BF���Q=lfq���u�pD��n���q�׳2dP�k�C��{܁&5��ݸQG��A50�c��=�a'Ѻ,d�:�5��
aZ�Ʀ��˲1nYS���Ę���
#Ѳ��LTZ��˚UE�/���f���{�Z�ƚ���'��Щ,<����y[3�Ϛ1��6R�@v0u�(���d�	�=J!>�Bd�A�~��}���R(=�?pO��?I�]��{�vhJp�*lJ�l�N��	c�=��o��F���g�״��2�C f��G��u�7���T[Ix�YOn}� p�	����m����F�Iܮ�h�q~a�NZ������_��o�C���
E4Vs�ZX?6i-۱�2���ŷ��7��r�Tq�͖���[6�UEb�8�\�` ���N���oz#���#�y:����^\��{�4k���YM5s� Y��/�q�Cp	}7�{� 1n��L�����?��$�#��b�0s��� `�V	gh���y��ej��R{B��߲���K&ƖdQ/��Q���:�=N�3v���b���L2a���R�4�2��̱&b)�1?j0�l��K�k6J[@�yB��6 ��q��B&V��lnk�*ۼ�[����%�=+۟���<8-�� xt9�S�.b�pGt
�X�hh���&g`�qF�0�ЋC�AG�4�ѹڃ�"Ì2ܳ�L#�8��RX�A�5�5�ѡ*�8fv��V�z�
��s�LRu<�&�>f�|L��`���(�|^�q�Ae"���z���P95��j��	�7�lO������U���dA��C^<���������F*C�e�t���yѤ�S��>.=�-�H��s����>�0��Fě;��wT9Wԉ�l��3��t����Z>\?���F�<�'K� �F�b��Q�lPe�Ɣ�4���.rw�?�m������k�BX��	��^#q�
��������Ą�Fa���h���l��X���?=Jr�o�=��^l�-�S|'R��?��y�UA����wD�Og�����WU���Sq'Щ{�<B+PNw��ԫ������������Jtj`�u-Í����`�����"�#eSp�����-@����TX�N��.\_�;�йE�Ԗ4V�_�'J���mM+(�@ 7v�9Y^L��JVX�qj�fuI���}�&�l2���A8�Eʾ���Y	�ˇ�>;>�K��&��&���|d疐�������ј/ϳSy�G#І��RQZ�n��E;��y�2������bw=��s=�>��s�;R���u�Y=�5m�F��9�%Z�qϰ~��{�~ g
bD�!Z`��@tt�v���Mv�2����$�w���x+7��Sx���fP _�@v�Q	1�UմUU@��
i�������(��G^W��K^'S^���ݩ�+6��L���d ��
S���{�C #?�{a`��ꨥL²��Jڼu�cP���c��v��*;�-� 
D-��3��`����k��x;QɌ¾g�� \p�l�N�< 5<�v��Ƞ����}µ�{~�pnf���n3�ܫ�3*g�k�&�G��";v�iBg�������E�
�*��a����Lu\�(�[�O__\��/���_�d0��,�yP���ꅏ���k�G颩�N�`����``ؾ�2���>v�ұE�*/���a�����@c�A�Al��>X�K�&��r��o;2x���w��g?�o&�)��6�;D(:�m�MI�?��	�Ǐ����w�~��q7P]��B��+X��aM,m��S���z��A8���ʡ�a���)�D{��c~�}�{4u7�3Ւ3�C�1_�jz�[�,�8����)2[xDS �p>�38>�U��X{r|�g-Ͳ�h+�mr1������b�R���Wh���2 �=���b��U?�4Д��;h�~�YH\I�5�t?�`Fu;� Ö9^أ����p������мc�_�Yo=dkYp8�3�һɱ�I: ��BGX��J:�Y(�pc�m�pө��8N�(�p�"z01��n����h��hL>U��R�jB�
%
nF� �����Y�|��$^8v�G^��KD�d�5�^�-��
��m�wu�:Ȝ�T],��>Tf_�h�U���@}Z具�6o���V#Ǎ��&/.�L����q�+����3�����NiMC3����.���)�X��4N͐u�>O�l賡��{�8��۳{�rL�g��y�_���Y"vySɛg0#��nv��nuȈ��lಝ�ͮ��5V�y�9cp��ǜ+��(�؈.1����P�e�b���i&��Y���-s��3Tp���4�?a4�N����I��	���O���[��U�-���\������/y|�=��AZ��c�}`��e�`P�@��X̚��<�U��O�23T�"|��,��~���ܢfރ�;z��
�<�� ��`?�:� �H�KC�3��P�)R�5�Mc��vq��H-Ƴ�M4P��S��N!dPjp:�ru�t0b1��dC�_
����
�İ�x�,c�k H�;��� �C4e�)#�g2�-H?Rc�Ö�q��Y?�n��c��?����?
X~�����Qэ�_|8 Vf�� `�w�{�@z��^���Y�� G�гM����m��zK0u�o��������[�!�0cV�e߳����@�]R{�9�R���H'4�3�=����c�M1���{��5ګS�~~E궂��}�m��6j�Rè��e�U�@Vh�N��.�4fS4����/�eu���tG���?�������1Ě�(�t��G �J������x����|�ͯ)@�����`�{�Me� nw��Y�#��%�e�l-XӦ��z�=8%%#�1������~I�;��6�΁m��*b4�TH4�XS)�/j�,�H�D�h9m�l>�m�d�`��R>]�����Q�=O�>vJ�H��?�k��{�1�s�|l�e��
x�d��&��(t0x0���Aګ��u�F�_�|��7�y�M9&���Zׁv0o)|���	��T"���6�5ێ��_�!�&���(h�"�/F{d���fų2��E��6V}��H���; �^L��g�yo���$�űz(���=>����جVK���`OQ̏��N޿{+��ޡO���)�IT�=F�D���(�Q�V�4d�`%g�IՀxRg˵\H��,���WE\�j:����ys�Nj�6��z��(ˬ�@��-@���[ ��_�^o=���p,�Ye�z��� ȃ	�V�7ު�5�&ME'��K��A�4���PT��Ib ���yl�r<��R�:��ۖ��lg�JB挴���{�4�`�&k>�강�����
�Z������bO᯼�>�ƴ�'�m�e0��ǻ��|8��&��.9&�"�a����wy��1˛e���C�p�������e��NJ��.�)B]��V�̈́Y��3B��
�]���Č�9����:�4Y��٭,Vf�28�E{0P����!�g@����KoQ,��6���φ(oZh3�H���e>ތ��ݼT��z
J�Mš� �+b ��J*7otOތp���5�2[c� �Bq2��*fJ�/}:���;O���0�ˏ�}m����_Ƌm}� �O�
<���d��"��M�&�7�um��Y�v�|��(9X�5�J���zf(F�5C���2�(�F�bDA!���Fi
���>R�Z,*R=�!-��h8`aƵú3���ht�zI������fź	��=��Pk��4��s6j0��FEeHcW8�H�݉��=�$�P�}�0�b�� S��b#Ga7����Gm��uXr2�Og��p4G��'/�?�#���G��ˌ����~z͢�� d��� �~p�@�YX��p�X[�lhv�7�J�����u��CaG�"���술�-rP�멍X�V�p%���)|vڸY��*u�(P��d�Ɔ���+S!�)�������ubM0�C̉����̪v���c��iِ9��|����7��o�9�X������O�5A� T/%�2^*X�u�u��o��3�]���7�_�^~��o�b�b"볹'xe$פ*��q;���г$�_����`��@�'�b��j�	GFc��'��Γ*����:���R���"�%3��nCQ�dʸ���f�p=���k�4�i�~�gL"3�	�O$�؏��} j�kC�Q�!�L�R
Y��@�L�*�7�`uLPIE��/� ��2��!�L ��p�%���GϟG�a���6fݐ�Ǭ���9v�� y+3�0��A�G�1�J*"p԰�X�V�X?ݠ�'�<L����
ޢG)�}���SlD�O�����ybo�Ή����5��.�&C��ŋ����K�	d��e���w��?� ��7yl�V�3�J�x�{�`Tq�$סq�5�QdY��"$VAV��c�B�1;�}���Z�ڒɟ�)U�&�C�U���<�<�T�ͣ�+�=0��OmK�R���ӓ��^�/����ۓ�o1��.Ν���%	�X�U�|!�����ۣ��ѦBp�O)B�_&�ֺx���I���O֤D��A�c��B�=��g�c2���V&�ɪ��p2\c�:�r"�MPT`v�#x;�l�����
�]o�3j@'y(3��RqZ�T�4��PNn�\t�����%k��*���������TK����?�%��J�:r�*�"� ����95@8��8N>�i�Ifg�a[�ٳHf�4���)�� ���c���� �]��u'�C ���JܙCH(j6m�P�	^FLe����q����tm��|���T��h��k>OǇ(N�	��\�QU5(�lr��Փs|_��:(��^�7�^1���(���W8�p�N�+c���5�R�x0�j�W��w���Qc�@�\/��U�}�c�n��lȕG�q���Rg�V�z�t��2 ZS4��+���9=n|)���i�N!� a^ӡ�D�A�Vc�`�i�@ �kuc.,��M�Y���:Y��v������6�Ҟm$N�ST^��:�W�De�,�v�W;���6OXd�� ��T�BZ�>+є��{�x�yȫH�?��A|��g�U_z��0
�����f��SAF{EP�Ez�����[��}/������D
�^�;�@����bmn�Z'	��Yv�����z�MR��E�(����fdjƵ)T����s��	��6�Q玎x����jpE���@���I��TĂ��Ԏ��� !3̒�
�Y�a��>���s��?�V����_��������B޾{G�����٬����bj�u��F3qbYr��B�J���R����e�����'�E���;f
e�罏�}�T����9hk2�����]��	�P)�A5{�M,8.Z7��}uu��!��@P+

//.duu)]��е�l.&�2pCG;���6k�L�*�5��w�P����Μm� 8�3����5і���h�uCI��h��S�l�נ����p� AV���7��!���|�LQUU����?�Ȓ�I�Rᇨ��,A ]��w)�ŒA~
� 4{����o��A�� ���^�i�>A�me,$�^��	���'S�����΂�(��2�(�N�,��	Z3�G��^�D�.�ׂڳ����������Oyo����O��G���?�f��4T��?ʠ�H)�Q�T�
�o�iK ��ٯT��	�Y}foR���F��VK�Cq��ĕ�8�\�L�O�T��9�>��H&������c�e�9���=�z���*�a�9em4��h&v�~>��zv�C+Yv�N�����߼h7O�Y�A��F�=���{:ܠ��6Ml�2녉�W#T4ǢD��g�Z�ɮ�<*��2�\�؄""y���[j�����D��\��i���7_մ5�\}	�76OPI�>���1j�a�;��R��Oo�)��z^�@-�l�S�Q���ΩMBCՃe�I�mZzg�9�nt,,D�3���0͆	uZ�-�i�T�kM�%*�a<u�� ���v|�q8^���B��ų3�}��}���' ZG��u)�6��c��E��l���,;�gr�,��S+�|N�l����)�:2�dw���w����� ���m�}o=8؏b�GfZ�v�`CH ׇ�V0�e t=�<�e8S?���R�{=1�lk1'5?2h<��ɾ�Ë����~E����j�s�{�ؘ�jE�z�jEe��s�����SOob��H2Jn���
�ݬ�nK��H���'𜡵���f�g&v�b����6����@��Fe���)E 6T���Yo�M�.i��Z����g�A���}6����J.������c�f����L}��&��=u�G� ��͗t-���jf5����2�7j� : i`��4oZ�#4&Dl���(�z�TG�����Ùǀ
nhz����GF�Y7�(.�,۟ q�EB�cǆ�I�ŇQ��}p�#s��Ȏ
8�=k!v|�f�5���?������ Y�:O���g��D����#�L�}�w�>K���6(���1�Ί��ا�Z �(`Q�����dP(�3;A�u8b�����v��:��f�p
���)���lI�n��
�Q8��r����#�ċڰw�b�ބ6�Ԭ�jC�᠙�#)�=���?��L�^�cNLM�����4qf���M|�4g���A�g���zٶ��<O��6�._(�P��F�9[�����@盯���˙,�9�r}q)��K����x)_B����&8�43���������ܾ}-���M;P����|���?����7��#��R�t*Kȼ��AFu�������A��20^�]jk	쩇���@��fΑ��6������;���{�B�9�u�q8t�e�u� 2?xm��Ы�X�.�wj��<�k�|�BV�y� [�������G���;yw�Nv�{�'��L�2����RX`��U;�ڽ|/���,C��.��� :(n�Zo!�є�R<���9�Z��!�c����f��/��m���m�7�M�1�65{�_�ǡ�l�^��v��Y H��4x�/�G�_���fPx��������_�6QA�����!�ƪ����?�z.IŚ\�Ag��v�K PQ�̬%eu��޿����]����wZ�����&<�od�y@R��W4�>N������`��jR@���'�y6�l$4$i�����]b0���P��2�������s��^�20��(����Y.Y��j}�10�vU�zw�c���m��̆6y?l������H:	��Ocڪ�r5l�F���1ϙ�i�j�՜�H3"d9�����)th#ݨ� ��D6���K���#���fRS��nK:P<�e# ���Z��(�jd�n���}%��R���O�s[PV!��F��|�|L=[2:��;r,�,�A'v�MZ����$Y�iM ��e���=�c��k<:<j4 X��&G;�ߌ�x�kt&F�	�̋q�#��mhgr��ec�I����{�9��a���6��o)������'f���Z�͑���wC���4����/�5X's�"����e1��R�{�Z;5��x1h
�����s�Ԥ���>{������a��P����`��۵��5�[i��T~/G�S���b��8-�e���0���ef�'��@�u:��0|b�2�!�&�C�xo��#�@g6s�٦��� �#�r�����J�z��sZ�Ė-硣m"I�o�c�-ApQ�Ų�y���V4��s-�f�`Sc�	���|�K�؈:; ����hO#�@��L%e�?)Bb�`T�4�f�Q��T�)PM4���EY�^��1�*2a����3{��-���ʤ>R�B�������NP�����'�;�_�C�0�O��Ga�:;T��cv�d<���`ak1Z�Á@�~����K�4��)��0ڭ=�hD��NX�ٞk��`�[�`�Pܠ�m%�f�2�+��Q�
�j:��q�zM�^��y.��x.{ީ�V���bBi�T�lb�@��~�
 �^\�����C� �ѿL�?hߧ`Y��	����?��������+y���w�������e+�q\.�(p  � �-T�p~Wo?e�s��eI��lā�Dl�5�b��+?|�GJ��T;����y��fqI��h��TFm��V*��k�/�������\��/Y�������ޮ���AֻMiGe�h�_7���z��7X��w�=
�f:v*G��0H�j	�T�w�}�o촷�yֆ���c҇)�M[�mJ�2��٫EiS�̶����	���'T������Q��x��-'LR����`�Zo�L���Oը��Xsg����X�T������߷�5�������'�1�~�N>~|O��M�~���r��`�*S ]ˀ�2T�f��k:o�Pɪ@?�V�dt�N���V^9��cR��Г��"����a���)}o{�2����FOdN{�U	����2Z��A�C���B��Kx�Km�i$Q�$p�$dx��Y4�Ds�A�-̦I Ȋ���8|&y� Id������je�ܞD����PTG�=fXɘfĉ�4�14�T���=�7�	�5R&�x1�Y:�l�r��1+m�@����]�C��cNw(����o���@j��R	��{ +�=���J5���0�&��̀;���^!Xh#�Qd�\���d��,��?�q����0jw��Ɇ�B��M`q1��������h��M�� �]��v��Od���F�њ�4��`t��걐U�d�C'VemxS�H@����ua���2�|�tq�Y$q�Y�ˮ<͐�~�T�a�FɁu=G��I���~�E����:)���LM�r񧠮�m�F��u����5����Ӡ��3m6���n����v���7Oy�NY��D��^���ыX�L�ޭ٨�Q��������҃�:e��:�4XƬ�� �<�,4 g��^Ay�Б}���{v����t���j�b���$��I�3OC��� g����J�l	�ղ�h��� J�M�-����t�/�P��ϳӝ�劁/���~��)��O����ޏBc�jQ�eD�1wؗm�=�H3cS�	o�4�v�M�&��߷'�X�����3�:��҃��j�p��H���t�aZ��4��-to��@7|��SgE?k�$~����@b>�i��W2��U�e���9�꯰��eʱ�M@�꘼a0��-�q��a[��W�p�~�:��M\o�1"{h���?���k�Tb_k�1���Bf��2�߼��Х<{v%W�V�my|�s6Q�S����wrww����CB�(����r~���!��î�ml�i:G(�8E����������IC��q>�w������	GU�����7�� 0�jJ�M;��"A>i� L�x�|��^�u��9�:2p��Ľ�6<��̌��;��f`(�_T���CK!��\�.�%����w�b�������L"��R?��߱G�W���{\��u��i�\�l Lܣ�b٘���`"!�;�J��9hd�G�f(%���ɏ�/ۇ�d������&��{*F�u�����nά�D�?�OܤT�)BK�3�%�0��}���ȷ���%l�-I�+9������t>y �1y��h>���u�Tx'��ˉ��κ���=W�S������
f��'�N>Vo�s4����>��폪'�PQ3��$�ba��x35J�7ڇ���Q,r�g�_�)�`����D��	����ТғJ��?i���KC3�����U%�Δ�9���;����-��8X��������:��<m�>%-RӐ�DM�F��ۊ�ra��|�{����<�0Z;
f4Rn����!9a��#x����Ngk�,�34C俣�CdŪ覾�d�r����e�ǘ������_���ҿ���(34�t;F��w:WB������vF�� ��Y�%�q"e���=*mF7ܓ$>g��C}���$%{r2��sn]%�� :%��_��������?��x�!W}����J���X�~R�5��)b�]"����;y�\7ߣъhyF�6��L�о���0������Ѡ�#@�ev����:t�XSer�ɲ����S���_D�jT}j_�����f���b���촠>O�W+��LI�
�<r�Go�[=dY�����ͧ�,b~@sKP��v;m�<��ܠKz��d�dl |��!�9@�8���L�+Ćt���甿�l�X�Y�Z�Z"����J`'(4�I�J�ҮE�if��,�`b���J�A�*:�8���̀�Q#�՗�U/��(*}��;1*]�މ��eK^ ����� �,5�>%I_�\��(l�ٞ���(@V�8B*�5b�$S��4���׹~\S��p�� ��z���"Jn�X�
X_k
a��Xw{wKY�ۛ$�����<��c]��
P՟Q�8�IL���2<�U�_���>�߲g�:d�
�=u6�l`�γ��v~!/����7�$�|�?=�d���"����:�&8���6�?��{A)1%� ���4�����<�.��9���yà���l�==�@��t����:#��d$0��A�no>��B���Hjv���(s �Ժn�Z>���M�M�Sֽ��!�;Ơl��Y�N�p9��9�/:X�O�K�3� ������J�2����t�̀*u�D�T�1�!�E%�c��K	ȡo�}�������{Y��]��п��h���ޛvI�G�j�G�G�U}�	r@�p��~���'��rH�htwݕgD�����aY�@c�/��def������������6z
��=2E�4m�]���L]P<���Kk���O"E���.���R���R����C��X�rB��-�g�Dū��i`2���@ cCY2kz�����7�n�E��&y8��(�AȾ�ޏ��wV��1I+�)��.�Z���TD�S��k��沪��)��CN�)7�p�re=^Ir�.`MsVf^[��w|�$e8|�����:XgNy3p�ǳ\��}��@IU��Xe����O��0T0�q�a�R�.< �[�\�\�V?ҁ�ACT=ϣ�%Ҵ;�f�{��J�n#\�s��>�XFWՏ�6Q<=��Z�՝ț��UO�'�%UEkTv���o��EF�dcE��cȗn�X26A������4`�LÕ7�Ø�ҦyBuR���"Q@D�|(nv��܁��14`S�?���wv��k�l䷳��`8�hn-A #@^n��C���;f�A���'�I���tP:u�A�A&��|Uek[�PI�Yƛ���ͱb*����f�|V��&�O�-֕�,t��S�_��3����^��Z���̶S�;sp�N�us�h��j�:�G�(D�`1���#:N(�^hmU�FT�Wpv�MT%�{��*�܇�޼�I^��}�c����\}�"�^_@�b�ө�YdW'nc�F�5�NJ�V3m��i+�
��^v-�U]/�<�7ƿh��z���qiR$��L`���衆� [Ț��)����}
��ޖ ��/��5�H�'��W��>&x5����5WGk�p�I�QK��r}�ԎZ��Jm�o(�j'&�қ`�G�E� �TD}�ΐ�o���)Kͨ�|��_R�ِv��7IՏ!�o�%�$��S�|��v�0�� ���\���aA+m^������f{+�o>>Τ�b}u�DhfY�w���\���L���}��^>~|�>h�6QW0��q���އڧӋg��������%>����/�!��[�X���l14��.�CPkJ�V��l��-�!�t�컂iک޲XYw^�0�2�,�d"�b�$�1�����f~����x�_QȺ����ț7?��A��F�Mk� ��F��|�,���ߢhba�
����㙀������&� ��8u����k��j�Q�!�y�DI���Z���t�-eHa�G�@燏�����C�#�,�K�OϬ���B=�r-h�s_��{f�H��d�Y�*�O����+A��A���H�6@�Ƿ���|�� �}��Œx� �ӟ�9g�x�L{b���	�Z�����l!^՜X{�(>l1��-k�@˞_��
�*>h�^6߲���H���u�2���坧�H�c8��G��U�}5�,)���:��^�"MZ�Փ��kt!>+�����h{��D���
n{;����棑*l�#J�{�`��MW�����;���6a�hXRˆ,b̵(e���/ћ������Q~�F"�]��.���A�d4�x�(�G�!f��F�1��?��b�� ��؂Yd�U�;(�����F�7W�n���HVO@��F�T��O�5�j�A֬K����¨�70k��Wk<D;� b������?�y�Os���j ����s4(8h W���UhW��,~`?K͜��a�1�{6�W���E��ۇ#�����hk�-��i�;u{n�1e����b2ۡ�Ś�}�T7��uF/��҄��y�3�y\��#�+�1����x.��R��(h�%��hP��ܭ{f}�ON�����sy��qqV/��OP��J���#��&:��w�����l���I�c�(jq?~x/��A���&��_������V@�{Fo����ZU��l��1S��/�M��J����"�tD�k�)��5���<���֬A'f��z����Xg��W�χ�ɶ����li�@i2�����r}W �����(����3y��Uqx_���#ʁ#��Z��a���< ,�q! ����Y������h��l<Ojs���GyI^�����M�?�6Ս6
�7�c�,��φlN��t��j$����g�^	3�P�C� ǕH�3�u�CmA��=��8`'D��<�ڀB#zLMPA�� �_=��d]��+�b_�/cs}s%��[J��v��(K��]���?K�����ڟ�z%���������݇�$��Oo�Z���<nT}����>�b$�����^k���W���m&�����������T(���\�r�s��>~�F���3�A��8+��2���J�.���-��ךi-��-t�Q�����MX)-u�����x@�hu�9�������L�
i�9�y�}�	)Xt���u���鋰�^ǈZu�L(�	����Ş[�ܓ�F?O�I�,�fR��J�#/sb/��ŭ����J'�0�3M,t��P���s�>�����u����ߒ5½i&H���X�}�J�s_�?k�߅��E�=���u]u�U	�r�-��)�+�'�YZ�'*p���,�p7�Et^v�� 0@^��3g-�j_������l5���<e�dX�+q�L�Dz{�L�K9�M�e6�E�g$�V��C�#=�8C;僻aS�1[O�}��� ����^%�}��6��<�W�^�G���`�.��<C�%U�/,F�-_{͑M0��H����s��� �p<kc��W�;S�3����٨a��rҚ,��6��f�O��2g�QnU�U��̈x6��P4j�Z�-���n���rWvW8 �I�|(�` U���6�d��5X�Kg偋8��L��y���8���f��-aOr������(��/�� '݂Rnм�����>e��+�u՝js_���&~����4y�����Jr�� ��g{�.�a׌�z@�FAi�]m�`����2�m��9W��N7p��]�-�Ҥ�F�;����)h����W�Y�J�P�I� W��С�f���e���5�5t+�r\\\ȳ'O��z�葜�����?D��P�x_��>q�V�MF�ϡs�۔A��t^,�Sȩ��xZ>��?�'���PA0`�NF@�AM�҇U�w���ُH)�S��¡���ZQ��M��s|oMxV�s����7:԰��8j�PK)�y�)�l����T����XJ��F�Ăs{V^�rR�qzvQ�my_���YN̉�hF��ޫ�d[AE<9D�NH~d p�	Y��W5ڎ�@셓ѹ�Z�:�dO���ni����?��5w��
{t!ޣ�'a����Y�Q��Y���u�W�D��le�H,,J�b �}4�6F�M�A���$3Ca��{��~�_<\�$?�r��7�j���Э�e���u��Ky� �OXW�꺎!�`���b�q֚V�����z����!ǥ3io+�Щ׻�5�v�BATGƞ�=�8�[�-��G����$Q�2�*�q�L_b�U�>�}Ec���1:�#a�؇�~L&����
E��!_�gl���!Z�κo�m�<P�������c��������IU�o�=�]G��x�l��l���3[�k
-$�	��u�}l<#�*��hD�-�։$k���G�)�Ï��6�v`�4��uk{=�ϝh_"Qt����%7�]Ek8��7��L�5��H"������Y�3�)~���枊Ӆ+��_&�9�RJL�Y��=�V����l���;�����N�Ŋ�Vw�d��\�`G�{�A錞���d�ul(7Z�7�u�%}҂q<c歷�8�`�]����0�J����������Sة
S�m�D���<����$ޯX�����{b�(us6n�b@�:wS�����&��@:�?	��GC��*8jF�4�d��O1�eQy�V�N���_(�Z.f�)@��p�r���I#��
2H:Ga/�#]��6�se)���ԞR��ԛbe�
l�*�e�s@YT���/����H��D.����0*#���""�}��ɨq�G�@K9���U�Q��?��t�4�
�r ���'p�>���Ժ�v�٣߷!��zTc�sE��Z|�7��<�٫���p @忽=S�>�C�Q*a�|4�b�Mgs�w�u�(ѰZ�s�^ݮ3It�z�]Si�ӂuSj�����o���ò�"
�Tqm�P�����L�=���Źy���)������Ab�;4�����.�8�� n�Y{ o]�⢗�aIa���@]>z,�����������e�|��1��e)3��b"�Nzs@)�����n�[@�׾�����S�b�QsF�mE���j��z���k���]��E��3�D�AoC��@UeS8��hVw%T=z�T�=&�^�(��iq����?��bO�p�1_ U��(�7���A;������'y��D>�-WW���,����sT����(�TV�5w�C,���2�����KY�)���`������IY�K����YMJ��Yd�[�	E&��& �������.��$�^����^jGq�u;�V"�l�֎�#�պ ����������D�[�e������s�<y,/_>�Ǘ�T9d{���(R����f��]�U71ѡ������Y;�l�g�Ƭv&Y]h�ɂc��K�z��Z�,��ur��Ā;�'�`�]2Ål�ݞ���%��{����!�m?RA�������f��۱+[.���gv�O	�����*%�p��=?^ �����b�;�ƨ���jE��gi~����o&�&�G���={f��ԧ���3L����g�,�l�H[��kN�@�~�k{�ϩ�	��˫�V���%[si�{?��>��~�J�[�ӂ�����w��:g��>m�(v�`���&�$�B)��w��yB��'К-�7��`'^��a?��iO��[�Ղ�o��z<�BN2h7+��m{���p�{���L�}^kv���� ��ww
�|y�=�=����e���U�y�~6oP��_��>�gh�*��hiIO�ɑb�~F\�;>���IW�jޛM�S,2E.���*����~�;��>C��F��j��E*f�N8'^�Q�51�� �~>S�VP&�0F&�\�be���fk�G�ͥ3����D��Mf���ؔ؜P���R�E��hJ����/.���G��S����k�u��%.��]����K�����Y�|����OQ������
��9f|���[1��ac���lX��Ҧ�^�T����ڳb_�S��y�VKE'����. }JQ�>��7{"��5x ����V7�R���tD��&�����갈ӓ5{5]���RU����L�?{*�^=��/���Ǘr~z�N@]��=�f������)3�y��4[��4�L��)I֦�lڨ�(N�is��X�pŇ�&��^�'���`u�l�FN�g��Jm��h�1�<�e|�l�E���m�W�����G8T�*$�t�#�]���Tֿ���J������ﳗ����/�8藏�	��Y�| �
_q��RNjŢƫa-���"���R��d�@���iw'���nS�e���v!�~u���:kh� ��Z�eMc�o�O������ ���� ɯ�z%��`ise��D����\m}�ހS�2c�q3����q�5��k׋��<( �@6�]9�T�n�V*PtЂz؃� Mَ̠�.����ޙj�4���4Z~��9�MՎu�,��A�=C�@���v�O�A=Wv�J�#�[�,8��:�~W��={�=�3�h��蕞J��������M�?}�����m[��wĞ������ɓ�p-
x�F{]w�s���c=�]��N��g�Qe�7�5R���?�C职�0�{���j DI�^Z�Y6�4�5��dL�(RA�5�uc;�m�V\��kj�q�VK0� 5��d{y�����?�w�"{���3Oݙ/$ܿ�b�s�S
V��r�o�������S{� �~��|��J�f����	�����!b�Nլ�;����q�@0z�-��Ɂn�$�H�_0e��W��T�ap�	�<w\Z��\Xj�0����"Y\�xVz��{ƝLrY���Q[[0ˆ�06b�hA݈Ҝ�J>`����,^oŗX��/7�ҡP��3W�&�Gb<��4)��T����:0V��}~a��Z��N	c����VExtJL�ۡ��G�����]1�ҙ�����ZlP����#�Y�;e��vƆ�ŉ�)�<$���ٶ�� �N�����}��-�ivD�Y3fT�lY.�/����6'�=�z'��ٳ����9�uq$k ���{6K,*���OA:���h}L���������^��������QAIޟ>Ԥ�G���DV��ȁ�C0�~Rr'BT%(9Ht���(? r��v��[:�;(q/41� EK�������<�(��1n�\����X'(Q���Ś=ǥ��M�&���\so2�n�;��s������(<?96j`X_�|��+y���\��R`�i�:�F/�F3�~I��z�}d�qn�b�d�ٴm�����T�旼7DY��8ro�f�Y8X��N�$.�ް�L��of�HTڠ֫�{أ��#�Vqj�������^��"%܄/�N�꿣�B�m�W��)��Y֧��ꫯ�٫����%��;�����:X�ԁt	
R8W{K��� R��qG ��9�m�����*�a�O��V�YG�ב�J���z[-vX1��[�s�f�i%� Ԭ=.@t�3��A3PT�ޝzw�t�AmLb��`����7n @�^P����e��p=T��mTcW����V�­��3Y���G�^��n�dv�,�%AuC�`�An7�E;9�WG1W&�A��N�E!x����c���Z5Ss�-��}a ��`
��⧱�j�򘕶��URw� ��\��D�c,nٲ���Y���0��I./Ni[���X�ݤ�X޻�N�p��q���BF~�ީ\;���)֍ʣ��H$d�!��ʩQj����l��k���G�|�}��y�F��=�,Wʦ�O���	���l���^W��z�Zf�����gQA�G@O�W[���l������)��̆^z|hvR�k��Ҟ,{�T�E�?����1�P�wi~����q^� �g�yf�R!�}��W���/��\�C�sޮh�~c6FT�������oBG��ձDD8�9n�F�u����ά]$ Y6���v�����~
�R����. �f"��H&	t
7�bu#�޲���3H�.:NfN���5X� � 0��i+��b ��8���y&�
��d�M���d�r�Y;k��}���6��>y��{eOvH�-9B;i��-�����CW'D(��N|����w֫!�{}Q��G�X3Iϝ ��_����"d�s������ׁY!`F�lP���o���;�����)+GMU��� "1��������A�M�v�4�|����=���%m��;G ��p&��̈́�-��X r
��g����)>�yl�������� �f�Z^[�%�RA��̧�Ԕ�ZG)���r[��:�\0��P%b�}}1`�#��]ҵ�ɳlM�f�pũ�hUg�������'-E��P�P���7�p�AMr;�� �r�̋��xDT�J,G�.z2���S�/�7)�<��KCAcvvzV��#��ꇲa�f{���C(j.�<Ԓ5Q�hr(�ݰ�r~y,���+����;���G��<��&��1w�>QHk�'<`Lt���y�z,�~�QL�8Y-��ꡘ-��c@���r�uq�.�s=!`��~_6�[�ͣ���sQHGe��2��D]���-2�-�O�;,��␽w�֙�ᬀ��S�[���-����~=���Pf��b��һ><�j%��o?ݖ�E�J�[����ӗ�ʷ����ꫯ�|�k�+t?���z�ɽZ�������\k��JީpK�^Z�Z1g�=�����|��Gy��{y�����9w���]�A�v�[�!��a����W��D6���S@8N�A@�n7ڽp�onM4E�뾀"dz= ���M�a
�GuZ����;�Afmպ��398|I!) j����M������@bW���7o$_�6���JUU��< M�7��V���-�@��_9��U'����TΕ7h�{L��U�g�-6a�� �[�d���o�(��)-�|�!������\{�����7���ig˽����C��;98�,���>�43@	-Y�����Ʀ��b݁�D'K��Čx��\l,��m�q7r0L���p&������rv�.��Qtt�D1��i���6���>&���ݎ*��Q��
`	�$Cٲ��4�E����]�Cwp ���B:B�j��G���(�Q BE����Q:�!�L��0/p���we�ܒ��](��ttRa���g�Br����Y���eVYrf|�L[�izFF�M�a�O��q��v\s�͞��YDV���LN�EvJ�Yk�T�JL���k�g����@0�ݻ���O?J�6���o�(S��W�J�,�����T���3��3T�O�9hS�>2�?�Ț(u��<!�� e�|qgbl�ECw��`���去�<u�%������]������dΪ�B#���9�bS�Q'�i�mTۣ�����B��T�PQS!���҃����2�W��o��� `�� �8�l2���&�<��H1��2�ܩO�p��/�;���بƿc�SU��|���zD��Y#������J�X��<+u��'P�\�4�0���0I��Yу��Y��p�:�0K���1/;�r=�r���-,]������F�L�"�ȩ�[�y�D�>?Zw0�
vP�E���'��J>!j��y��2��ˇS�����{�,o�1��ւ!����,���ZFM�(���w܎T����=�����M�WĨ(3��(���i�Qi�Z���Ȕ�9[A��^[Tf��]�_&2W��82�	�/\����SU5m7j��3݂0Q�*�C��o��F���7���s�����M�v�}<�:�Dם4�?G}��� �Rd�?�����K�z����7�`4�e�J�QdTtf����b!�*F���zcu�(�����wZu�}�������W8,r����uB�`�]�f�w�@*�&W�׃�y�����^~-��HdH�2ʘ'��H�INR�4�
�)�A91�������	�2j��'��B�AB}C�2�w�ؓ0���ق{��:�(��m����9-��-A��ω�MWl@����PUa�O�kEPggM��42��l�ɚ��yGt_}����Ϗ��H3,�CM�Q��T���3wwJM.ˊ  �g���=K&����K*�q�&�P�����4�����u��_����� ������ƶ;N���Ě�Bx������-{Qݳ��=3Wo0��4Z��4H �ʞu�ҫS�&�h����xd=V�PqgbB�
���@yFCȹȩ2���3c� x0�6�0P�V�+�b�|�<���(@E�Λ�Z��s��kb�kd��	h?DfA�X N��=!ڻ4�{X#W=�Z�*�V{�m�����Z���܇�zo�U����;�F����hꡏ�����E��e���f�4���''��֢-��`o$��@ߤX�c��]\��G�7��}�~z���l�l�J��k���X荟��o��~���k���}g����$�2Q����C3��p5��Y��]{���$-�f��UX��ʉDg~�I3��i'��2�j`ܙ!7|R�6d[x(0_(�oޛ��>��d���J=�)!���@&�d����p�5�ҼvM�Pr��w�lQ�Ȧ`�d��dU��\)��y�i k�����&��Er
f���UM�2�\�et���~U<�m���T'1ل'`�5svu�Y�-|ŧ:1���:�h�X�C�/�1M�*<�Pm��}�`��R���sS�<��~_0�2g{n����_1�b@��� h���k$$7��0���Ek�$����ȸkZ���:n��"~�Ul��c?���o��Xr9�K�6JW�J��n6���7 VC����ޔm�c�\�J���z�D�\m�<�t��ϔ�����g���G��d�+}N)��~��<}�T���[�MX/_�`����EFC�=9ծ�-q~�à��+��A��^�����R�F����K��@�x�����L�={�\�Y�Rg�3�f�^�@�Y@���l����뻡�|V����8�>�f�u)0�z�71�`W���5�@#��� ��^}]��K
�I��j��dbEa� �>���]���|�L��3@(}��~y���%�:>}@�e\�p��6���p�e�^�`�R�f]e��8d3��7^l���}�,F؋��9��ƍT��0��o��\��ȣ�c9:X�:�I}�m�<p�{��߉~M���}Y�
�&�qj;i� �=E��� AR@e�nP�1
�n�6��?���_��:.�:��A18���<�x�>S��x���8�6+{X>����.�'��2�]�VEș�Pd��sk��
<h����`D��!1��s���R�&���9�?�vl�^�9��3jo)����{��k�Vt�k��z괅lL<Rᨀ���g�a{�c�YJ�)͕/�Q��J�	�{�bR�qk��y�'��)9vZV�gat:�Y�����Sy���B`��Wii��X�Zq��o��"�:!E�1P!=\Z=��X��r�dMdu`��_*�B���!���O�G\�������OSZt0����w��v�l���B"Y����$�R'xM�丢J'�g��!U1���_�K���G�aB��s5,I�V��@�Y��0JcE�"�nc��x�8��dè#�������3V��.&�;��5��L��-2Y��'�ff�T��ˤ������/&������<Mw�����|��=��j;c�����Ľy��`��N��^�-{n��{ϲ�t��s�@Gy��b_�HmR(�H�9�3�ڴx�s��lO�Μ�Y�G��g�*�k&��S��݆t���r�S�I���x�(|	�f��e�c��Q��������t���8"��O)��]\�G�T��t@�k�޾pd�~?�?c�!���n/���eٮ��FX-d(���L���>^Ζ���m3!M�-a�D��Yk������VW��NuXR�}-����͛���͛b�oxNR�;�Nl����������u,���w,�Gt�5��5�A&�u�^W���<�����Cp�Z��}�-�.���`��ܕM�Iq~��G�}���I���o�na�(1W���4=X ˕:vhl<�}d�kjv|6F������z�q��vj����*��K����i6(�h�������7��W_'�?-�bey˰�')��<�&�T�^¸��c������>�4I��z/vxxB�J"���\O�ui���`Td�7��+կ��:'�����n��6dh��Ḧt�2�}� Ԛ1BpԦL�X�.��7_ɳg���l��x;-翥��"���_�D�w����T�r�=ؙ_cYj�ٕ��ׅ0*�!�t��{��PҲ��n)�1˻�e���MX׷SrG�����< ������#@�g�#�n���Ь̤�0<Gd� ��B��9i���蘩T�lR�8S�b��7�jw��?YR�@��zqY�-��=����k�@��2�*(�d���&U�_��(�����U�s�=����8nQ�Fj��Tj|����|����7�����e��@@}��"����e�P�d��@A��eR��� �{`o�����0P�R�,�1֢�E�an<A�N��5xFL�j�^���;Ȃ�DrPS�L����DK���Z/ ���qr~J�����8���)�#��h���|����MDI�����>@����!R�b���+lkY��7���4d v�A��α�%mF��A�"��E�I��os�}�ȹ"H�RD�HI �l�I�(��z1��,ݭ|�F�<m[��vP��n���8ږpξ�����p[0^ǥc�f��O�/M��9���ʤq��\�����p�;��ͤ�o�~K,�U^����9�Y���lT��� G�.C��A�ܤ���n�s���)�T��Yh���~���Z4�{J���"*3��½����¶@�ǹv�l�����gG��%�{����*w�s���K�w��f|b<��4�l٬zM>��`|ᚣ�D��>��R���!�O��TgB��e�S��g�3׾;<~�fj�4�!�Ա���(P�B�k E"����My�R|�]�jX>���ȕ�s(G��T^�f�������������Mq@�	wF�Ȥ�LlR�:U���wT������\}M�uqqIP�~7&��[U;�RgX�n-W�w�ƸY���`?B�1)`�̋ٿ~}$��˳�������2m٬�tA�`�x>�ޱ��iA�Vd��I�mF��y}~��C�jU�̩���Y�ZB�{)T���g�X}-�~�;y����S�*��_2� F?���&h�r��َ���ط|K�ȉ(81D��
Cq�?Nl"v�be���{r��wS���ǩ�Q���bq[���Y�s}}#WWWZy>�Zx�B]�&�nت���\\���HP"�Q+�wtt*�xl��W	�&2���ݤbO7U�c	��3P�g���l#��tpt&G��rV�W<���������v#�߽���;�����>.���˿��r��ب>S�׷;�v uX�8�O�D#S*�Q�PӃ��"��-cY(�H&���@
���T�LXK��Fv�p��ݵ��u������LĞ��fp� ɎJZ�4G{�%���nŹ�֨���Mz����Q��L��@�1�r�ӵ6G����_��o�w��G9, ������������Oe�F>Xp�&{0�)���(x2j��̀ͧT��>D�\�O���+
�v����˹��ތ��J!l'�R��s�>��Ku3�I�� ����(�� �ZG���[���T�������������93Y Y����&Z�@0�ӧO���[�����r�~���vE4U�/�A�zp�IR��tu��y���z"�S�cP�|`d���7��}R�$���F���#�h	)'��o��u�kf
�x�t�LE\�Æ4�7 f�.9���Zj]�5���pq��ױh�CU���7�*�*���!Ґ���;�9��t�NM��Nj���d�����ԺQ��Ҥ���sj�+mX�_\%�qp�]�;`�i(@qp�1u�YJ�3F����Z+ب2�>�F��s,�}Q���Z��?�����(,��'h�����`�R� �.�� ���i�mn��gk���\i5��ϩ�����)�}\�T���]�����l��B��a{��[߃�1����,_�R�̾p���Ј5YL��/3�S_z]�ݱ���(�l�'=?�S�杣6��&���dJ�ؼ(��i��Y+�T���U��餇ЈxtSm�g1h���9U�� �'��7��ŋ���P�%�L�E�锌��B��|u�j{v�	}���g��j�NrA�h-
�:�x*��Ei�Ooe����z�Q��P�X9�&A��%��en�5��>�h�S4�g��|a�����s�*�k*8`�ҠK|E�!�W��>�/_ɳ�/�h�_*4�؄ZZ���[�~7���s}�Yۏ�?�
��'����9zj�b��`{�� �Yv^��;Ĵ�S -�&���2��2*�D��^��J�3&n�Ç���;���f�؅��G[:�~B�lZ�ܬ�Y��2�R{�u���Um�둭�B ���@*�Ԗ�_���Y���z����s8���~�t�l��ɥ���;���o(k~us#��G���;��G�~����$I���܎tb�h���8������l�!�zp�H^�y���s9)��7v��	b�hpJ�X�8mw�B��y��ѿ���3�q�y�@Y+sta�1��C]��[e�����:�V��[�~}p$���W���J��[Y_�9{�(Zk�YO��i<U��Q�k�� ����;�o��7������w��;�
���T����y�>��z�]�Z NUW�4�?�3m-j�vcb6��R���S�w�h�=�0ؖ�N����4��l�|���M�/'M����i�8�(�➲\�֋}O��,;�-�}u3�(A	<<:�^���R�\��ݚs��䈪��Z�ޱ��`r6���i��{M���}��~?���OIF�(���Bk�[�&�f���r��4R���I�����u;Ō�eVg�?H�P�>-��L��<J�à0{�}j&K}�CW3Y���A8�q���@,�����hIH4Wg���EQVj�C<L��|��I� R��x����� �N�^���f/����ݟ8�iGι����?7�[̃9�׹y��A�g�d����d���7�v����Z�߈͹R���0��Y��^��o��L����ך��g��]����¯�����H6���k�K�T1<�Y��>s?�m	���߻�K��ϧQ��l,D+6�`�q�^�_����f�|je��M���o�R�Z�����"uA�q����UN[����~/���v25+���\"-�����������~Dϩ�dF֕�2v��;�y�P����Ϟ�����^�
T�B���e������?���*�#fX8��������Ã��k*N���T�<{Y�ʷ�}���i����v�gF����ةd�F�%>Վ��\���I�Iu��z�mu���JZK-6����e��t|,��g���#9����6Ŧd[���{�8{g��.�������mBj�u���T��܋��G�hu˾8cgr~q�:&�,� �6!�~[�5[�A����� ��Ȁ�S�_oj˛��J�#�;{��㘩�ZiP���ٴ4a��oG�c�>T��ї�x{Ap��4ؽ��bI�I��:'�s�g�����BU��D����O�eq���5!@��'��鋯����=�/ �œ���d��U~|����?���G�n�r}}Ga�rY!,�B�]��Q��G����cy���tPOD&H�6�N�i�c�kΓY�GO�ՙ������G!ȚI%�I�ʀT9|I�g��_a_�_�-��d�����4PWX>{��T=UL����)��Wy�@��zDu:�UL�@8.�����o��W�� Z��(��?>B��%�%櫊�Z.a ����ބ>�PҞ,�µb�*�&�LE�E䬊� H�v�J�>L����^1I�5jY�_�zCn�����&⢭P �У/Ԩa�x{�շĞ���qy�M�] ��5����1�c��j����m���4�}u�����zf�3����x�y�ڞ�2W&��u��鸣U �q��ve��r��.K���T,�Ҁ�=�n�>O�ۙ}���rB߄>�\}�܈�D�������`D�1���<*�l?�WǢ�����sL¶�y��"���ut�������V��C#��=%�qrpA�r ��p��ƣ3ŭ%\���ߝT�I�V��Ȝx�@�X��ڥ�z��s��,�+��z�*��f������C�f<c�k�+��>��?�xꢠ?g�����goƻ]�����N�ٙxֻnn��&n�O�`�5P�����	T8�>��ᒆJY{��x �{Q=��/׀�_T��O����?O�,��YB�܊t�nG�*�TZ��)@���񆾍��nL�T��� �
�Qs�6h	�[�A�{d���j9��-���D��_�����wl=c��b2��Q�5bFۛnW�UW���h��k��7�����o6���X����eƱ<~�\>~|+ן����J�W���r`�����.��d�H�e��k8���y���W<��K6�K��ۯ��|t|"���]����A쉔r�B�b������9��E�w���)4�Y��>��:M�R���]:�9�2�z}$��eʑͺEC�͍t��O�Qzz�d/�L��������l���±����74 �B8��r"D���q9j��5����K
�R��DGLfG��:;���)��{�i��{����$�~��4��N,��qd�@M>=>-�)�����rT�긼.?�6��.��y�����n�����ObP45O�~g�d��b�:m�o����O����ݽ̻����ē8KƩxT[�}�/�7�6��!���� *���p;���P��j������ߎJ�Ml��v���"O�(���)*c��uHg �Ѕ����T�h�2`|d�z�`��\M�$�B�jړ8�s���9{��RI]��<KT�k���E��Yb�=��%t�waݧ-��=e�ҤA
�'@�Zګ&D�xF��)�UV�,������x�:'h��f��w�^u�t�=���R�V���N�w���k�{�w�L��76��A���@����j�:)�����b���4>�s��>�7�����7��Te0I�t�U�bJ46�F&F�0�9M�R�%2`�Y�������gs�5T���ubϮ08+�5����lZ/"8Q^��7�<�����'����u���[��)Ա�ӧ�\z������\RS����U��Ţ�Ցwu:7*���Ȣ�H��X釾���!2�-9�S��1P�٬�u�۩����Ʈɽ���\_DX�J��w��9������������m��д�.{�Y��*����_'�� ��~ Z:-����
���Y�NnlS����~���Y�)l�C�k�:���9�_�����Zb.(��T���v�7to�������1i�o�U�m!b���0�t�ȑך��qO��wf�'���Yur| O�\ʫ�^ʷ�|] ׅ6T7g4��pP��c=��v6׋�X����t��^���� z]�]<��O����|��Z��=k@�X�&n!.,�����xR�J#�}r ���&h�%}f�~=�Gu�M�&i���e^�v�����C9<Z��_��ey-V���S��Gx�q�ʙ�Ϧ��q{?o��N�l�}ߣ̡���Nb��D�YF�y�(��5�J��L�z�s���f;��=��WVŐX炚�)�s��vG��Z�l�{Wkgݣ��t/hM���]@�v��#�zv.�F_�K-����%l1"Ѵ4����N�xN�C,��H2�3�g�T �G:�l��i�u�=R�l��
"g/ĀٟT�UR�\�F�q?|����������rc�A:�N3�f���1�_�\�������ǰK��o�=�o�8ժ3kbY�R�o�Yc�f���mWd�_v%�I�)mM�2��Y�A��BvÁ�W�>t���0�4�0O@Ce�
�se�l��և���*⍣��1{¹X�&�f�'����5�+0M0�̏��~ ��p/�zi,�L�W#LW3���\ɰ�:�5�b+b�2�z��Wj��ٕ���m٢��R���m/���+��@Kt���H���,wcm%×٪�@��K�{��>s��}�#P�����&��HD�c1�RY��']� �Q"·Tt�Yo�����V��\�]cDdM
���(�i��p�Mj��Ȟ�>���γ��h�xT]e#I�K|��أJ��s�m�땫d�ß�U�}�Jߓoj��'Vj t��iuPg�O�MeN>�r�2���� 5(�-'B5�nr��?�G��Y="� [�T�M��U C7nG�y��lҌo� �<�D�U{q�u��3<8�(pcS�U�*�'5cs�z�ώ\o6��;����_p`��a_�>��zOq��k�K���R��r(�
��r�4<�*�x�Ѕ�=뛲���A����C��޸E�&jv ���JS�x���l�+�v�!�]���d��"[�id���� �G���sy��4��f�e-���k[,�),f[�}ۃ�s���̴:�$�����l�f��\�v�H_�)@��&���3�>c��i�9w>������\��L*����n��C���51�Nj��ډ�1���[:��t��<�Y�9�c��Q'"���猂��� ������NJh�}��Z��rMjhCh� �>�Gts��@� 2Y{v&q���쎘�\��Fڹ�5�5��q}oz��ĳ�!�ӥ�_|����P�����~e/,�V"Q�"d���Wc�S� b�q���[y��-e��PS:#%ߋ���AD�,Ț�h8=���
c(�=|2
������e���;�|�P�P�ޙ��ĠՆ��!����*����9�P��g�TI:�rr�VRb�A%;:<`@�3�.��`���Nvm�Z&���,�����k`Y9F�η��Df6�U*"��q
,�����@~-�?�,���xt!x����_���s�~��	�&��v��6A�I�hDrg5��~��(��'��~��-ܟ��v���YN5��[��7�c����?�;�o$j�.l=�F�MՇ�+Eu�d�=�@G��f�܊$�i�j�j875w���4+�{3�i�AUq��b��B��fk	�@U�����d�O�C�^�!y�(_&S��@TE�r!;p�Y�T�B�j��*-�c��l��)�C4!\�$�8j3¼[�B��	Qj�вr����}��=tX!2��bD4�@��ⳋ�4w�I٬���f�x$�5�Ɯ2'd[��rm��6&FE�
����YPұ�|�t�Ns<ub��X��]�GM!6��3t/���9�� �_KJ�h��nTC���I���1�z�^�����pe�Ze}S�J9?�$�g��H>��b2���ih�K��:�
0tC���9�H�j� �Yu����k-���Ӭ�̟�l�x�J��s�Ei3>v�]�^-�I�����_DL!���Pr����LS(��\h����RD���M�?��]52}�Tzfn�ۇT�����J{��+�@��vb;�4(�i�t]��T�>�4��3���yK���5 ���g��]Y���6o�lj$��3i }��4��R���v4�#�XL�Hw�@(�0����O��꣡�9�5��pA^������o嫯�+`��s�xۇ"lD���_��O��q�����d����c��l1G�~��Y&�FҲ�>�X.Ξ˻��r���7֠�,�����F;\����	T�m�����Z�X7��J2�j��|�Ty�?@��x�������b�j=m��垏Amu�X�1@�l)%�滨	�7e>�i.�"P�*{oVaq�H�Li�j�.w��j�>B�e�hg��b9�t�sb_��)ڢ��ڌG������侇��=�.�C���R�2�V��rn��G��a�=���2��%v���+n�W�7��E����D��d�Tij�t�Z�Z�Q�\��Ή:��*&6�}��my�/�.6�����iq�7z��:��lj�`8ve�G�|w��M�@��3V�5�&�a�>B�=�?6���]q,>����z��;�S�#�<o�~��=%iX��#���؇���5�(�޿���f��vh6�-X�Sx��8�
ا� v��h���.�ݙ-*svBM�z%��SY�ɲ��ږ��������õ���^������C����h6��ӫʓ��1�W�)�gt��y��^ {Y�����E���<�<���.��bͬ�fl]\�������o���\��� ��HI� �ĺcm����㓓2�sf�.�'f�'�8�\�	�X|lPD<�Q����?[�c�{U���J�gMt�����rgtJ� O*����,�zRv��A.T���e�?��S5�!@0������I�3��F�\P��1on &�=��uf�&���!��gSFƕg���Po�\�l�T?!�_Yy_�OKd��t����/�� ˘�7d�TYfs�,������e{� FX�#��%��L�Au��M4|�G�_�&����G�����b�m��x�p"�H0�4�w���I�d��v�9����1mF智��h!�D���.|2{5�a�� �fʏ����Yd?�"�g���v(�q��*L{��/d%rؤ����k�w�͝9����N�y��j����d`+�]~������� ��\I�Q�1�v�����p��G�;v�_�Y�p��tC�q4� @�4������q�qm�)̋��M��x�2�{͚�?�g��N�"���U3��9?��zbf3�q�i��?��8(�IB>:|��8��w�{m�ȷGD�o1o�^:��Y{��nG��:��M���4�"j$�fӫ2�M$ڨՊ���z��� ��9��5�q�r�+�3!l��8;����rN�zT3�i��4�:�u<��W����|�g�m'�=���T[Dtq�If+4B�g��=��[�8��W����̬�J���:�Ul�>?JFC���h�~ͱ�c?�>���e?����S��_�<����9����-(��Y֖-T���� �xM��6��wR�Q����"�Y�S�,�~�}�`��]�~z�� l�M~ݟb#�ł���(���a�֎�<��}|�^�����X��fcʺY�a j�v���8�����;��@�����}�Cg�4#Kvw{#'�'r��q[�|�����%����l�R�#���Ϡc=y �S��6��ˮ�<������MˡҊ舩�nC��kD��m5Qc�6.���>e��r~8��^m5`���뫛2We,�ɺ�nI�+��X�����2��0 ���#�C�_�
)�����x>�g��ށ<y|!O�=�G�.������<8>:f�D��ӓ�����vs�z�G�1��9/ټyk{�H����f����|�^�x̓��b�����_�����?+�_k�zZ�+��\kn��~Z]��F��=9[�y���U�I�\�� �Խ�AӾ��-���B+m��J���7��~�q��=f�:���������9����9��#����y��� �����n�)l��!��YO�b�4z��X��z`�a�P��\/h�1a6}C�2��k�*��z�����(jo��:)��9y��̘M��٭J�#���v�*0���Jw��ͨ k�Q�@��g���|��M�f����P�t
^MzXD.�D6K<�������qH�*����?��Zp���j�T
�E�:�T��[�#���b�w��ߵ��E!�?}L]_����T3xfT�	k�c�<��(��F7m�ɯt���_�[-�L���p>�\m���TR}F��q��h�\���:�v��w�����s=|\���L����Rj�+5�F�Ѡ�=�eS˲ِ��YSC7�i��&��5Nco���
��6峃^�^�a��r�鬗_��T<��(�

r�
�B��ڛ�w���>i]jfg����3HE�yoVy#i�@�7l� Z֧�TR+�FM*���}�>��^���Q�^��>��<�U�[���I�Q3��e���]ظD7�iχ�%��Z��	���j<�Y�Zź��8`�,��ӕ
̜-�	�7.�(�@�o6Ƅ��]]P���PU�?�ٮ�3�����ac *�ۻ�>\����@��� \wduf*H�uy7Q<J}�����i�� @2V�߫����O�U�RE�P�=.=��/_�����EP��}� �L!B�kR�� AӬ�����Ʉ�R9'z#]\^p�h$˾[�
��e�"�gF����_Raʫ�����ᳵ�U@�gwwI>�����#�j��i�{ (v��Z��ψ��/�f!^ٛ�\ǽD�������/�DL��т�	
������`h��c�򻻝lFd�(�RΔ6�g�!|�Lq!(�<����|���)�~���9n����|\�䚳ϯ�k���筡ݗ��l�G�%J��#S��:Ν����+հ����v9��g�l�� 
⡍Av��0��R�C"\ck���j�ic�y�5�:j�:˺�i7f���&hЪoT>��P'e����_@��j{O�C��a�q����CT1*�����1���H�h$3^�T�i���j��JG����U ʴ��s�s�nD�� ZF'TL��H�/˜3��̲XU��g����G���~<�v2G$�4�Y��~3�����r���iD��*������c�x;�䑅�� �>��A�T�ܹ�E�D8�9��a�yd�QH���<~�`OO���Q��
EuJ��x���>�$Aߕdq�������@���z�g��z$�W��)�WZ�{���c�C �pc�z&��!8����&��@�q�])�S���o�r��Z([Si��6q�X�����=��S�]\a�����E�?(����~1��ej�������j��ug�MYµ�2�x{�����M�ܗ�s���8�FBqޓ�S9;9g�+�U3��]�6�e����ڣ�3(�=�\7/���s�Px�����|T�m�<����sr���]g1���_A���ث��}�]�vp�Eƅ��_{�:�U~���w{O��9���V�/��{���~֫zϮ�j!Tqaҭ��}�"��k/��{�"�0سP&�_^R��0P�U3�����y�}����B������?~/�����+R7P�5(��H��`�j2K��+��jϦt˲���������ȧ�t�p;+�ׯ�uvϯo(t
 {��ʂ��2�"b�&p�s�2V&p���X_48���;*���6@><>����7�?��3�*i�>�g*�d��|Rk.@���F}Y����-�N槀�}W�ɧk�d]]]����@) �8Z		�5�eZ�#��sVd\e*�n�{�l"���y6�ԉ�>�F��p'b9p?�?Y�]�+�XQ�c�lX6�S��b�=��|�@^�����|b�/t$H{���NE���6�Ȅ�����k��ut�ۚr�I�/���L�L�D��P�m��T��.m>�v_�g��`���L��[��_��b�`b��@�Z�xO��ʝ����.
�"$cv*�}�=3i�V��f�C�{��� �����7�l�1E��0O^�YeVzA��j$��܄�?v��E�c�\Dc2lԛ�;	���V����I	Ny��<���9� ��}�>D����.�`FYrYـ�Q�9��E���FH��
��ި����dlm�ʓe�P��o)7��(~���ؑ)�e��Z�ǋ��o�J�W�	 �Z��!2X�'�LFz�+��:?�ʩO5E� ��㾛SsF��d��AC�(���믋u�TqMih!2�$([Ɂ�S�<�����,�)��D8@�ť�Q�v�z���Е�86��1x���mwJUL)�>�É����0��?s0�x�9��{�
|D$ސ���`���`_�^ǯ�Pџ��(LY
�x���N���O~`�l��l�r����_���6�jШ4��?�$�d�>h��.F��zf�:%���Z�Z��ᱬ�>���vM�e_�?G�l��/E[���? �S=����Y�Úa'��"�.��3[_�(�	�q9w�+�k����mǭT�_�����2Y�>R?TD�\z��fUf��Z�q�:���?���>VŅ���z'}q��]D�ToL�{9��?W����7���/��k�:�<xUo)����0�T==;!U��M��o	j�)� �� �����~).�A��n�?p��������7��m!A=��2�o�Q��x�%0C�n;+k�6[�$�nd]�R"����M�5�{�������wpzB����R-���gJkTf��i͚o�ò�]q4W+f��Y	�D.�:DC���2~��g/����Q0?f{F��s��d�˳\B�@$�G��;�_I0��9�@��w4#�71�E�*��Q�U�q�g�OX+A��ڣ'��^k� ��}F���O[�zl��M�J5ɤ*���㼚r�ޙ��TQ<�9"`�5��*����)"2�G_p�ɚϝ��p�8m;�]�ŵ>���8GǙp=#�����,�8d��ss�gԱ����A�N)���v*�[��V؛T{oj�Μ�.���*����߳�P��Iݰ��XE��j�����d+�@���G��p403�`]���GI��,��9�.��ua�K's|r|� @Z�@\#�{t�ĊE;:�J޹�dW�����0!E�[Q'˝n�JRITU �Y!w!�eG�v�,�i��<����ɴ(s�"�J�hz2�D��12T�b��;70�����}H�'�m�=~�ؼ�(N�R|^J^��W�呆���p̶����ţ~uR,l�6���d����y�'Q|��_�l}�w&��s�#&P?W*�3�!�g��]3g���~R8�m͖��թ���i��0Ek��)�0�s0��:��hC�, �ay�Ge��V��<�
��G^��1�i��9�Z�@&��]��g*|������_Z4H�ϼI�W���u���ȍ�p�gVl�6ť�*�ϭ�a]�n��C���sA¦(���*w�n���-l�h�I7b��$~�)御�������+گ���d\����|�Ŋԥ��C�l���:$u�7����}?���/r^�QE0*�r��5XK
Z4
��$L�����X��f���X6�\�f�_�6~=D�ap�>K���������~�"�lԝU-5=�����+Z�%"�ޔ��sTq�ۊ�w-��Ņ��*2���k�/�=�8�� evQ_ͭ]�l>�ڵ^Ջ�T���_�p!�g�O
���d͞��[-�_��l�����?����O?�H��,��s��o�H��ܹ�Z�)�־HUz�+��2D�*���������� �~z-��t�"{L��(�M�jP��lo�lIdp���Z0H_ ��l�P�N8=��b7O�N�����2����N<7]L�`u�AEy:J�@�-���ڟ���E^���������7J�BM10��;�^�S]��p��`{��9+���|�fS@�튾 k��L��z7()�c<O�D�Iǵ���Ӭ	@
h����䘊�-�*PS��i&+?c��`�9��L)����7"�l����z�uQ)րS6��|ϷCs�|�}�R�{jcX/m�8�2�\JӝB�>[&�Ǿ�,�e��V�:OV?Ϭq� �[��`�ݔ}u�we}l	�t�o�X	
�����U5Mec�@X�=P�j�M�+[��M ��e���
�<�3��ql���H�����+bc ��E?�7��Q�Z<jÐӜp��R�㑓o�ۚC�7�]�{�wk�����}�Jm�D�
 �燾B-O|s�����ެ�+�g`��]��%d�N���.��2�4��Z�L:CɏHB8Ǎ�܄L�Er�(��ek�[�3�7�,����57� i;Fc�p�Y���I�]��b4[lNc��i�xeaC{��- ��r��٫���>���F��d�^w�Y,����bqT��h�2\�^�(�?���$��y���?��������֗��c/�)���g�y��	I�������_�\�<#ѭ�p3W�h�Ƀڐ�=�����^Ё;ݤ�v�6¸�x�v�Ԭ�=+���F�:$�L;4�L/��<����Z��cS���5c�Wk4J��c/���;I�z��<�U1��?����_[?�aLͻ~�Q�=��s�.��R���kY< �5��t���$G��mU�Ƴ�]\o�H͵<������R�j�m��N�5'�=�j�݁MDW�hW��cv��V��l���~���_\�<��f��X��Z�*���Q�Z�^�iu��h��	F�i�h<WR�%y���wl��lV��l5��sfS~�x�s 0���ׯ��� a�N2,��������,ɘձ,s_l�2;U~�YmR?��b��"�;��Sf\���,Ӏ���ͻw�ͨ]��O�*"�5�ّ�>]ק��M���ZZ�jzb���8����"�R��wk�PiD����D�v0,��g,VZ���/��B���Μ���/�-�|=�����nHY��#*C��n�4�����dB4��ܗg�!;	s�q�~I�!���D
઀:��������7W��?(� �+����v�VBԉ��^LQL���	�^gm�4�51�Z*��������W@���Xe
��g��,�E�B����?�c�p��ZCL{�f��cW���'�vv;�ۮ��Z�\��g�k:�Y[��D ��r"�X�m�Ѹ�?Wb�z�^j���Նy-�ǎ��ΆE�t���د��������!v�ǥ��쵶n�ym���Z��:/�g&��hA���(S�:du!`�M̖v3� ��y;3�����6	����k9��o�w -{y�&�$��Q%�%��l��L��{d�D� �4C���{�ı�`�P�w~?ձwG��H�Vog��ŜϠ6�g����2[��:|��~���y�3�Yluw����at��p���g���F؊hdO���k ����H8�>m�?��~ƻ��v˩���q
�'�:�i4��Ѱ\ύ� �Y�%��y:�� �V��7F�L����Vx#ƽ}���z�%@�3'�����Iu0j�����b�{�e�oZ�<sr@]zvPn�G3�n�s\W�,!����	�9mY/�}]��OJ�5��e���@�Z�/��I�ߌ�$�6ś'R�h��6�	�(��8��N�Zg�c#�kܩG��)��v��	 <|���h�#���9�g㞇�
'����"���C��&l�8��-��Ю��{���||��R�yf�ú��W&k��0D���1ƿ;��KuV<H�$��9�۹�ɟ;~�
��Bb9�m����F�;��v��8mI�X��8��ȷ��\A�FX�́��iW�&Ev��R�gc����G^{n�sx{{g=���Z�<>k�P�� �x/w�3o��uO*��f�ww�,��Л�ɮm�rpo5�ڌ��Jݚ͈���A�z����nF��� ��rQ�,*Ou�I}#=����^�9==���c�mW徆�|_ ��n�v�3�0����O����;�Q����d]�u�cS�1+�c#a���:��-���?|�T�����h�#+�{����k<+��'��Y��2�<w5�HȺg�p��i���'O��wh�qp$���d��TY<, ���Gc�M�g�D"`��A�P���e==����/ 3��	k�F�KxR�����*|]Ɉ��_�}�Y��GreX�m7�B�du�RcK̯�^�a�[��}������Sx-�[�G��/f�<&�c�g�+O!T��褨����|xm�.k���t&��g���f�=v)}a�} ��hpfd�U�����P`=ˌ/[7��Rt��"1�T�Y}���:��=�\iF_�¼�L4� 1c�����i1؄����& �S�j-�D2���h佯-7;���l���F�*G�"v]PD�bӁ�+�d����*�X�ĲX�/�֭Ԛc-٩��:�����A���5W���Y�b���׀0��6�}��M��h���H}�7 +��g�R�Y�u{NR<�m����"�s�ID$5#��f,���cU{��}���dͣ]�F���ňK��R� $[@�&�����ψ�����%׈M\k8)�H������PK��hr�h��%�+��e��Op�hM4�s��Z���㽰��p�N|������{vɒ$ׁ�)K�z�Ո�$8\�=���������E���{���#�^O�  �;_eeeF�4�k�Z�7�dՊa�qk��^�if��a�&c���P�z�Dk�u)"�!����BA��[����F�Te�q�W��^��� HN9T$����u=�`�y��s�w�x/�Wq�|%�066`Z���n�����j�F�]9�������������Zd9��)V���0mX��#���a{�^~��$��D;���i=�ek�/~fM�a�i	�hh|	�i��6y�Ɂ暹F�YӍ�o�ę�@����z(����P0�4Ѡ�:#����|��R�ې�����G������@>���	?�<N�(�ٷi�=%������;zĢ���5@~g��"mF-��i$�®��M�[��(�ͽ��>����L{�x��W��6�s�olOfS�~��] ʸes����� �޽�>ȏ?� Wח	�-�����gys�'�dY�,�>�������L�*��l?�q�zx:��<��t����D�PF���f}�3;�4��`�S������1����7Grqq��5��?�!�a.��Q:GƲ���AP����Q���3 �z��`�؞j�>)���[��KgJ��	�^_]�^��c�lX�n��%��.t"t���Qy_�q�4��5l�Pp]��D�C=��7}���� �D"A��fT0��ɍy��_X�2(0܏���hL�QCdGX�Z-�=�/�b��<;�$�<��jYy��렮*��$����*:5�5C��m̸.�5����$&Ѽ��� ��t�r���l�.��ʠ�O���n��Rs�w��R뽇�4V̫�c�{��B�l��l��Iρ�T�|P�$�ܷ�YDc,r��nX�1�cY��3���@!\Aaw2sEJ�Xϡ�X�	��k���&T=(&�F�21�q�>�����V��6_�Q=����`}��[��9��\�� ަ����s��n���X�E]�U�o�2|t�H�7K����h�\�=c�c{��I'FO$q4�yw�>O�-k�l�2/.�2�ɢ3���~L�y߈�C��\F{�;�pw������Tժj��l~)������_;4�ٗu��0{nP~�f��6+;P�:)䚚�ܼ��S����x�p@���lbTL�ӡ���z�k��C
��&'䂠K���[����p0F/}�_�@v����8�X8��X-���G�{�����Rs� ������d�����k�J>��Py�]8���+B���
�=��'YV�]�2N�]p�?�R_C�}(�Z��0̽q�_3������� dP�0x��iq�S��I��'�
���}sL���ь�q,�
vߠL�S�e�>Y%�pyy-�}�}w�Yޓ�����n��C�s�N���2��Ś$�����~5�֧�O�`!i��	s���m�s�b�:��Q�ײA4Q�����Aw���/T(��A���R����7r�qD��Q���@����O?ɧ� ?'�9S�k�uZGU�m�'�Z��3���E���" Vy�G \cu�N (�?@�]Q�v�pA�Rb
�K�����,PoJ#��H.^�o~�N�����ߦ�o.N�X�ό�Xt�O@i��;�?�»��C���`då![�WOOO�u#o��Uj�L>}z/?������q�Y[40~��͇�F��[�?t��U`���{{-�˜ʝ���eߣ���B��@�KjPe{$���"Sh|臞,�,����,�9��j�qKVE�##�?�=j{u4�N&�ز��H�۵'�Ғ*������[���b:���U�BN59,��#u�s��GD�D�ک�=z~UG޷Yn�}��j�pcaSGU�~��B7?ߠ�L#u��^�"��z;-��H{�-�J�L	�k4q��.	��*U��%��hnx!evk�}�ejH$�#����6�h9� �.�mzo�^l���>��u��k��6k�_�65�V�|!Q>�f�Z61�벘o*�p����Ҋ`[�-%�jG��͝���h�g,����U
�^���2�+���V,���9X�ףΊ�y.�W`�wq�W���*?m{т� H��:* �xG�v6�y�p&��帔�]6E���V���^�ԝ�7�歾>�Y���A�a�mshÜ��p��l��J���f�!RP�{b�6�<�}&=r
�e�5�,�8�Ep��V#�PS&�j�w����h�����
���t�UبB�Q5��F���|�y�A7 @��G�iB��=�*ܮ�5�N���N4�^��b��I���Om�"�r^Ы1�P�dr�: �N�aZ"3T+�8GC8���ԛA�8R�����y�x)�O�z*����~-w��.xO�t�]���Q�{x�n���	�o�M����K#���5��7��������,�n�aM�
m��#�ðj��s�_��jP\����a���5�>�I�X1�m����,eM�HC±��>�FV����:玒4�͈�5����|�iԵ
��Cͻ9��s(ӆZ���F��wy�	s��s���ó�n&K��J�{D#�T�,�,i�3��Ԛ'e?��䕌QȔ�ǲߎ�pOi��x�6����jfX���g�Ʊ��Ψ��bp����?���Te��.2��BF�D���A�̓����Ꞓ��iN}cO���W��Sրl���$�e�b�^�˓�,;RD%� >���H�d�)5a���⨕/���n>��Ҿ�tk�d����7�K`�i����Õ|��`h���/���y��AD�M��*��~-�ܶl'���#����\���PB��@�$)�(�~vr��rƁ]&/ �2��vq+��#��r@�d��gg"�{�̔�k��D�E�M�Ԏ��,t��@w�H�ZN��Y�
���EyLJ׏W���㍬�	T��2> �&j���S��y��A����r�X�f�g.�."��*��9��a;m�X���� ��0��0g.���W�y�=�����s����_����������w�ͯ.�w{���\9f��&d���=g�C� �7=&�O\@Ο�>��7�ҭۤ��rz�ʫ����9�o��&�m��2W����J&���x�����xȚ��d��p��(�c�����D+�ϵQ#n(q���3P&j$�h:�I�5M6�#�N^Wvo�W�U6J����9��t�N��a��)Y,C�\���f7O{2��}����������O�wL�K�zJ�5�:=/���e�p��^��!*�;fT�{X��H���Y���X�,4<��q�a����.�õ<<���cZ����_<�������B��2��Vqw3�C4g�N=:��219|,Z8���H��Gc Q/
����xp�gG���Cw�#�(n�S����_2��2·q�O���/U~�)6�4���w�t=q(4l�+�>fv�����0*�E#e�D�2R���'�k�4����,Y�/&β$w�߯�!�;��1V�ە��|?�kq���$�0�yr�c��e�@V�L�u(^NS���Ub����;�k8^������Kv�Js�j+��1��s�r��u��J�߈y?x�r<�t���;\���h5�՗�LU�$W}	e���֦����5��{�3�<!ፆ󕰝�3owa"Ł�v�rYX�{��I�/�P���3,Q�xxUp���eXZaA||L��ݝ<>=�y:<%�D���R9���:o1�����*r������k�Ƥ�w�<���(�lD@1�Ő�h!V���z��+�����,R$�S.*Y�H���?RG,��a�()��g���G��;e��K%)\�� c �Y+��ђ@V��՚FѨ��2W�!���Y��d$��?����́���XG���%�
��'��3�v�[�5	2�qPJ�8�T=�ai8cA��	X�I��.��>�i9䭑LA��`4��&)z�Ղa�0�b_�!)���̩����H���Vn���X���ͽ�(i�Xm������XE��5�:`�>#z
���*���l�7ب&o�@����e�+�'k�������n)r�@� �ԗUR$�Ifд�A1��
�y��<�-R{`.4��ʰ�W�2�b�)�N:͇�;�2���e�f��$ܓ�s������L�������N>���D4�v4,DK���IY3�^hЎ�1�5޾��o��R~��o��涏����}iMm����Z�S��іƛڨ�J�����a\k&\w�?lR�^���u <3��Z��Ox�	H=X,������,��O?2��	-��1�����zNi���u����}}/;��?���X��"���\E��pb,pf d��	M�X]�)�[OX8{�\8�*'YĚj��1��Z�q�� !��|1M�u�ɺj�_�Z��*��^BYѓZ/uCQ���0Ya��2�췞��@�s'�7�Ck��6�.�z�x�$��7�>��]
 �+!�ui:
��t�kڡ��E��a�r�b����x�+?�|�`��>�aط9�6�:UKuŚU)�~�BibA^~S�K(�ޛV%Sܩ�Xa�h�'H(e�B4�F�w�Ӷ�?��x��rc*厀���f4�l�U�6>�l�YMY���"����a���U�*{�=T�&Pպ&U��L�J��C��C�ߒa��ئ�ƍ�'���
�ʂ��yT���	Ӷ8�k�h�A���>Ժ��=��J0�U����~��������2�Ny�D;����B*��0ǘ���5Ro����qXkNVk^:�^�5��5�����G��sP/r�k-�����8�u+۠d�G��-��{&�����_��Bf�y��|�e`��j8�UP��x�fH�I����c�{�o�jͩ��Z�͚LVL����h��M:+)����u�4�ۓ�=f���Xy�����d(�������!(�E={��4Eb�>�G�x�60�@oD-;M�=5�&�YRz��Y���	�N/V�,6�{<S���j����#�ܘ��Ł��Hhh��sn4�>�~^Y5��
$۝Fꔼ�rj9͵��w��@(0)�#C��7KJ��ɉ����L�VҊ�z HMo�3*��td��b:�	�Mh��M�
{N���@���#Î��,�kG�x'f$�h-��4�!J���@��r4�7��%�V05b�}����1-���	,��X4 H�r���yR|/ ,�c5İ@�ab���ZSG,�h��W_�J��N��I��Aܓ�˳c� ��/�J9ˌ�y�^��atv._}�N~���"���ޥ1=M�="c�O?�(�^n.e�|�w^�Q{�c�] �#�ـ��&����w<��>L��b�"�Cb��?����5��7�b �CdD؞�7�Q��FI��~Hҥ)ff��߻x��JL k)�g�H��T�ʺ'J6�W}����Ϯ@g�z��Ld���.��d��������)�,�J�e�< �����  
}�f%ќf-����i-���ŝ�K�p}�{��i���ؗ=���i�W<�g�'��5�	��P��߂�c[	��(��H59��3-�/�0�}���F�NɨGK+ɏ,sg�/6���p	.&#
3�-X9�qC7+����C�D��g�2���w�6i�tʊ���8h������@+2i���{�x����Y��I5���:H���jomk��ht��GK6�uK��w|nj5��e5�����
~�Qd�i�g-��R��k�a��J��z���L �0��)��to��"z�BȞQ��w���T�ԁ�)����Ӵdo��`��벐*JuVW0U����{38U}v�U@�3��2�_u{�>	���U���� �Jm�w6*\꿘W��0�`ޫ�I�����s��Ǽ�Q�Cɡ�u冐�8#����ӳۨɍ����3�փ*XY��
��N����y�L}�5�L����z/?~�o�-�l�/�E��y�].7��]�2��QQ����?|4�Q�{ F�����R�Z<&�fE� ���Y�:,�NMM���jg񠏵�]-���[&籦�"��D���Og���O���S��u�\C�8X�޵0b��{EalX������=	H
P�kZ�^��͕��w��z�֯��|/2�|h1��&?u,�� �V�K�6W�^k��C��k*�5���ԉFkoƨ��D �@�<��Ue�I<{���o���^ߥ}>�ER ���Z6D�P��t�@k�'�z,g�G�љ'�=Z"
`h��}��9���B��)D$x��/� �j��m����@��`/�ZW�Ր������.��b��e����q����C��˯��w�^��z�z��r$g	d�:N@3��P���V�>*�5�r���Ǖ���R}��$K@� ��Z7f��Diӡ`G�����];9:��o����{��39??����i/77��� �����5�2p5z�&%LiS{�A��2�b0�kޒћ���`��>�|t�m���YZ�Q`'  c��n��t,�w�c�� {z��&̟cI[����m���^z3d��8�S����2i[z����8+}��vʡU�@��g�+���.�o����w����,��A��It*OV��6i�x��2dN�e$G>�����0��l��ԅ���{�u�J�ƀ�3��2�\��ڜ*R<\�g<X�$��A_)Q�OnM���)�x�T��5�Iw�`���LP9�5�����3Z`���SC�*q��tU�G�וk$�񜰟Tr�B}c{"�{� ���$c���uccYY��u��Lc!;I(v-Y�4^TA��	����5�j��*:��sn�(�uy��	�(Y��	����9��\�gm���+~^�������m	�6�{Y�����%T��?�>�J�����z$,
kX�T-�/��|��E)\Q,��@sԤ烮��{h�d�W]��tJP�+��W�fj�/<|d�����e��9K����91R�Ɣ����'��/+������8\ �g!Z��
`�N�I����"����@����3ZE������Y�P9�vF���~ƃ�xP
�O �����^�G�aT�ω�"CPi���B���Ƹ�p��E�]7DTb򸘂���K�d�mRv��p+������(ch�e�Q��ɞƼ�=��[��d42B��|sH�&�jΞ)��f>W/��3�c�?׊<�v��fE��Ai���k<"�8��qt��$C
��"W��i3�{'���_d�k�B�V�`jh|��;��m�ˤTo����0rR��d:pI@�ѭ�kxOj9+:����s9NO��AV���I�ۛ�o�?����������k6-X�
`LC� N�g$�8?;���T��^�o����^��ޱsN��-��n�тl�����崵�f|�˧�� �r _
:��h�(딂2}Z.7��Ӎ\��Q!�q���	$ _���/�x'�߼�?$�Y.e������Zޤ���0cn<J����H��ۥ���VF�O�L��(��{#��:�a������0VG��[�z@O����d.�|������;yu>a�M�݆9�����_>1Dp� � 0����<�Qt�埂�vİn�>(Ad����g~h��v��\�+�
ҽ�62��|�9�0I����󮎏�i~&2M�7���~GX����\~����dR�bt�re���5��Ѣ�	��jD������)��Q��)(�s�XL'�|S=o��<&�$�R?'46�5% x��Q��	��f�2mS�'��5�+�۫�S}X�
�}����[��Pi8!�Ź�{e���AG�����G�!��\,.�p���\W�A�~�ĻJi4>K3\�Ƕ��v �� b�k\1� ]��9H0	P���::�0���B<S�� ������M�Pe�<����Z7/Ԑ���wa̰��N%����7&��X�~�D�\Y۞M��L�k?������Sj�L|`LQ��2R0���-��`�4��Fr7�/C�"�s|�W������<����ǮR�L��m]y?b�->�o4>G��J������Qj��k�؋���"�Z2�Cs�B��T�\*úQ�w��z`m)K����B��m|�Q��S#8��o�h�?1�W�Ѡ��gJ�����P�9}��2���%�g"�	��A���&{��e�Z�`��Y75�B��
���52Ku5�Qg�vLC�<~�C����#^��'�?ؾ�+Zf4c����[�1����4)�٘�#� ��mv�%妏u+Wt�ZیN���s<^�|�^y�&;�O����6)(��
��Q���ljn����CI��X��j�l%'3�b��a�A`d>�W;�����2�X�����=�:%d��� K��cR�"�«�I����O��+��5LT�(m#���f�����/Ƀr�_��3*�!�Yٱ]� @�S�wa�,ӛ�[��Z�M#O����#��`r
v"����˫�9{�J&�#l�J���3���'i�_�]K�́Z����x>���S99J���DNX�B	�է����&�������X�A�@B�^k�\!�� ��Tka��S�	��=$��(�t�	��O���kh����Y+ƞ��ܟۤ����G�:�Ӟ���r|t�{�����9uJ��e,��E����C�h��0T��S��r� �� �H�͂�
�X3������:ͽF4AO<M�%���A6�4���(��4�g����1k�����mMn��M %��i9�c����C�ϧh���G��q�k�.1酞L�U��J�'���i��}�_}%�/X�+�������R���#=��g��ka����a�����S������Ԟ�ݑt)*{54F�=V�> pz��\��K��dG�o8�I*/��h�l���]�3�(z9�P�.k~D����''�;R��3�9�~�
��TkP5Z���یJ��A� * ��Ъ��{m�v�8>����[ZnJ���JE8㡒�)(�\��sp�Z�s�uؠg�=0��F̛�	��� e��	������%�,��y�Δ�>��U~��ؗ���łoy`�f!;��?��X��8*��Y
�-V7\�
�pw���$�?))�g�,��.*�&�o��]��/ K�W�kb/����0+7�3�eJy�و�����,E�Dܙ������5�B#�����ӣ�9��ٷ����b}=��*'�&ThZ*�g1Xڋ�C��Y�N�C_���x�o�V�Z�ý�(|8f�B��p��zԆ�C/w��P�7P�۵q�z����K�	1?�5�Rċ�r����G�ڝ݂�u����+��K�S�3WD���R�S��d��rz���Ԯ�7�[�'�(��&�U��5���}g�DAs��Y�-$�B�WG�k;���Y�{Z����?�#k�̎fr܎�1��<�qQk�dW�a�AY�C9����y~���fr380L�1)���y��'*�Z4�	��1��U��݆���jI��E� e����
�_� W>�\9��.��a�,9?�����A͟�/��5}d��g9����Z��i�&��r�&����F3�G#x"���5U���$�g:��-ʐ���i4�W����޾�[`-��d1�U
#�57���`���%߲v�/(�s(�� Yo��$���1r����{�.P�W�/�,��k	C����<xg�����G���ݠ@m��O*�؞���"9��
!T�ѧռT|���RVoi/�':v
�x~F�i6hs-����� `�M��,�o^�K�$�8>>K��1�
/ ����َh�-_S�����g��q���B�����YS�7G�N�x0ڄ"�#*��o)V:�p3�G����ǬJ0r��^%y}BP�Z�7���P���b�"�܃�����g"%�Co.�X� �yO���% ��Ǐ���^�>�~(~@Β���G�B�I,.�|��������@�>-���,{�c�TAꎁ������I���iP�{&j>l�w�=fG�pg�Cyk`q(K���>&zG6�uI�#�y���>J�dc�v;b�=滟��`�;l�1�3򭐃�{5FD��!��s�f��<�~�ެ�;��,���EoI?�/��7�Ku�X�Jc)
b�J�"�3���G^U:[�_R�����r���������� u�i�1L<6:Ыc��l82zd�:Ҕ�u�L��Ǻ	�<r1O^�N�z\ko>Z��yp�"���=�����Rɒ�;h,n���ٴ�S�j	�di�� ��!�j��W��݂"��#�מ�]���i(U�y�Vot��k�#SP=_N�!Vĵ׶�`�����2h�Y�cp՟�xs줮��+6+��AD��,/)op�g�UDr��^����u��1�T�����
B�a1�9=��byǸWqxN,1����E��vą��n>�t�wQV��Sb�Z=�ҟx8�
!��^ת�ƪ�?w���HV)C	��P�:$�"r�1�G�c��Ɡ[�`�o��>:�����nJ��*J�
d{����� i)��#-҉뀹�O�==���lF��uzz*�'�L<7��,�ю����:Gݖ�?������w_^01~2�Qy(�.yϸl�	+sg�A��#�+�|�͝XiXzb�
�Ý�\_���me造����r�D���Z���l����k_��T�z�c^�zf��c��%�`ya��_��%����������s�s �c)��&�Ɇ^��!�k�Q��=ʇ��$�e��sۣ|�F����Ϸ�s��z!@!Jƈq��	�{������5��z��(`��|,�{Y�A��+���P=��,
��숄��w$�N��Ę���	"' �w(8�$Y2&��g�S4���ig� 툦$���Pdo��f�8�"g2�ڇ�ȥ���o`l`@�ӓ�ř��.5�vX�vJ�C0*A^� >�Esgf�eԨC0�	F��#�`�tY)�`.����<z7�u�$1X��+r������H�� �� s�^ш�hy�hc|�g��K;�m�caX$�����rz�f�>���o�0Jj�HV���V�Қy��ׯ���u Y�|�����OW�';?U��W_-_|���J)n� ��V��W�7������;�8�����|�tGO�(,xl�>���2�z?~�$�;���h����� �C����:gݰ�x]��oL�Eux�b3��%gg�G�d���þ���6�ZAp5�r��Fn��w�c �b�5��j�����S4�u�-�/�R%*�>��T�Ò��@�8
1�Ө�(����de�ʗ�5���ڞQ�;!�8&�C-<�Y� ���+ �1��F�샩a,�1����$��8���jlU'���/�]�S�*A�'��5Ȓ2F�q-�)����	�9��3к4e��HO�Dkd�ᦗL�7Qť.��Zr�hQ>/�G���h�����/����!����c@�9s�G'^-பW�BY��~o,N�R�Ǭ��Qr�hu�Zz��uwF���=�y}: ��7fe�=쉇��G�[gd#ѭ�ʤVX�`i���89ȳ��lr[@Vp�� �d_��"y�*$��j���1������*){V]�����2�v�!U���]1� ��f�(�6�Q\��aƕ'�p�R#���ǝ����-��>�'n���K�6�PCE�5ގ
�~c�)X#�׀�2��5�h��i��I������׌��9�CL�P��յ���I~��7��_��ٹ#�G�BX4��-�j�����?U&���>{�)��=XA�lq���
����;�������Aq1�����m�� ��t�%%wI���p'ԥi���`�ͺmul��)�C?֋���Gm��։�=~�W�ޭ�����
�[4C�<���}ь�f�L{o-m7���`%�aa��zPy�L���?1��o-�F����l�v$�����L���֘���#�o�UfAҥw����T�K�I��1��n��#��5�x̢��u�h׃�עlF�F*(�:z��$P�х}[�5�̕Idt����_h��+{Z32"3\t;=/A���H�E�A���e\�</M�%+2�M��HI�?��J����#]O���C
��}�Kc�6!S�:�aoN�ѩwcЀ���W
a��nF�m��"�1��}oҪ՚��j4�Ԇ�r#�%B�P�,�Ó�t:[ߜްh�%�6O�pB1X���M-��0�Kk�2� ���$�'c/7�|�Y	=>�-�l㼾{Lkd�Ί1�Xk�浣�Oruw#�u���r	 uMV�h�����2 w���k詚ع��=�:)�(�E��}�.��`Ώ�̋�ά,�*��	~��;��}�]5�L���������!�, 
��h�>5��z�1j���(��wv���_�Wٰȫ�{�_ڧC=G*�� +O�uɺ�{�X��6�����*�U ���ˊpA�٥�H8�J��V�u� �m�jɬa�M0���� Kk.��`�V�`�Aw�o՜��GS%�-��~����[~A�}�̋��P����@ dEMF��Z���<s��,,�`��fMH�̮�G���ݪ}Ydq�<��4�(2g�qb�\Rj���.�h +�5	�l!�vP�A ��{>TΘ�W � �Y<�t`L����{ȣH��)�g�l-7���k�uS���㡟�H��5d�h���zb�XzH`*#�؁d�,$��Lo�'�v>�+��%j:����u�2M\��g�Ԭ���|�2DJ��T��}�j��+��Y���]��2�B;5��[�9���ql��a�%�j�x䣇
�'T`lokB=�m��j$����K �.-��_����h�����z}�C6K�`2{H���O����r}{#_|�s�#�1ךN]<xݻ= ��!~�(��RJ����9@L�x����9n���N6��8���D������=���uR��i�V����^e9�B<��D�X7�V��Ó�t������:��� �,�3f� G��G����:���Ѵ֘��ؠ�G�#d����vȫIj-,%�����g;c��V�y�<Q�YC��Mٮ�4��d���ub � �(Y�X�F9�<:'���`ax;����߿OJ;��N�͛S9N2�r�WEk���}�7��u[Z`m�gp��͑�e"�Sk�1�o��������X�X0O�������i��k ;�r��k�����D��cPe�ۛN��>Q?@�ℹ%�#G��i�1-(�k�P���~��X�S����rv~.g�@5JO�:a����$����i�$`Dnh�W�9��t�2�q2�indg:�7������X�Z �N� ��e�d4#��q�c�:־��i�D-��I��So�����W�:�ʌ������ˆa�;��gD���dƼ7�؇����'�O�o�\�~��&8g����N��2���j-���,�v���0lA�����G3-!����QG��nZ�T
�ߎFD8v�����$��K��������ܱ1|��ɘ@�����u�&����YL����XT�댝�����(/g�Tf�^?�~��V����E��\��Po�Y��dtYm	�"��J��x�;�Ԏ�F��Ieuê�-����ԏ�x(��k�@v�Ec�se!ZYA @:2� !|�Q����� ���=-0�����:�[��ڐ�f��PO
Q��!���YX��Mg~���PA�&m��V_綞�Ã�ژFtRB�g��~EM@���E$��Y�oo�I�37�"��� �Ӑ��AZm����21c]4� ��@�����%��%��}o��.*?H��ih=�DQ�G�`��z�t�Zi���|����	7���P��ƽ�~cnom�`���s{!dm�N�gfx��2�zX��m_�*��Lr_�h�Wl�ҏO�2>I::$���FS(�G�ux�����s5�`��ƪ�m�k�!��h�����0�R��ԍr'*� � -��$��������F�^�b톔GC�j���<b�|�%��AaJ����ێ�R1�Uz�Vci�Z6����������j�)�b�!�i��iR����c�� �%��	OOw�\<� �и�zQ�d�'�������4�w8�Qc��6) ��6��>ȗ�|/�_�!+ֱY#Uy@��<��H�!{��-Y=\����`I��zJjmLqǫ�D*[ht�5gskY��$W?�An�/�y���1KWt��i�xZ�P:�$���; K3��rq/�~��|��"��,�팊Q^V�Z6���iB~2TH�K�f��D�L��G��C��g���!&��S�,�W%�����>Cb�4)���!i��k�'=���#�
����(�l�0�>�lX��d�4CV�@�2��dY���r����]m�'�{?��dn��*� Hl���I�x%��KY��aƈ a�7>�QY�BR���'I	��r�� ����x��Q�~�S���N��S���^=�o��Z�������9N{Y������c�3�*˲�t�uG��N���w����$2�
�	�%��n�7�C{Y<���pN2�����@�	(���4��ӵ��m�t^���/�ի3�w�|���9C[��c�,�� ���T {�ў�1�,���C����s� l����i	�.V����å|� #�G��g��\�s��z�@g�޸�SO�;�{�c��W!���m����}J��!]��������ߧ���K�Hs�	C;�J�pW�Ñ��QМ��,0��Q��J����0R�C$����e��IZ?#��mǒX��������|H��kR�dJ�k/�٧%ϗ~�:�>�J���	�p�����;�:�>���Cc�3Y�b(�(����喞]0mB�@ݠ���w��E�pGj��]j�4�JuШce~����b:B�3�qE�S���Ϡ8x֘#c*c��E���^��⌢�6����*Y�}�4E��x�p�ʮ��>Oل�2B (F1i�o�Z�9C��&�7r�,�jM�:���2EWD�ZFe��f�!<�d��Ж�\h��,� �=��9,A��d����Ԟ,kB-�eGo�J��
{���m�W�Le��;�\���Ў5!3��,VǑ4�lO����d�h�i$�fE=Rm/:��1���`��[��m��-/���g�V%��UFB�3T��4<Ӂ�Ȫ۷7�U�l���%E���N�-�@��Hm׾|/:��x� >�!��2�ޥ=<,��B�9b���>9��QC.ԫ��%�g�G���Oge]J�Y��|�z���^��s�����C��nL���D�ޢ�E�{�Z��DP���t��P�r��,����y��f�
�l`���'YC��^�Qs����IO9#QC=�� I%�~_%E��q)����?� o/^�l2�//.Ȭ���[��u`J9�*�^�Q�,�U��f�\�K���ZQxQi��֍-qOF����Or{�))��M��>�M)�<�s�/2��v��?=0��/~�[���V�ŉCc�AZ�c���vU�����j���/��g�����P���^�{�FqK��ɘ@�zU�A�Yx,�S�O�DMhh��Ы���;.���`bƗ>C�� d���@�$z=K���>��#�
m��\,(�0 �[5nԣ�F`��Qyt�K͙a�Lg��x�;>e�5�������#�2\]]��	]�}��!o�>�{)���Ч���;y���܀8?9�S2���^�W��R���O1G6�=C��Y��L��p�?��b�G���E�Tj0�}�wU�g��A=-Х�8�"�0f ���tnd ��������K��j��ʫ$�޼���u���V���������t}�~����VsZ����%i�8g��'AGd�1z�1��f�?<��?�(�G��b��뱜��bN/�dŵ�S�J> ���۵XƣZXn40`�����H��L��1��6��n��q��������_���Γ.;���ݧ�#���Qc��J]���,�T�U�ҁG1�����z�Gj  ��L�g�P:�k4:�v�P�T^��J�ZO)����$R�"3�f�*��r$������v�)+��&dpϒ��M������I*�ꖍ�y{�z�ٸ_]'XJ��M���1�0:?#�/��U�H2x����k����R����sQ���>�V/��C�љ%��|�>�����m���AV5de +�L��G�mAٙ�����刪Vh,�<=[�c��'��埠*L=�w�0��j����vd����z�]}sH�Ƣy��a(��1�;Z��CX��X�o���dC �ʭyC��Lx�Β��ѫW�59�1Ss:w�{B�3�Y��u_��(�Ȗi�co�jP�ﻸ��`LpՎO��;��
��F�Z(B���Z u�>��}���e�>{��@�.�b����=8�
�T�?Ǽ�F�J�BSR>[���ʲ�����!�����ُ��s�������x�گe=�A������LPj�PC6*KX�=��
�f�3?=����Q����Xv����I���>���Q�A�����[���[99>V�x4c�#���[I�_j��%�0G6�Q���!�)�F��mR��t��=	/@��1Tu�ZV��J�����7KU�4x|�';�SRzQgJmE���l��Wh���z���?\~�1.�/e�����մ��$�x�smŦ��j���@$!����2I k�r� A u0_!��<CIk����Z^�(�Ԓ,+��L�S��I֋%�= �6�-����Ez<�86�e�$;f��fC��@�2��eRV�PO쁹D
� �9k==.	�v`i�mx2����,�#��u~rF��iGP���B�7��>�=�9��%*����An0!K�\��5<�`1omϜ���>]ݱ�0��jo��N�Ӡ	��A�	�Q �	p�;��K$��#���uYwi��,*<�p-''XGaz�{`�O�@xd�V����h��|5V�9�Q�
���!t���E�l����+��#�����o~�M�cQ����bF��#X�SB��/`�enb�3ʹޤ�}
�j�,�nQ���3u|���F�JC��w2���c����rys#wi�m-���D��&T[ɜ �gM�1�-�fyBQۡ�u-�4�>Xy��92D��5j�vc
Ec$T�6�����a ����z������|�2��u�"��F�����d;��:CE� ���58*z����Z����D�^�xf�U}�ڥ�E57�T���7i�G���F�ߠaV�
A��q�^�P&7�h��ZI4�L�z)t�1+�,3����N
s�)OA�u8I;\)S�%���&%	�o�z�$HV�Ռ+��&�»bQ�<.`���U�eNJ,Jl_y�
�k}���¦�Ձ�(8&�Q�ɼX����Cs�%�e�)kC��ڃ�Y�UO�g�*ZM+�����k������ d�^��ܒ��0��v���+��yYM�j�Gi=�S@����l��;)!Lk�F}��H�5�o�b0�]'Ŋ�ݏ/�5�w��>�Q{���X	�X�<��h��yͅj߄"$k[R��\P��!�;��`3;�1�g1�r���!�[�&���)_�cdy�b �[��QgV��dJj�)tP� (�x��jp_]-^�����\]��?NZ�FBj嵐��^�1�O�=���}���E�á\|z,4,�}QY+z�7n�{�Vw���-�t>]�C�<�>���u�'j�b��q*}�r,�yhf�h�ہ� ���yR$�R?��T����e��g@+�����/�8��,��G'~���%Ca��dm�J9�`��D5�� 8�8&�a�&تnWOOu��,�냴W���B㠇���Y�2�р�:���K��jϺYA�&�v](��� YC2���.*�Y�
S�p��a{`��W��� s�-����\kH=>>I�^�N��J�ms��Qa����	Ev�҃;��-D^s�>��O :�4����Eҋ�I�-)��K�'�_ǱQ�4=�c�1��
�x[��H�0�iօL�%P̻Ҍ�$c�щ� �K����"�
.�<l	ܠP�i��d)-���x���ӰR���ݫ�V�+p\��7�s4�|
������ �Bw�e�"�@#OOVo�e�o����I����� �2�	��EM㱮V�
��Ҕ��zIY��w�3M�Q�U�_!'���Vn���Op4�E%��9⥅��A#.2Sft���oX��H��4CI6�$�
�zY ߙqX˶(�C�1d7�95r]�X>[�|�|�3re�1`����5�_]S� ,���J'��(�͇��秗�%׉�v>�J�E1ÌEtl�s@ϲT#'�Q ���q�2��C.����#Q�W;I/�DB���m%|���� ��E��b�Y0[�
��
eJ,��z"�

��^C�k�.�:�����}S&v 4�T+��=%���0]^$��:��z��luNޥ�e�m��zo�?~��"�z*�H�Es��hy*���r豫�R�^� 찊Uݭ�qׅ���b�y%�V����T �>���钷�}����tM?k�	^�ږ5�a���Ê�{Q�Xh�IQQ����!�چ-B�	%t����\Qn𙁩��Ց�on���1�UB}/W/@�h��w�����G^hq��U��A���l:���J!�#+`��Yإ/�vS���������˄.¦��;qr*'ǙK����ǧ'z�������D�%z昱�QA�c�ɧ��|�x#S(Z�F�G(���$���v��Z12:R�����ZݣYO)/���k�\�O�W�JQ�n+���m��+���r�ӏ� �&���AA�Ӈ�tDj+�e[��{�?�8���Z��u?~�Qf�G����D���hU%;XA 1׋��O/�?��_�[%|�*#bQ͋#B��IY�W�!)���� �G��uR�7+M�'�k�"P�sm�M&�����h�9hC�T��� K�൪x�&�P&�f�G^��d�B�����}z~d遮�0G��-��Q���ހ9@�Q/3f�Ѥ��Ë�5��2ax��A�Z���7̉M8d:��~��t���d�-��d{O�,�e��z��G�B�A������3⼂�|����6�Ol��K���v��j��8a@��Ϧ�{�QBX(J+`����������ҲfӔCL��!�P2���ʖm�FJ��h��@Ly7jC�QС3��H��{<�џy��Wgȕb�$c@�q�~�Mߙ��N`��z[dzt:��g!_���0��k��#�$+C�����#�z�F"�=�!q.	o ��цm�\8P���-jсq;(��v�f��$����rpݠ�gpc��X��]������T/w��:+^�kx�~�<b)��+���"]�-��~�l 0LN���z������E��T}Đ#�>�p�&;����ϝ�5G���}5�B��x���i>�As�+-��r*�F�_�2˻50�����sS�-�)/z�|��l͚�kzᮽQ6ƾX�5���I]�~;����
�L���Dπ��`�?��kI��K�t�� ��+��r�nw��S��0�׌ʚp���@+�f ��}(o��bȎ
�D��=d���4��]�Ԡ��J[wb�"�G�WW���<r�	�[�?��u�4!�H=����lK�X�{��N�a��(�ZQKkd�;���Ƭr*�bUʔ��^p�^p��ϏO�l^��
�_������}�ha���O����U��	Xe�8�J���hD2��������1ꪜ��,w�o���N~�(���1�3�"'�]P~�`���ф��P��Ia��NW�.��Z��1�V����I���������$�]���<)�����_������t��
-���#���i$d�k�f���{�22j	���()a��Gy��N����d���Ǐ��O}��;W֜ib�w�	�d�2f׆�$� Zz���O�Y��ݛw�+�˴��((ӗ��=qQ�pd�%�>(���1x����C% �P��.e��g�H�I9���lX��Kk-���Ձ�ڜ�}݃��K4�gkAC
�Ӗ�Y �C�ֽ���)8�SI<bS�ŭ�\�����o/�x�v��[���=����!ȁ�p0�1�&:�PP6�`FSx��Q$�Vhy�&�u�}�[$;��u\��Z��F�R�VB(��Y��C5���9�q;M����[eDM'��!����u.�,�M��cӏ��b��Y8}ƐA>��-d^���m�d��'���	�0Q�=r{:%�����i���3�y�ێy�0RAv�SwO�i�iabqR/Q��+)�=�%�@3�D;h�R-=Pf���#���_����,���+]&���EN���|�F�>�$���L���>h0��
����g�t��yQHР]����6��䀘�a��X�FZ�kE���h!�n<�����$���}�n�����b~q'ZC�ɷ���(�ޢ� �J��{Rk���Υs2Q��/������\�h^���𨑲�k���J-�nkMb^�9�tmp�a�9E�%)����T�T���(J��%�B���l���\ $&�b7��(���0
t$�y��M�+�x Z¸���[��gD���Z[Bs�8tF��(O�g��Xy�ie�e�	��nJ�u0yjas��#+�W���P]!߯b�z�g�:�$���b�k��Q�y����,�l�J���|��1�'[�?��#g��Fg��u��i�t�.H�M�M�{�U��%m�K�_�3��q|�s�)s�����d�7��\X��m�Y�wO�|L��6h���J��Q򁪞��+�{�L��6��@����ӱ�X�t��g�9{1����X_k�X��p�d�{˃�['�l> !jF�Fښ��aX!C�Iu�p�������Q #\�A�0�зr8x�,���L�c�s(2�i.�����
��P!�W_�Z@i0�M��"��������x<I�DI	���}.g'��@Hm��L��-�޽�bʨ.��y?M�pB�Aq�� 7Wrs�Q��Ox� �����B�D(&�1����	��j�v4>�`T��InT���-��ЬO�.,�=_#�5lD�p�B&[�>/1p�Q������޺y�!�)#�ޫ��4��Z>&���2H�
�S��2� D�����0���h~��h�_���57AB�(~N� ��)��g�Q��;�e.՜fD#�Yj�V�/?������CRr��X�!xZ���cڧȑY,��f��m�:L#T�5dh�_��dxr�d��j�b�lbe�Vj�u��v�&�
��3�O홐d!`�����]�^Աjӵ�@�z� �f($1��O{gQj���s��D��}0�s����vȓ�q���+�a��(?��v.�fB*x��-Uo�ŋ��E�ݎL�{���k�����=�*�4S�	�:(p�|z�{GH�`��׵V�!�2��FQ2�t41�5���t.��_����o�����L�[ 2X���2o�^У����vg��U�g2��pi��ͷ�@����!�Y���F	���8L?N��$��)��M��s�8�Wg�����$��M0J���b���$�b�x� ���k�uZ�)�|B��K��L���k����G����o���� +Gx�9Z�z�|�{��<xA�U�"��;MԞ	�|v��?Ti�Sn�������qP3:�wL��P(������+ �w�K�j\AV[�,osV�=T�S@���.��YS�|����,��9�/�l�#��C�D4�
�;��IeI4��N��u-�~W<6CI^��j��SR=%�p�O���j��y��{�%�l��1Z�j� ���%`�tj�3p(�^{��7gc���P+��o��?��ʵ�=�_�i_,yU?j�s V����ů=���7�A���.\5Tm=xfi?2�M��@��Ec��_���;� ��B �(@�k��g=�D��Bx���}˵��Ù�}���8�t�e��!�p2�M�����3�:+�;ˋ�<l��s�"kȴi}1TЍ ƺ���b43����+��=o�nw;���ek{����Q�9t��z8BRZe8��F��h29���0E3Z���X͞�����|��:D���=�zq'��g�廕��_0|I��dFO>kE@1��+/�̥&�]D��슁V�'y��%!���%Y�m�'
�.=潩���=6>C���F���GԶiJX��2��a=����t���S9;{#�T��F�}�fSGYL�e<����y���cEn���K��!�KO���6H"n��Bi�,���Ar'P�K�C\j^BdP���L�_u2?��"��a�־���B4�|+�<<��}c�\=V1b=Z�^@֜Z��]Z�W���G���1�����m�ߚ,ߴ]5A	�@�p0݁�`��1}	����y1vc��������im�=��N�fu ��NUqF_����T!v�9�5a���=�'���ab�YO]�z�4�Al�5v�FO@���������wV"�̢��Z�A=���9�.ʾ��1��pbӆ�!��z9 P�&ˉ�{����y����}�1*CZq��Ȋ�SY�v��n*�.�}�D�l� F	�R[v����1;?�ɯ��B�귿J�e"���� �4������� uJI
��so -����czs��6��I�bL|dP�L� ��M9���C�/��"�|6��Ԯ�E�#DE%���酼y�:�<��dJ�?�wJ��I\ҫ������K"jr�dz��(�+�zBc5
c� 9�ǝ�����(׃y��o�K>W]�IBy.�שʥJ���9e��Q�8)\��=#�0�]�1����Y���g�6`���W���נϯg�̟���N�
�Vg�d��������k�(+i�;�X��3;�bq�t�`��gi�+�d1�f��N
��1-Ȉ3��ZZh�R�P���A�@i{�p.
� � U�z1�I�\X�!u��WNLS V0䖙�*To5TZ}q���
��U����e��#��P*���4^��x�i�y%Wcr����˪�)Ѱ��	���|�:���_6���P(���ZT�30@o�7�������`bx��?��ԟ|�+�b�������Z�����܋�8D&ֳ!�q������h�ZϺZ�G7<����Z��P@y	��y��W��w� 8Y�pi�f����B��پ�Qͽ�>H��ʎ�jzU�<�|@͏F�?x>�vL��F����{c{BsO�(q��jb=x׃���� ��GY>��<���ݣ�~�V�_]��+�G� ��AC �666�~PZ(aT�&ݲ�rDHhq{��d��g=��f��d�k����e�b�:ދ���ېs�@+�2�����y�����㇤����S�*�(e�2���״K��ܽ��ܿ����=�`({R��Ƞ�nM�s���#�����Q%k^��%�2^A�5�16;���+tt�H�[/'��G��|ZR��¥`��t�'5ȲHj�A��Ń�ޡ��Ń�_����$Vyx�"�|�� �,�^7�W��Z����N����6�C��N�����]��] }@�G��4M�l�R����P��b�#P�'%u!���t��B�r�v 4P�I��BL==v�Ճ�Z8�r8RfT)$�{�x�����՚X�$æ�$?�Y�i#Y�z4YL�"�ᕞ���$�g	$�S�Hy�@�>ݿo��G�p;�O�{�ahZ�� <Ӹ�A��������#xv(�B&���`�y.�3�dP�y�9.�^k
R�E�X���/�O���4}΢���p���u�}��;Y�u�O�I���3dY�)��z��J;�����E[pʽ����܁�q۠ƖL���cF�$�o�d%��@�I������r�q�HI��B�� `|L;�� +�]&):�@!,�MG�4�3��A��y�{�C�h����Wrh``6�4�L.��LR��<���1��+'��M(za�/0��*�5��~ѵ��4P�9�9G�uJ�za�[J�t��I���>��@��S���W<*}.����� ��8uݙB٫%d:�P��Ua�Q���[<a׽g�&c���9���;@�'�}��R�V�gzq�)���a0AR&���j^�`���mP/UVX�f�I�WX�Rc��z䢟W>��r�m������y����m�D���2���[�k  ��IDATKT/ݮ�hno���N���a��D���֛1�e5�1+���G�[K�`[�o����4U�V�!�L;�{W�1����������*��{��E*oLo�AJ��{�]������)���i`��z�3��C�V����F�wu�B�D�kY ����j��yt@$��J�6���� ��s/�R @��f�d�ް��k���x�; ,~d��`�����Y���;�64
�`ؙ�54�)��#��(y	IK��!�;�������cؚ�����eRB&#Xp�'s�pǛOWr~�J^�y#o޽�Wk~���'d%���}��\��ڸN�\,�dAr��,o?�CW��LJv���{*�jȊT���z!����W�1ו��]%�=�C����[ �7[TT�/?��2?:����dFA7�Ho��֧���)��`���X����d�J���#�A8�#W�2pN�TF�{ �>��{\�׽C��&������ɉaGjn(��ݎ�K�WI�<O��,]�ѺZ��R�<���dp��gQ���g��� �-��ۻ+����eVO�����+)��^fr(��f�<���U���H<I2h�c�������|��~�~7����Bb\�i���'c-�Ke'���޵t_�'AW:�<�̩u��A\!�Z ���`}D�@��D����4��I�yu!5��f�V^�:fAb��@__H ��� �SQ< �h<��@�?A��XQ_�Z��/WY���9�����9n��w�	��W�,��V�iJ"� �Z*���z��8��7e�#=T;�>"�`f��X"BT՗����i-�9�i�����[�P4�Q��0��$�J$䆣������I�s;E�U3�9n���]��5��t�WIw:" �'B F���Ғ^Y������Ju�6bfxVU�0`[���!|�0�6*�m��<�a�d�zQ�P+�'
�L�iL����Q2�H���=�Ub�e�[�a���˦��k�/e��ɉ��6�*#'H>ڡB��M�p�S����)��˯.�.�|u������<ݦ�[�!~uL���U\�A�"�#2P[�*�%�\���r�z�c�:�l�A#7�Sk�4m��фL5}KĹ��@�Dq�3y7q�Xq�	���Q!f8G�n�7��[���:�4Ym��Z~�{�W��DFE$����j�����@���]W��zn0��7����
�s�F �U�ࡱi�%*T��;��պ�&{"ܫ��Y�$姹��� ��b[��h��~d 4b��;������eR�`̑ōm�],�ռ�[*r�`�:2�g��ݪ�ky��U}l��xK��q�PCT�;�0=ؘ{Ϯ-�p}��`� ٘�{Js ݡ���:�C�Ҩ���t��gJ�-�Ż�@�b�-՜��!��lmv�og��rk�G�#�l�2�,!���Л�,B�j<~owdXk:ô�@�I�Mj��7ov��� �������M�|ڑ�kE�a�Z!$n�f��P��P�a���+k�e��jŢ�8�a]!�"���lU�0��|��S.0<G���2e�8��^3aXq�t<t��?��FfHRFm������R�o&IA9���_%%�B�O������GV|tK=Q���e-��G���M׸M 9X����P&��G(.�ɘ!N��=P���%	�,�C�dYDC�p'���������2C��S'WI��%��t�}�d��w�dx��h$uB���ޅ,�F�]^���;Y�ρ�bn҇n�a�$�qt�1�ݧű�gg�w���w��$��Q��,n����dqw���yXc*�P�7�5����>�����7�-(פ%\��>��ټ������&�pF��5���!Zv�K��1Y���<�K���f��m�
�n����^]�f��wޞ��V�I^L�*3�y0�4&,LmEY���������I܍d���>�<�F�����u�&��@��3�y�$�r~>�����������WI~̵H��Q��S{R��(����D����,��6��܂Up��1gs���'F�J���T�؏���Ă���3�^ec��-	&��Q���W��w�����(�o?$�p��ւ��Gs5�@a��*�"�'0��������̪�7w�XГ?y���|��o�_}C��Ï�忏Z���mҵ�������8��i9̔`�gDt�m);j�D�<�8Ð��T�6���d6f��	�@۞��"��p�(��]A ���i`���z�j��e/ߔ2Y�{�ԲB4 g1�t���9�iM�#�uLr�I>�p-o�~h�S9>�y"iL���/�ne�F���'�����5$��k�FB������"�D�@?�f*�n�����c��鄀�kN"��u��Y#,����A>�$�{N=}(j�c�_З�L~}dO�zJ۸>,9���pV��G�SH�K��?�ES�^��_�v%�:u͝A`]�:��EZ�^9�2a<��IfP3�'�i�����	��7�*�=z�����t���u������{0���c�:,|JCl����
MÂ�Xb�U@�J!_h��'Ӓ�5���)���g�MWB�bn�5׬��DC�R-��_s����0t��!������ ���]?V����ߟ+����v5��1���*jo��[�c�C�Մ}'�g���7���n"��+�Y��$nU˥V7��uU���x�Uׯ������>�_����Q���u�%�×�����v{�Og��y������q����E�?���do`��������y�o�zo�V�z�V�u쿇�s����7+w��`�b5.�W
(���A�BP/S�B�J��T�ٚB�d�^s��s�k��E����u�h������j����BnPy}wG� &R]G� �P��Y���oZ�g` �z�ZJs�M�nߛ�JJ�rs�Z�'���i<�Yad��g?̧�Ӥ�"�%������-����j�LV�u]�Q(��Y��H�$����wfVVuW�|�3��}��/�����twY�~�N�������}��UL���  3SSQ��G��.C&�Ե�=�~CS�����ؕqb:%��F��7oа��.�)!��%lT׀I�������B���B�}?�+�������ۆ���!Ɛ]�I��������~ ި�C��~�Y,�AN�u����m]�n�(q���B�l=��qZ�od\ק�齠���ڊ�P�y����Z�Z�g{|~�ۇ���PqC�����Q����A0�UȂ��<b� t���T4=���^����QI4��?�&��eq�N����Wl|���?�zuΠ�3�k��,Ź>���K[w�bmFC�.�]e%Լ�c�yfC��-��!
��|�o���~�اϟ��Ǐv�U�=2��a�� ��wuy^ �+���r.X���ޞʽ�x��~`S��9 �N��;t@ۓ���X�w_���~�#;�=�o?��;��od����ҁ�+߁_W ��&f�HC�LYO�Ƃ��4M�L����ֹ��L�-X�qp���Jj���?[�l����LV@�)s�eP�L��z�8:�D`:8\c�Q������MS��gR��S�1܃�����?��O����iy}�Q�>//c�ȞJxIT^z%�j	z��Б�)&��38�2�7N��41�jK��E�#��+cVJ�*����is���ɘ<�C"=7fs�Vݝ�&����}N��69מ՚��#L����˞<�J!N�3cu՜.�t�Q����`NQ$���U��AE[Q��}*�4�p�q��_�݄p*ZJ���W���pXv��&@�E�w��c���Gl�������j�Xᴽ�z�夏N9�(f�,�1�������׎�k�-2?"^ϧ���&�� w>A�D=�}���;�tR��;��49��M�8������R �a��nk�r݃�KP��xt>��H���
�*��m��&���s���#�`O�j�@,� RA�{8�� ^>r+�H�2�׿�S.�P3a�ג��Ə�f�n�}�W��_Ԥ�<U4O��p�p��G���@�?�k�X�	>�^��(���I�h�x��j�@T�8S˖@Q��[�)�h���M�@JH���p���
0��7j�G�����n�#�,��)�]�>����H���3�lY$긖Х�i�U�XVfW,'�vRݤ9�W�B�tP�=h^h��m��Z����Ɋ]��E��d���(u��3TP�*�p�#�u"㔦p��T�>ٜ)83ͭ�8� ,WW�}��}�S���|bM��D0��cwj�39�jw���`��6�����G����F���[+vp5�P�{եl��ᡀ��o���>��I,J����hn��V��^�B�5=�Ɂ�Ư+f[/�
jP�<�dD�.pbc��]-�٫�oS ����>��h�gP�I�:)���.3��-RP��x�<�k��`S\��}�uW���i�Y'�W��:�K6�!��и�w�������?���}W���Y#x,@��g;87�u^���&�&I���˩��%��/#������`��?��9��F ��K���R����垬�5��j�$ծeFMT��b���'��!2f��=Z"����4��g�wۢ��]�����C��}������S�y���w����S�|ug��X�U���͙Y��[I��8�_؀=�k2a���`���V��]��'��Β���.0��,���H�Mڌ&�_�^�9�	�[f�Z(�%�	�F����DI��af ��_��?��&���3�Q�W���0�T��O;QCGm��F�����NG��%����S|�j�F`-b�}��t/m�}Z���`:����LY=JܻBnr:�b[���y��8
�F2Bo�,�!a߾e��a웕�/�Ws����p�������+�6$��o��¯n"�'�LZ����S�}'4Rz��-��;���9?{^L{�����! (!M���'Hu"���:��
ʩ��r@;:: �������Tk��*���<�"��j�8D]Ǭ�v~�{�������K։���+�z���w�;N|=v�	�U��_=��*S���?Ve�������oC
V�uX]C���ñ���HrR}Qf�^��Vl�ߊH��ݰ�<H��g�Y�n
����Vs�O+���U��
h��_����)�#0#/�~���1JS.NA	\oW?57�Z ��+�^�1>��V��-����Ͽx��L�+�[6�����8>��"[7��1Ò��eaѵ^o��٤ޣtR~J���Q=��ݦQ��g%�Π���W�Ĕ�6�<><�ͧ{�VT�����tuui�^����+"�>m5�ˍ��~�����Z���8zcQd���ڳ�F!A��� �ۺ�b�`|�8q"��N���5{����T��u�M��{�̠˦y��p6i�BѩmU�b�R[���L<d),R{8��2 �����..���}F���4Y�-uN��6M�Y�$<���w����=^d��5�:�4\�g<@5��^���"�Z& o6�ƾ٬)� ʽ���9e��1X��%|i@�"�-���0���������%�X蓴d��T��䬖V�>g;E�I�{�m�+Z����[�q��@�m�,w�,�iT�K��RY���5����6σ�;s��~ �Iw"!�N����A0�ʂ����®__�o��{����?����S�o�����0�ϋc{�L��:P5��L���k�jX�C?_I��Ye���Q�E�k�� ߅뭀$�Y]���[�;��ހ��������� _�Iy3,v~e�K�z�~���}#0���Usk��ݛW����,������/�������޽���W�p/��GR��	Df�g6h.�eݷ�S[4n��k����f����%ڰ������'��/�����B+��A]�օ� �V)[���g`��5��_��[?���1�{R��&��+�w�S6��u��_��V���|�T�}�z:�<�u}�e��^�I�ՙƛ
��O�\�5�#��b�����!s�;�ި�/�������=)]j?o,�����+�Ιu�ng���#�+{<g.}e����k3wE~��Շp0��5�w�Tg��#���Ҝ}�q=!��lVG@?�iU�O�Q�m�:��pL�,��}3W7����s�J'�ӗ���2N�\ܞh����	B��i�9s�&&P9�(�P��UMӽY1d����m��a��*$#gN�|Lr��x�o�́�hڝ~E'j�T�"��t�Z눾�\{����.��xq�- ��N�PQK5z�cLc� �g��oҢ�H&4Ef3�݁��)z-9}N/�	���X�9�S���b�x��%w�&�6E�}�g�k�p<x�!Q�����7�p�œ� ����N�h��Ѽ���<=��䀅q��<|�k'�an�r��ά������7�MtA;2rfV��1��O�W��M���`Fqgǜ��P��7�VΕl��R9�$z����@D��p�ksG��������Q=O����B(�|�����%�0]\\Pq������/X�L
�S���Y�*��8:��3�N�I�&ke�O|��u��x�����ϫE癶�-pK�Y���RX-�VN:���uw����[�}�QiF�"ٮf�tR�p>v���!	)a][�[��uSp����ӯ?�9'
����@�h���c̍c:�_Z����?��+�7��S ,a��P��.���ў���h�h�[�?n�jU�R�zQ�G:��
�s����]�:�����:UK��=���8�;�еy���ꚺ�t*hE�#�߳f��Ӗt�}9�g2�7����P��'����h��w��yJ���շ��=ؗ���h �0V{<�=M�/_,N���͖�Eq����v'd]�o~��~�O?���CD�X3�3u셷O8{(�
�����Oi�Ձ��@0&�������2��Q=3[���]-�}Df��}�%�/��K^��W1�^��v!5��j`��͍y.EHL��Gr;j&�L��nOWvq���`d�����ݾ؞�A��[p�F#^N�*�IBl��N,3�+�ɥ�����@��cp�]ʾ�����ß���/�\��o�ym�IC�fL�8e�3�d -�G�P+�JnP��tLd?��]��E���_��آ�
�3(��IeT��˦��{h�*�n v,y/�N{3Y���R�����r�T�D�����4�U�7�.^�7d�ջi���я��o��'�̻� IRano§�="ƣ&�j��OI�㲁#��oYC����ώ��׾�ο�����L��� ���P��N�4~,�^AeY�����.��H�ٜ�ZQ_ܴ�9(���&����& �(Y/�O88��,��	���!�a��b�)����U��͑t�7I���)(�4�2Y�5�u��&K��d�?f�aAK�	<w���^��w����WSp��JGT�ʝ��bm8��j�Z֤EEm���~"!��(Z8X�q0_����6������4Q��	9�TS��GӒ��;n"D"y���*�Lv�]�d~ς�79j`���;Ω��<�Y~r����y������,��Uv`��Y`�ͷ�o���{�:�^�.�c�yz��S��N�L]���o�%p��˸�����K�T�)'��S~z�h!"r�b~|�!̡v��B� "���6�(B&�J��r0:�E,˷�q�R�߬k�BP���Z5 
,�>�,��"�=�sq�PbC7E$��kE�l� {�q�N2�봕Z��V���#�� �ŬT�Dg`�Q}���,�r��U��p[��{�L����ʃ=o�˧_�� (�oD�J�Zφ���G?^>b��O��������|���F�r��{���ϟ���!��hT��Pf�#�t�ۨc2�ց������Ε˱+P"�W֎�Y�(#��ۓABZ���t�L����R��  -�<��!}������� �;��9�g��V�d/@�귭=l�������Kfl�~tA�5;�M�z1���3�rz��7o��ݻ����9U����ԫ���h�����dl���Ȟ��;;o	Za�P������������� U��-WQ\��q�1������\�L�*z9���w}�ʸP�� ��@%��� d�W[��B����	tυ����c����QŴ�SP,E@[5p���*6<��g���~R夗����
5[����Od��޽��7o���;)����j�����5�����_�6��X��S5�kB�A~\ro���C�w���A#?�s�n4I�x�R&Tle�����3�o�~dT��k}���@t>�;��;���A����7
ʵ�)����iL���̛U�W�+�%s�6�<���:�y�+���& b~�4v߲��N��6ޓ�����U���J�N�89��$*;l���Ű�K��u�7E���[��I�^�F*��^eEo�����̢�=�ᨆ��:��8��u�JǇ\��p�:gW@K�ӹ	��Y��AE�4�"�R�q^/7�4;�u�D�C��u ��G����hi�sN�k�Q�1������7�ۏ�D�_P�,U�|2�he�%���2:��9���H�P�c$��}V�@W���g_���>$�g4)��"P�*p|:���V��"'* ��&� )���D����t:�u-��{gw6����]2����X��i�GN����h�)�7 ���+{S�/[u��d�z͟�:���ɣͷ�\���t�~pś�H�5Oy�u���wў >;�Idx�&()�9ac]�
��E-{�u��gF��~���DM��yM ����Ơ"y���gg'�	��Z�bD��Y�����͟�
�]�O ����ҳ4��TC���jF�з5�k$q��u�2�DOs��6/1���'Hy�|�d�y���~�Z7�+y�#F��n��������	�F�:��MJ�ؗ�������)$���vV���=�P�F�Lӷ���gN��{�xñ���KJ�b����N�.�ў�>��-��/��F"k0�!%Յ��!%M���LO4�Om��Y�;n"Z�&&�L*�&)�`8ǞY!�Yʎ,�4�+2ɐ�mH�ڣ�H���<m5�ȌKN��,T�z��iq���hI����+!7�k`�vPC�,������c�
�������zO�}��ۧ��~z������@ۏ{��</`�}eo	D@��t���X��]R=�P4��|����G�=c/n\`AY5�J*N�gm��>�ZAPtT4����\�A��b�N��]^\��!B�d�BUت`��ic7�>�����=d����ř]^�r~�{ ���mQd��#<mY�E�>��QC�ƃ�S.K'2z`ˁ>����� �Y.������]��|�_>~��b���:�P��䬵��+�~����U�/mS�
�$�%�ٲ㩜��ԅ6�%��������;rH�Ǣ�����M�GP�J��ehى򴱳~m�T^���G��ܺ� ��������m{r#Zy�e����H���3P�[�+��( t_���-�?��f�8&�H�j��?j��s2�a#��r�y�w:3hf�[<�~�ַ=�)����?3m�I����u.�o�?B����v�����-�eȟU$�o�n�,�M���a��	��b;Q�́֜>h�V]�I��ս�^{��4]^��������O�K�g&��i �9q�Ù����V���pƦ���ʳ!ٝ���������̢e�ˁ��[�/"|Y?�1��t���c���a�NQE�rj��jTX�Á=Ib=(��,�����j��(���~��Xk��0d��x��u�h��dP�<��p)oT c�
Y�n�oYG:`���R�`�: �-���g
�Sv*;����G�1Svz�Z�:�3p6���L�9\�\�oN3���#�r�ѹ�|��g�xv��Y���3�ߙ�����w���߇ɮ���HP��;��@�b�E�@R���>��:�̉��+��E>�����'���k{����z}M����O��_~�Ct��U� Y(�n�[�L�nF;FD�%D��v{��I�uy.&���yoTa����u8���m�D=5O�]�ydr�h����vLs��xt7@��t>�/�s��uf�OP��i�����`׀>�>�9iY3�>\�)�u',H7�Օ1��S��#�U�}��x��{��B&�m7wl��p�ޢS�Gd��;��Gѣ"5T;k�I�# ^�Jg�爂P&���@5.����A�吘"j�'29]#�
s�2�A�P�cny�c0]��M��߬'i%L y���k<>����6{RrG��:����uaN񵺖(�=x�����Ԡ޶+���?۟��G�o޽e��u=?l��1P�=
�_��FuMwwvsS����Pv�4��ʦ��Y��ʌ�zƚI���E�?��{5 ��d����Յ]]�S]����c�<b[�ߵ�	 `��/����}�����z����ia;pO.�qу������I}4��MO�P�w¾y�)G0 <������2��ō�5�&��ʣ��q{ԑH*�-[��b�}9��I�PyY�Y����^o��6J���i�Ĉ�r��f}���je��O��!�U��i�F�j�ٕ���y�f��2s�$�SmtP�,�){�Խ&�z�ki��+��5M���e"����vu�yqR��Xl�g>�����(X9�O��K)��b��L��K�R}O�a�#�s��#��K��$��_Ǟ������kKq*�����9�?z��$�����l�τJp�=��U��kMc�Mj�ǛiDy�iGhr���D9�輜���gɉA�;��1�����륒�R��b&ɺs#����1Wh�?ŠL��}�Q'��K\�R8gyr_z��0��@+���ߎ����왍�;�5}i��f�ZռM�����O��e�F�!"���R�l�?��v/Hq�]5 �@���9GZ�*j��+�%ZU�)���υ�A0�Ni�'�dU-��]P=����N�p<3�f@���hu����������&���3t9W aѴ��OT�	v�3$��� s_:�����>�Y"٫��Ǿ2���}��pF�'����L(�^��g�7���Ϣ���V�.Dv���e~�R����Li3ïQA[esϼ��"-�l>h���ۻ��/@�l��g������� �	J��ޏ�"�f��ŕ�Ҳ����ʶ=5;+(h8��9H�+*�<�0�2�VNXO!���C]��`��[\�ͷR�L����@��m>4���܎2�k��b�ECbf�Y��f��-���!˲��eqJMMW�(�g@���Ƽ1��gzL����xƻ��v��-�	���d})������^z)m�&ӽ�uN�M�1�=5b�aES���)��h	�U������FA�#e�_�)#��Z/����*�}�H4̢j���ڏ��ނu�����)k��~k��bz����nl�,�Ǫ�P�-��kGR���Y�"�]dް/��3���������@A),�^ŖK�g/�=�"keR�Dj���%���
�L� �LwrvN�F�1�2U@4g����+yp�`� ���ر�+{��`� �����<k+���1?:�{����ͯ��O7����l!��՛�����J��)��Wx��7߳5����l2���=�Y_#�t�c?`}KY��H�24�ٷ�a���^�s��JȾf���f����N���͵}��=�V�U'c
��Act���2����k�J&&gG#(�i&�����`�j��{��ڮ$��:.S�I	��N�H�s����)�9�$�����U7c�5�I`�R�
٢J�n��!�� �E����*����޽{g������˞�K���j���'��T@�����<�)`{輌@�����Xs�4�w���տ��z���ܰ����-t=���n����?�8P:>f�0AT!�mU���ZbA˗1t��a=���@���+���!��~DS�o �
X���8��ajP�<ˡT[�,
��D�fb�٠d����U�A5��c�2�(��iӚ�Nw
�魎�Z�&�W��o<��&�ɏ��s�(��[�g<lrn�K<���iG-� #��K��9�Bg���~�Q�A�a�lְ�B�����	z�j��Uw3Q
�#`��Mm��
@��TF�PE�44Pj$O��a�!Z��_�����c٤P��c/��f��C9$7;~Bʆ藠��޺��e�8K㑼�o�~E#kl8�g�x����N�6L�}>g�`G ���c��	@��Z�F�85E�&05��~��.�(�P�?��}}��Ѧ��!����R�kz�t�S��+��uAʲ����1��1ќtL�J�撵�Ka#�����l:W���{{��-i6p"P/�l���#����fJ���^,�H�2�޴�]7AF՟�������a(�{khs�<[̀.7���Vr*��+���;�^790���N���ܬ��^�Q��x��REN|��P�#�� ő�גxM��3�y��MyF�xY��ՙ���Xwbw��F8����i�}�o>�{Ac���/և;�\�L�����>@@ ��}��Ѿ|�X�ϔoG����.��vR�pE�� ��q6u/���:�0jB"�j^�lV��a����U������	�����5�s�J:RF`-O��X;��o�l� s�T@��S�T��ۤ���` $Շn���f��q*�I!���k�(=�'[#,������g�姟��#�#!�����?����Q�(��Ԗ�\v���E�#)���=2xD��1 Yp�˱!���7&����b X� Y ��Z��9����ͧ�uЋv't{���;�pM��x2[hl{[~�&�S�U->�w߽���3��7�0R�a�(�g��bC_���X�;�h�(�[����^5 �8�k� ��(�* �2P;�/�.]�����X&���?ؿ��?�����eôA�o�]2�s[��`tt�����1Z��-�9�7 }&a4� �r�w h�_�ER�r?P�38s��r��]�V��$��u�'�-j��c���l�9ja�4�d��z��Ţ�_��|HJq��w�F�W?�����������/�~���_��>c�?QhNmhrMz�)� �qeD�88�~RMdپ	��x�����+�g��#�0�_�I��O��+�g1�A�7����YA�	�4�ޡw\Y/�
+�F� -��[:��e�j[�?�XP$���qb�yA�7w�cDG�N53L���m�zʇ��;���9P�E��	���(�+�=�U	�L���N�'t`z�>�.{%�(���/Gd7���A1b�ҽ���,��Z1�b�c�c]�j�н�tlD���>_���s����I�|ǔ�G�]��9$�O/��g��v䜫	Y�F;��{'_�Uq���B���[�� U������|"6d�-�KR8�&��H������&�=��t�oNL��2�-��5�Q�$�pu��A؈&��z�����P�Zx��k�+60��Ɏ�����V�'���T�p��zF��gQ��biJM��ńF0 �+�b��$FL��q�76/R�(�K�E�pTwt:PD�"H����z��"�\���H�0���
@6�,f�b�J�ˇs=E�=3+<�dvG�C.1=g?v#ʆ5N��:	�݇A;����|���{��{	;�R�,�LrFGϸ�t]�"KJ��zVH��P�Z����:{k��KJ1o�����)�F6�lTK��y/�c��)b����9x��Q���eY{�`����l�,m4�<��@��U����T����Ӕk]df���j_P@��ي��qw01N+�w���y����G���w�;U8o��r�u ��:R�vtA��u�{:�jv�O�{Q<��9t'�<NyN�2�{;�|[�ʒk�v����=3�����:VIgDYM��PU��_�
�ܸ��<���U�l�~�9��Ծ��_Rq�.�V��#d��1+��ȶ.�C(dn�� (hǘ>���8��vw�kX.N�/ű�����w>�q\�FLL�Υ�;�<0��A-��
��4�<_���WM;���O��ѕ���9*Sܔצg�R�d�aP�5�lz�-AݪY�|k}Q�*j5a7�8���y�P�O�b�˝}�C[�3�=��s)�+ ��=�~ ���@*a���RȂ��:�8�}�Ý�O[K�����r�޶϶�lH�ܗ��8~���3^_
Ё8h�����8�-�V��Q���Ȇ� �P�vT[��4gHG��u��64�ʂ��:�ɳ1涎-s`ò�	�!؂���e�M�Y��f���P��q>=r��z���opj���*��ߍ��z�����^]�U@��[;�s9=Kemc��)8�u?.[�/6�	A^�l`n�{iN�Vvvv���A5g}9���b,�]�����~g�����
���l����V���/v����������%�n�T+�^\�.s�}W1��F���3��N+��	�Ц#kz~��z�q��$s��S>�a�-6nSƯ�8[�s�S�V+�[�D�|>�q��ðs���U��m �^^q�q��g�����w�/ֺx���Qg�����×2g�/���
��Z-Z�y��������~�[�>�h�+;0|wsc�7��<Є{j��(��.Y�!�u��K�F�m 1ȢV)��"�����t#��L��ݝ��7�����L`��Ԫ��X��k=w���J���Yqo��d[���m�O�ٔ9D���<.�I3��G��9��H��BM�kcq�����?JHq ��=Atc�f��){�h.ڥ���3J�[��S������k�~m~���i���9F')�7���T��Xu�c�gD��q'sd�I���U�n�!r�6���7��%�:�R;w$��դ����*QC��F� ���FFd|�:U����|c9�{͈G����ѮMT-0�6r�̵ ��C�0�8׌�@W�"̔%��Tub�M����#}h��e���gW�)�MnmR�D��D|č�U�%6���G)/�T��ī~�����u���Q���?���������G� ��d�'�ڬ�؎@������U����?�霢_G����מ"z�N�'PE�;+��c� �i����ݱ6�FkA4ՐB^2�C�����f�s�'��%mג_�<`��%j���+��!���]Tbt�bhY�I���4���2��J����� N��}H������ߩlT��1���.D�m�G�ׁ@�8�a�AZ�S��~�2����#�$�[a�s	}|߁@�1��Y8KpD �P������|7���r��Ĉ�Kh��S7�lHe��4/� �e[�M߯���l1����4����G�A9y�i-���$jk�q����&M`YAD�n!(���|aC�(�gԜ�E�Æ�W��e�,5��#If� �랷*�F}�j�$V��K�J�k'���v���ʙ�u�I�!YP	H����u�Ae��:8�T��Xk�Rgpe7���<��� Md�;��:�V��
k�3��i�.A ˃tC���=kdD�]tq�&<���$�7[���jh��#��P
Ь�X�/VU A=K�e]��4e�j�>Dك9�TH��y���|�%��k���ƴH�/���5���rq(kw_���Vj�YCy�l��x��_��,"x��2j��5����"�V�Q6g_���	�9z�uw-i�tv�AF�8��a#�@3��*�h�������s���y0o�}||��甠����K�V�����{W-f;�욖����m�3X�`j��<@!�
6c�^��b!�S %T*Ѥ{�j��J�Jh�<@�=�Y�S�m5�$��e��P�&���Y� xzjCϘӃ�(�٩17��9) �����w?ػ����=�w�^����MPŭ����5�pr5�ٝ�I�8��yXs?:0G��w��ER"XG5�U0#P�D�ԛ�����g�S����,x�Z���I���#��d}ؤ;�Ŧ=������ �Y)W�V��p2�̀�! @��s�(�j]&�	�N���6B"J㙬�5�!.k�d�Lyv�/ 7�٥�)0�ձ�$��_4ל��TU���{�1��91m��:�ܐ*`�&�����|�J���r-�g�{����[�?�{�P��X�"�����#�x�@�kܨ-���jX��F�2�;Eɂ�Z#����֢�qV�Á!ML򦅘�ThCDv�){�BV��r����qe]y�+�k���uDi|vIY���ѻP�So�aE~��^W��c�]%��)\2�����l6�u���0�:ũ�0�@DE#s~��k'2�Ӝ�y>���Jߞ�/��o=�)[sZW��0��
�<�G��J%���i?ѯit�������P͢��YRTX�
:se3���S�uP�6�u��Y�%��쇑�ӛt�g޶�co��jw�PmW���L�С����L�U1d�[�x�Gk�M�<>�`t�:��[�4��$y�Z7�`�k�q:R�U-��Ha�ܜvr��Zem�V>A��hѧ���e#�<ޱ>e��h��A�|^�ӭO���`��#vs�=���sk�*�fP��~c����i�O{E=��s��<V&�
��8�I��f������~���7�tkw�?�uC�=�W웖4.�����
j|z��"b�����6����W��Z�� �v{� ��=�<Ξ���}����'��$�r�XW�Fs]��CD��f���4����<�@�n[��2�@�CO�A�k�^nZ+̈�$�r6Eu�ߞt���Zxq͠��r���j� 2hE*��$6�ခn���5SgM,������;D�e�Pہ=Υ�c2S���4f-�3)F�E��hX�>K��Ŵ��ř$�Q� u�lhҬAY5��=��2���h*��C�ab� #�f��q���N![I�q7Љ�ga�A��.�����2����G{�j%�pݺ ������y�FvK�t����w�`A�R
$��� #iӸ^$�����"������
T�ڧ\�BF���0���9�i�=�
 *�C��Y" T;aP[�s0בA�.K���t@Ei�p�2��]PQs��M����R��:!3�;r�������]��`o>�`��y*@k|z,s�yf覒mFQ��fa�f^����7O�	CW�e���8����3�~
qV{y���ޚèV��Vx8�DK(���^��Rd -���=���u�����ig��'�k�&'��m[��i���k�U�$R}ɯ�qcƈ�rI'i���SS�Pj��M+icD[�iw��1����ɜ��ɽ�9��.�M1�q���&L���I�o��ș}��@W���Mr�"+�4��"��@�NG���=0�pl� �v,�ǭ~�
��
��O�'�vC�D��f����`N��t^����JQj�t5;��F��n[� R��?p��-}nOh���N�Q��M�BM!��F�I;6vl!�!�5'a
/����9at��&}��6���(5<�׍^�=O�hn�|NcK�H{C\�u\��|��9��1�룉�F�1����S3�y�d�kl��8��y�ά�4)�Mʳ9��}�E�����e�J�Ԏ1 )֍߷�]������><�°3�2f���8)���rF_7mmg�`<pL�$ٳ��� Ǳ�)�u]��ձpeT|I�m ҍS�g����48dO�
䝓D0��q��6(@�=p|ػA
]T(Ħ�N��Y:��WH���7��~+�ÒE����J�#�c��~b!*R�v��cC�:��D�<���������6ٚ� ��z4�ڐ:Cbc(�����d���Q���i7�'
c��jh���H�i}3�ۏ�k��j���ʘg��dڻ���Ё�t�9sz`x&{�@2X��@ﹱ���b=`���\��.��..�'�j����'	A��oT�M��%�!��RH�#;��|�u��d��*�d��lź0)�QԢW��4#�-���)�����*�6�x�j�� N-�:��n�̣���>t���3g2h�'�b�5�o��{�$x�����i����	)m �b�e�E!� Uܦ���b�2(l�`L�!k�c��,c��a`�t��Q=���"�@�I�s�g�vS���L��1�}���Sv<Ӷ�<�� ����իW��(��#�v#�0���.L-�<[���m�w���@���R���e�Oh��ӔY5}���S�<��v;��'�c<�^���Z����cdl�A2��H�E����ͽAUf)F+߄�	��|�k�_R�L���$[�0s��/�1�!B挊䙩&��u�����d{�}����Vo��2�Fm�.�d+�l���n�A�D ���gH��J\.��v^��UZ�7l}�@5l�6��M�wr쇪9�UR�s�4��>E���������9���p0VW
`������<��Ef�c� j�Sd�Q��<-7d����E`�V�u,���`-�|�M���G����ؔ��|���E�*όRuL�nT���tCc�iBµ�:GӁu0lJ�3��>W���gە�?�+FͲ�F}�V���֣y�0��C��7��V-�,�y����y4�K<�y�?C=�H����EV+�S�$BZ �*;={d���}{*�F���֡lƻ�9�D)Pס&�]�&��Ftk_r���DQ)�,�s��MŸ�Vʑ,��)�-��旌�Y� �U$C����^s�)	8N"}���	�%�k� Y��=y����8t�hi�Ȫ�x�"�H΁��l~q�c�����^_k���q@�.�fIY�)33�`N�-D7�h���ϝ��s��2��f���k��q����8���q��,O7����rC�.y4=�^�y�p�a�̊$�ϣ;c0��v�c�>�W_�`�/��l�w��lEFG�۱�ɝ7^ܟ����.6�V�Mv����U
�
�s��{��û�3d�V����|�b����>[��^��6K���{���}Z��q[��6�<�JJ�JL�M3�G���uWƺ+T,48h���~��:�Y��%���K"�;��A6ܔg�����!��_[9����u��x8A g���/�T���"9�2us�YpTS5�S/�G(�G�zE���7e����~�������W'ꕋl|/*v�ysg�����������S�7�a��G�����v~qeWo?���+e�@-ŎhÉoM=͖:�r.m�v�N�8N������V����[���,1�q�:�ǆc޹�%���y]�� �p�H�N�7��s�
p�s'�=��&i;弞˞���`���}�0�j��虫S�[�)�F*�fǱf�5&A��S������ Ⱥ�����+6&U�Gb3A5��s�kE*ނY,�f���E�sG�!��sos��B':
��62��V1�L��4F@����W���}���0��-X�qqqɦ�������H�QB@��%�hg�Q�~�\��
��~<1I�7tL1fk*
 �:���z��-�O�>��h��t�${��0mt��a]�%�v�*�[� ��b0z'��6�U>1�X+�uӲ�׍�������`5A�����:���;��z9��㸰l|�~��IP�l�5��u�9ܒ���S��2�Xwɢ�������脬깝]����7��<���\	\6���QcӞ�kjR�N-�����8���FP*���o
�LB{�J�5ߥ
h��㾒�xG�+c��/QQ-FFqfcY�je5�5
Ta_c=��C�^�p�=Q#��N ���2�t����զ��ɋ����z�o9u*�� JHa8棚����:�#B���f�~��DU�@��;��ݳ&K�8ƹԄ[
�׌���5�ӂ\j�y롵���b��I��4�w�����fܱ[E�s���f8��}1)���g$9g_����	X���� ���I �׳�7\��p��<������5%Qѫ� ��������j�ȅ:N�q�@Nw��h�����&���Sa)�B�^N~��$�$j�P�`9�F&����� � @V�Bz �r/��&I{��M)"�j�Q���ik�Σj�Y�o�7O��@y
�n���*��y�e�䴙�+�1�'���W�b�`�dT,��W���J/ڨgmG�\�@�{p�ѯy��T��3�5�����
6[(+�Y"6M�Dy�ܴx�4�`���>h�"��^/�(�"|A���,��H)�;�%P�R���HՃʆ�� Ri�Ж��	��A�hD�A�>�A��7��
�#˹Cm�+ o'P�D:+xOW�c���s�!�Q⸃���oÿ�݊J(����TC�r�I��m�� �A�������5c\��8Th��=pJY@z�@'u8d��J ��J�{Ee_�}~��ϙT4	 0Ԍ[[]�P�㲜��T���g �=$�f�5��,ZG�'�&��xT
�>?��_/���U��6˲U1� �aO���k0�p��` �{�>c�n~�ϟ?����b��~�D�Cuz��s�z��._�-�w�Q����k[���&�PfEs-{�kL����xǹ1 ��A�)̂������T�<�%���]_��l�a�F i���Z<F�Qˀw�B��nʶ"��:_\YNYfe����M�!�X��۲��=���y�R'zcE�+彜"ƀ.2H
"rfX��9���I��k`�z݁׀ϣ���r�!��57�	Y�F�B�[���;�ô�8[��⣤ؑ��Z�(ID%��r�ܤip��ڶ��fW��v_���U�@=��1�IJ}�s���B�,砤�3U7�'���戞��҆ʋ��>�x�1�� d�A��`�ꠞW�a���э�N�iX��=�Ⱦ<{��ۭ�Pb�<AU@n��B��dQ���ш2��u���LZ�t@��te�>Ė:~P^nİ�=]�E�U��g�jH݁�f	И�|���a��\.$jB�6H�� ?�fk>@o��jN�C։c�^b��w���ֲ�{�yH�vs��� E��A��lc���j���f����������i�u���+��~k�O���T���pM�6��G�H�^^���71�&󩲐4������T��y�C���QI����ɧ	p���&�E8�q�-v1�r�}��ZB�U��'��u�g��B�d��&T�ڊ9�͂_��}���_q��V��3;������E��8Tqv�� }�w����v��^O�h�^Gt�1�	p�Vؠ�hD7@�c㲠*NN�
�S�^=Br��b��������3:[s9�I�vڊ����9�ܔs�$'cD�S�
�t���R��X�i����n�A����~ ��-#"űB������޽}��t'hA9�ey���N -���ZQ'J �{�L���D��=��kM4�Ӽ����|1����Hg���j�15�sG(?�}f6*tc��EO~3��Pו�Y�|��<�c��i|��1&��|.qÚh6u�_9yd�Tl�~}����B��.�Ms6y ��;B�T-��8��/�W���0�CU���^_5T�8���@�w�^Ӌ �%�4M���m��l�\s!�~��_�[I���*�Gʵ��@�A瓏�*�c�x�A�$��O���mZׯ��& TZF�W�_�f�M�LꎞEԋK�$3��y�>^��Műؘx���ݏ�x�>r��� ����|j���"(Qٕ0�ȷ�	t����� ���+�c�\��g�>/�97��I٨�����Yo�=ڏ�P� f���2�OOO*���b����S��Tp�]�����*���z(��8ǧ�ה��P���W��F��S�i��>��2����8���6���4� Z1W#R��$�� ����ԓ�oQ�P�9 �헏v��_���l�>}���O��S�c �8����w?�ή�|g�\��Y�0�%P���, ���>�0-���� ita�,��)���∴�R���� -�@B~��`��v�3A�zѲ����,���C�� ��u���3�����Û�k���gvC����>?<ۗ���Q'Ѳk߫0zp�I�j������f�XH�3@�
�&� �s4����{ 2���1`{��Pқ��L)��5n߼�M��h��'�������@Q��}KW]��X�׽^LL��8-�QC\զ��(Z�α%P�
�Q�̒&���j�H�M@P{�h΁v鴀	�����I����
�^Ӿ��������/�J���7
%:�Fg���i٫Q��8��b(�@~??��� �� `��|���~����}�"5�d4C^���� �S;�@��9�0G0"�xI�C��۱\�U�Mf�uY;�0�;P=O�-���2�S�"|���=Q�����D.�����ژs��҃�]^��C�A(��:՚],BQ4������Z�f ����]�y�@ ��d�<��������|�����~k�߼*s����� u��\���5�3�H Y=7ց>��}kΨ���)#��Q4�y��W�_%?V~���60�6�`�-N
bc����K�B�<X��/�X�U�QoVR�P��x������貵�T�D'mw�#8Y�7��.�fQ��k�6�9`ŮxN��.7��J�;wC��md�Qt���~D٦�zU@��0����nO�|����Bd�R=�T�%���~i2����qIc=㳞Ur�/zfE!�6�\��ɿ'���s;����g�h݀m�eY�K�Dxr4Sv����V�k�z+�H���������Ö�	�0�������޽����}�恐]H��` �V����
tY�
��r ����.�u���� ePM��T����N��B�	��s�q8��Y��X�ߊ2p�Gv[g�J\�h�xA���;�6O�W',M5@�?���	��PL�����h�i%a���L�*�D��W�q��LTw��M��et��h���7̱�_�j��}�<�g�lcvL���G�B�QF.۔�"�Я�k��ee�Ɛ7��8�+伓�Cn�u��\��}���>�l�޿��Wt��?C?��4a�u����A�h�iU��W����Z�r��g4R�e��z-� ٣����V��VJ%�Yl(�<%���{�풦8I�?�w���ƌ��U�� V���O.��^���5�y@5kN�MXvt<�Tv�^�B6"�+v����}���N��\���-)uW��$�`�-;�����������U9�WšQD�y#�b�W��2��j!Md��<��j9���T�D }u�5;�W���1���n��nY��� �Z��B�{�P�˧����?��_��g��� �EGj������</��[��0�c)��o'Z�|#�j�h�~���*��F��0�z@�\��
[����C��Mq��e~�t��nQ�WST�ե��C�){�A�l�K�':�*H�R�� �ǲf�6d�9��64��9�O:?��	����WUA�"��UyB�7�k�.//�\��x}�����OT���<c}�g(]���N|�7H�g�J�O�+�Nዖ�C�g�{=�@U+uD�[#�yT�hjn��0{����I�K<�硵�?� ��E��V���1˿XЀ�5xP������͵u�d�ݢ��M��������z6	��e�G�m��c0�2���@d#ň2��A��x�w���;������?�)���v
���l�P1|_��?��oi8�<����h`ݹ����FX���pF1�,3�%T�쁺,ju����h��sE�j��l0���p h���2s�@�-  �æ��깖����n�%kuq��1>\�ggTD��PĚ���:�?��H䔾�Ð�S@�o��`߽M��Y��=6�1�(jP�E��8�y�(c���Н��l)�2 Y^Zb����������Z�'��~�}�f���t��ņ��ti����/H�;��	�C��q�K�}j�Nm%�p��]W�+þ�ܣtJ ��Z�U�hJ9�t%w�����i��e�X�����(�ّ
(���#N��B���bJ��l��*R�R�u`�~�{*2�=z6� �SiFI O`�d�(6Q�Q�l��dl�3�6�p����,��:9���/��\u��N�	$�Lc��^W�^�vw�����m��qG~�y�%���E�8޽�`?��G���wvyuQbH�f[��z�[q�Y2B�S�jM��ʵ)�s`4��4��:���z-�g,
o1���}�/g�����+ӥz�������u�9��-���ëk� ?܇կ�zw��31�{I)毃+OeO�����c}T�a 1�J��� ps�'�;��������2�>�-��M�%��5^�7Q�׏Ƞ��;���1Q�U�Zŕ���
�浠��P��F��g�Z3���Suo�4?��B{�� �>�b_��Ɵ�N��������󲑯x\F�R㍍5��\�i�Z�Le�&���ʳ�"I�6n?��zϨ6z���ѷ����z_�2[�v�� Z)�q�#S��B4����J^{��v`�9�փ�P���,���溼~Q6�S�'����,�%a,(����4����T���Xo?��rO������a �=5��6�������
�a�:ҫW;9�m]Ωa�8ز�'�R̷,�9exD��Q)X1�g����i}������ȣM�].=��]<D8sW����)�����/&M�W�-�S���^]]�������[{��W��-v�x��Xp*)����@�2�q�ju�ù�B^ڋCl��*i��B���\��,�y��\�RN�'l8�E����x��xɃˏK]��G�a8�O��}��/��}׫�J�2 �3�EF��Պ�wL�
����N�-�= �������kʐc�D)Cq� F���q�55zm��*fBp�;ͥ�='3�q h ���n��G���`M���p!q �!H3Wn��f���N���V3ֽ4��]�D��]B�34HoT���b�Q�s��Z�-��D����1U ���iS��D� �b&e��H�u����h)���5�/e�Z�Ι���l[Cߠ�q9�O�>��o�b?~wn�ם�~u�O�������>��8]�51�$	���r���Ov��^5�!ZQ�U>�ޝ������u��h�p/r�9P@��ၾ�Qˑ�<�t�R���J��fc77��� $�+������ڕ��aߵ�i4�@1���A34Z�t�Ѿ|���Í�F��p�U��yzv�� �w8>��U�������:�J�,d��w�-Ѷ��d�Wʸ;�w����w�{��)��&^R
��]s����3L���?yf.��f� u�/&B�JF(&�"��`"��=�YS�� e��F�:�b��ռ�!S�+Տ٩�����X�#Em"Ǳ�z}S��/��ɪ��ށ�QϾFJo�s5R���xAk��o�/ޟzE���h�\D���W��� YS;�A[ج t�2�.�`yJ1�]��{�we�K�8���^�P��lÞ\�(ҎOϼ�#�8T�R�V\nc���_m�{ ���d���1��J�~�lXb����9�����c�	Dl$��[S���)/���h�ݞ�l��ҙ����c�#
F�kW���'�f�2\�QLuE�����Ȣ/K�ҏ�T�q�l�
,W��g�#�*!@��c1r]9n�W}/4��\�c.���%!E�kf��B��y��XDv̹_u~T#�s�"��s0�{Y�3b��@~�ߘwp�8�:���5?�:q�f_|I��B\��1���¬8N���̓V3��������B���N%��'�>�@��@hZ9�h@i٩=�=�����|"ا��jZ���ʴ2����
�7�^�E�U�܋��#�]�C��ܩ[<#�I=�@CD��MC�bY����-�� 赭S����3�'�@�e��5�5�r^@���^�/��^��,6$6^V<͢�u��8���7�)�����>�������v������m�Ɔ�N]�<Q�XۡikY��r�m��y����2.�(̂2�]@�:��9fW�l�@>�+8��Ӽ�#Ğ8�0��l5�hM��4������&��KE덁��G���/�ϟ-��a�E`/�2G�.������������o���3C�80�O�XEդDPJ���K�=
(�1߅F�f٢X�H,�iM�Hgx��P1\�gC��]Yg��(�P����ҹ����(�>�j�D�Qg*,Wp"�6�������̘W��]��ƃ����.@	���A���b=��b�N�`��g�tޱ?*��L`u_液9O���Y^h� �ދ���zz;���O�'e�.�ӻb��p�5Q�R��xM�곌F6��<��o��M@r�/0�$�w����X���@I罥E����c��ȟ��H��E?0�ϛr���X K
9x]&�A=4;N9�����
4���j�k�^:�Q����K6e�%�`%���Ӣ��å���ޗ����	p0���[ҽ����< ����y��������K{|��b���NX����Q�uqqƞU��$� AY�,>�����a��N9�g��y�N!�$��Ͽ�jw?[�y.6���o_����] U�k	4��
�O���tsc��zew_�p����](���P���e��o�Ӯ���I������Eʾv�<(���U����6�x_��`e�4���v7(�V�-ΝL�܃�~X�g[��'�=��ό=_����E�f�@d���Hu��Ŷ�Q��t�֕�����*J�}�\�M�6��J�կ��D����旣��{G�R�b]J�0H�vj0��4�)��;���V�,�'�aL¶�;����l(e�BE�T��:*��Z���D?��F�WlbqnlU*u,�E�S)��}
z�~�����.^H�><�Gj�|����	G*��a���N3MNE|ew�*��u1���R���yB切��@4����Q���[F�X��+sE�o�N���so1�8?�W�W������(]]	d��C�FQ4��	G��B�����-N��/O�,cW,j� ı % ���=ت���^#�褚�9�^\l(<%��S~�M)-�l3�HX�E���?=������ئ���yB��ͧTR-V��1����4K�����i_�C�Σ�f�k��Qw��j3�Qg�u驆�� �^�>�:�{eW\̢ύ.����s�Jg�8e�"|Yh3�R�����2u�����s2jNXX�cr]��Q�^�;�"�⶙G4��H���4�c��=7�޶Ł@=��$�0A�h�aⵎ��R��=SRz��336��F��DDv���\�m�v��=��w_�kS�/�{ ,j&LΝ;2��,3���{�����[W�35��$qX�_�cS �b-J^Cb�d��l��u#��d���Zr��Gv͒�R��b�C�+�ɾ�+����|��G{�݇�`������O�'����@� ����yk.A3��J���O ��%h�?��������O����?������2���d�:O���l���:������2�=
���񸵫�{{x�hW��۫�<+T��"�7i���h�Np.1{]�y�j���ڄ�$&�
��\ �jD���U#is0�]DG��:&/L�*��a�lEq�Qw�o��z���n��Z�hyB���Gf�0��h��5�A���؛✽��{{��o� �T�\��,�YÎ���I|�L��3-����(��>�i��O,�zoQCI��Z�'��8�����W��B��P������^a=QZ�?��aD�������:���l��ҡ�	2-fiVe>���}�˓=ށS�)��KE�Q�cN4����^�%�a��Q+E*�V3��t��g|ѠF��h�}lX
!�{�xS@��?�����=���eqh;�PPI �,��)H3R=O��#�A�?��O�	�1��F������a0��@L�n�_K����)��y�-x� ;�e�N��jU��zY�����qC��=�����V�Z??/ pM0����Z*q���;q�����2�V�����y_��Ayl��q06Q������WG1�ZC���o8�:���١�%jiad�f(� �[���ʡNO��9U>k�4��?A���we���~�F��ȗ��;+�>P|�G����ig'
 ��v�����Xw�=G���ρ��-f����(�sU���� d�.ΐ�:���o6;;<����`O;�n��+���ʼ���a/��Ǿ �{��lB����Y��H�U�
n���ޞ�>�ݧ_l�xW�=0�Z����D����N+���[��Ƚ���=80�3������hj�k򉧐O�l9��׬�03_�*�"9��7i�ؤS��q�h�;�ڄb�U�J]\��!��WD���eo��8l�L���[77���QCa�*.x�� {���M�
1:lJ=��KFr倀E/9���z�XSެ��C���5����L��5|���;�-Fʉ$����+��Q�@'��eC�"�i�=y�g�{7�o������XE48'����	-i~A�L	|�;(��=�� U�=<T��0�DhW�:^j�*� l��j]^�wN�YC=GW�����d���5s+��ޥ�j�
ifz�О>kx��A�'�3�j���ʡ�s��~�z�,(�Ko��
	D@�	>������wRB֯��@gcl�*���AߠhJK�w���U��4_�s��e�%����v@Vz�,�=���j�j�e���d4╀�_G{�����e�I�s1����G�X���~�M�S�Lfp����w+OT�z��=��UH�{��ެ�X�Ú��mI$}��H9J'��z�s�/$WSc^޾}c�^�b��y(N"�777�78�n"�n�D�L�I���I���<�Κ�a =2��{nl��[�ع("��(��(&�]��j7��j�`c[B~��q{/���2#��߾����o~g�߿�����Uq*^���Л�j �Fm�"��T
�	��i�E�{��sU�>��ǿ��>�},�uP�?�{���<�0�h�,Ξu�3Дn)����{ʖ���ll�b��7K���Y$ԃd����lee��6.��RЊ���b���i��bm�%P�;�.F8QP�+����8�v_���/�xc�_(vad�NVj�1ܿ�D�*s�����������p~$�ݚ��������U,�4��i�N�����7�tS�oI��4��uR��8���[f()YM���N)'=A�;�৵�8�,���E)ۗ���i_���6O��wk�� 
�g�I��`01����JL��5N��{&��l8�F�E͚��u���c���� �x�:c� �[��7��!p	��")c���j�H~���~��(#_�в�̲��'m�y�d����Uq-a+/.ι��S��za��S�L�I�K�k�.$�����>/��~� ��W���F���~�L������_\�~�^M.�/3�9��ᕻ(a?�F?#�������%�R;�]�bUl�+���T�[������9ؙ�7>���T!��>�����Ś�}
#��u�g�L�^�| ����V����r�X#�hN���\��7d������(�#M����.!��`+[�+���\��~n����i٬p���.�,�{y�o5M�1/@;��[�:��C�<T����ϬK����iޠS3CKs���T�1~�9�ݎ������|x2k�xL���k���_�bǥ�uw\и F�zR0��g��� �m�-��H��ev/�
�E��2��3{-�+$�>Y~�fTAV��D
Gh��\h��&@�xeGrU�]bl��V�����A:�`�)��ߢe�����[�lI��X�S�4��d|ȶ��H�o��q��h�	g�|m����c'9��i���h�Ľi�$Ǒ%���q�Y�u@�İ�w��~���v�EvH6I(ԑw�������{d��H�L@���nn��O����W�^%ٺ<;��ޞ;(	�+��f��ߣ�h�����c��P���h�����>`��!1�>74p��v��כ����lK)�Ħ�&����C��%j5��{ �mp����Z���f#Uf)���s�X&�Uj=w,��lﱹ�9Ȳ�IMG��$��pyQ;|_d�K:���Of�@�+?˞��C�m���4Á(��x��������>ᑃJ��7��r�P��ߘ����2v�k^$�{����������op�[���$R<�[S)��Fo�x�m�V��-�<����D�@���_����e�i"P�}uuE1�GDmN�ZR�ȹ}.�D�Y
�܇�������3���,]+H�"J���(�a�0����D���<��m��ٳ�\��ќٟ���V������͗r��<ͤF��#c
$�K��\�31�M�PUź���w���Tv��(:?W��v���\����^6
�������n��>d: ������pj� (K�ۣ��39?{�6�T�'Wuj��\&�����[�yL�:I�5P5#��c� G����P|c])����}w%�7���������u.9o)RԵ��XeЎPH�v'P�:՟��>�z��^�K�cO)ALƆ�\Db鰦�7c�ux�����#00���uWh��
 �J�U� IWC`M�_���ų{�lM|I�l�:�����wv�W'���4܋������%�g:�h!��e�F��)�p]��¶�~�s"���6�w#������:�mP��{���u�C����"mk>�ˋg����re��Q�03C+ d �/�r~<��/�y�~��f��3sJ%�#�V��/��)����ǵ)1{]�V��v��~�P͛(�H�@��~�E������q��uMo�nJ�O9|:�Nd���z�%��o�������\^�|�v�B���lm��"��g�b��|ov��u:��6lP5��M8�sI����o��7��J^������~2E:X��{��&�ڔ�Y��ó/�}��VkIZ�/�]��Js��=.*���%y ~�ś�(j#�� Ȕ�[�s��[Pl��km��=m̃謬�o� �e�*���D�c�&k���(P��k�:.nUg�X������qpMP�ŉ��)�:,&c�3�+N�wڳ�6CY;��QP&l�(�,�OO���ul;Gj�w�F��������Kf��w1���~�끵�F������_���l!q�k�ـ�1�(�s��	q0���`0�V�uW�8��f+����!�D���oE���z��vvq��fr-� DOG�����p���:r�{���XT ]j�Dd��F�q��)-�ߗ����	�Tj��>bcn���r��Zۜ��EX;5�-D.��
��|d�a�3w��#N�k2�.�"� ��^����;�;"y�=@�e�\�4�1Ŏɢ~}.���Ŝ�uȌBw6��a�'P,<"�u�K��>�-�����
�����MWQ�E@����J��̒��� D&��;g%J�<�^g��)�-݄9��!����6ЍF$D�эF��	��JF��n��Q�B��d�K�����	�sz\*�D�m�2�g2��G��T�>>�C��̣��J~��oOĂ2���R��S"�.(i�hO��@�+�%a�y��z,ϲ2|C�f�|=�P���	3���  `�	G	N����m���r�� lCZó�����I����NP	�TE��m�uBCp8�;9]L�w�7v��1�=+�"{@1�BC�2 i*�������o��o��^~��wrq��TI��0Ue�5վ�0 RPk)�[>�2A�$����rr�6G�9�����T�
:�ݒ����z�C`���p��l�ٮ�WB?�>O�Υ]�>8��
4��3e�N�UEFG�Cm���C�fX6vQ&0��0��e�����Cv��Ou��� �n��)��Y�LA����[i4�(MԹ>?;��Z�Xmu�lu\ ��B����~�[}�|Mu�����;��uŃ������x�D��X���"��ސ�k�D��sOz^} @�j^�J����-�OL.[�bj�e���pJ'%��dS��*ad����r����^�&����\��@�*����ĩ��))W��VoY[�C-,)�Y��  J����wo�y�� 6ߞAB��߹٬���������Ec��*��:�u�O4�-��\�>�[nQR����������,@���z����g���k�
���w�.[1+G:���@b^u��
Bp�7d�qM���db{�du�K�RdK&�F�kc��X��}��<�|.��[���, �ǻ."h<@ׄ�Ӱ�Tcu���@��Ĝ�zm���x!o����W���3f����ϫ~��rͺ��~���B��3f[�)��îA�{�i���	��-0^A,6
0v��u������[Ǧ��;�������g��x���A���S�������3LN�D߶�����-�&�[�1�8�lWM�󠓯���x���9��39>��o�%y O�%��v���?��8�[2¼ij�r�ݧ�%�E\�.���K�^����'�%>���������N��(n�Ge�w�}s�e ����2M�T����L��fJ�f=���czk�x2���	��8�'V�qP��bL�Z_kˡx��J����8:O=�o1c*�
R;+�t�d0�7�@�E%��(2�����%x¯8^�h�1_2�g"����ѵ�F k�����[��!��!�	M�n��K�﷚ ,�f@-�C�}wO�շl��~2��g�^��T��4uPجw[Ro��	�o�+�E��(!-��Ų�|we�D��Fq���1ӯǝ9u��JACz�Sn�����;y��J����ͣLԀLhM[DtC^w4|x���
k*@��ln�e�D6-s��BX�1��MF�c�z��ߔ��E��xP��`nts����IΑ+H�g���6�c���ǟ���ÿ��?�P��H���E�o�Io	�0KR/�5GG��}��+��hF����RD;8�9JX���\�Cct��%��SAf�jW�T���:���h$)�z|4G��I�j 4�g
�.//�t�ՑU�=���Ϻ���,�5g��G����a���n�}���k[���`��e�^�qiQ�A�����+Nw��W�/��سVK�Z��^�x.�|�������o����/e�%^���7�VUn�$ҘW��ͥT�dx"��u��� ��:�$5��p�Y-ϳ�;�rM�V��������nyAV�� F��C���{��P�U[s�/�k��>c18T� �'�2i����2�`X�����e��N�� �r���c��
�vP|]8��w�G�>u�oo�����bo����l�\m�B�k(����R�����>n�2�1�|�J��7rt��}?5�R7�hyM�5du+@(���"�{ԯybo��.{�׊�	�n�_����:9=!�g�e��%Z�x���c��A�K`��Vg	���e>*ʳ���|X�����f���i �5B�}��d 歷���S�T*xټ��E5ͳ4����Ц�e�̣�>y3���)&-��T��G&.�}���w �#�k�.O�\DB@����i�,(� �oV�N!Eۓe�QW=E��V���D�	��Z���!��{���9vk6oZ݉Lէ:=�T�����TC�����K����3Y"Fk���Ϭ�Vb��O+
]���Y-Q[�ӎ�m��Kvkw�AD��;3`	a�P"�J��&'�����˗rrvdu�؟�����?BeCۂڬԖy�iO�cN���F>��3�A'G��� ��W
ht�f��ڷ6�S������`bO��8;���S�0&N]��l4��{Xʏo����5�/Ξ�Ź�Ι/&��o��7׷�A���w
�W��� O�B�xi�Ĺ��+�c���o����&Ȃ�������K�m��P\�A!��Ȯ1K�,�g�XK�xO�*��`]�J �SU�r�����{�Oa�(��|���aG���#Wn��u��0���;�E�O0�6���(:��6̈́ XhS�:q���~��&���鶡����%�T�7�������bJ���d'o>~���C_%D{n�-�̔PUT�Svz���ڕQ� ���f�ɕ�
G3��3ySJ���+s�_�@bB��!�%�s��_z�����q��6�mWF�h*f�:S,�L���W�����u_^���H;���UH���,QF߂�m��e����G�	�f�>9�+��є�<C�uN��8�m��M�X���la��0�'�3A/��R(����c���S��R�ޮ���gDR]��>�g�f�Q`Y���X�;{�MZ+�~G�)��{�whY��3��ʳ榢_�Ȃ��d�ź�{���d�ۢ�2���Z�|B�6����<����=�.�>�an���@(��Ħ����1���^~aM��r��d�?����[�{A9���g��<4�E�	�]�-*?c�wd���o��c��Ȧg���pcdOm��bN�}W^�~M��ۛk�kv��{�q}�
�>Wb����uh���������J��l�И�f�i؟�����:@��5��L�����/���W��V��qGcL< BEP�g��IF�rjX��rq��_Ϟ=�"*�T��Y7q���o� ��c9y�3������Ln���n��c���&�#�[�O���F�K�Tߩ=9e؜��K��S�����3�iy��[�H�H�A�K��/eΚc�,(��I:蘹����j����^�*#>@~5W�w�R���z��6�P̎�/���F�����f[��#���J��^ʩt�?f�+��9����>��_L�R�ڬ�b��aPuV�{�=u�T��]�F,UOzfϟ����� &0G�*U!�k��mmW��J��NL��^�d�6p��bYA&h��o�r�8,��b~LP�l�v۳�T2����7Y��٭�ɳ@\8X��Jt�9==�O
]��"(������u���_Ij��޿�A~�A�����o�_��;yyy��A���G��F[�������Z���E�^���_dU@���<���\��Su���+0��	XNtN�����W����N�ߑ��@��?2���i�>a-�1(�"sw����
� �ι��؜�X,�#j��a��/��b1]�x�5Tj��:]ۉ=�`r@�n�o�X�1�bkS��z/tN]��lv�z)V��u�c���^ǚ���՜�r�[��nuN�򷿾�?��o���[����痗���O�X�6r��3-��`�?��?��w���"77w�G/T~���E &���vG&>��V?�g���;��ϟ��߼��|��R���N}�{˝���?��统>���=m ����K��>_+���][�g�_�䃞��?����O����uVx��ߞ���h΀|6Pf�D�fb����~8��}02�� F���
2����[(C���� 	?��@�����I|���-�����0cu���ܡ����bV���~#�O��щ1 J���t�,o�F?d�g`��b�s�FS��҆����v-ّ1ͮD��sMm����4��כ�7�=��B�6���2�Ԗ�)�����X���L9�ޓ�*�~ON7?�Y� U=X�Z�Q��D����� m�ˏ��$�����&!)��\�Ū�ݪ�!ci�GC��uM@Z ���{��b(�0��-JC��<,}�(��Fs�s@��4tnGS��3H}%��O,*)�>4<�5�ݕ��g#1D��t��9
�hz��	��
f�NhtG�]�h�z'u��M���$�����J	��8NI{���c���)�f8]d:YCK�D��&n�[k�I�3�so�-N����Ұhr���T��5d���q�) (���0�|�:J�X�4�#����==ίM�Tw�R����K��2u�F���t��o$0a���aV5bsJE��l)�+�����x3��6�Z&�H�{\Z���8�e7��4t�/..�����X����x�	 q���=2%њ�w�&����h�ڵ�d����!e�=�&3�	���(vъ"��m����b\8�_�_�V^�<�x%�:<�P�\�XMHp(fB�9��a�G3�W�5�����h��Xo����U�@�0e���:&[Y�@�Yy#���ĳ�Ƌ�,6��Ol�z/�խ�ݼ��"�|��d��,2�P��>�v�h4���e��k�6f-kIlc��=iC���B)m͆���iZ�y( ���2�������:�����|A/'�^>�s
;���T�X?�/McBF�	 z����=�S�Ch'J�A����Ϛ�d �쓅%�
xe�	l��7W���:��u<��y�n��h�s�$��6ۈxo�mY�p����n+W�{Y�l�0{�r�X�9�>bvDXGdN%�/���q۽�7X��r[a�i7 ��Ս�n����2���-w|��*�l �ۛ+6굜\��W��R��_����ۗg���	�ط�~#��/୺��@ �`�Qo����f��5*��AYxkl��ԛ͔~���gg:7�(�kzvzB�9�d����K��~�ѳK���GJ����� ��m�^�ޛ,�HD��xf�)�u<��[j~��z����^�����`)�������:�e"P�������f�=Cۉ*��
�o!]���k�ᇟ������5]���)zVQ�#3��5�L���[��w���;��ߟ߬ՆϤ��t���^.�>[�6 �����/|?�a�_�`v��v����B?�R��rus������!���~���ڨ���������Y���~����[2�fj��_}�w?�_����/����>��r�`�����~�G��7��������x�J��9��iY6��[Qc�;�l�j�k�cB���_ğr�N����΃@��y1��f��G��G�2"`~�(�R�3O>@U<�.Hb%O4��d�[z���BL���\��*�޾�""�(<��L�}��n8���P]0)"סq_�q��F[0,��n���&: ���h��ʼN��4�Tn(�P=�7�r��Q�ڍx�A022�rc�[�Sz^D���~������X)�{��>�lR�� `I0.FH:���g Y���O.oOs4 ��(��`�"�d�K�,���#�o�D)H_pp*d���Ⱥ�g:+����ڜ�I;#��N�Ǩ�T����"s#���=�C1mj����$f�=��PV]��fH"k�hױ	���	7�W������3�m����с|+�)�ڍ�\�n�D��g��Š5���� �I"fO��1�H8��8��>��b�o�sf"�S�EO��g��� il���}���mXʟ;��sAy�� z1�S�r����ʱ�a���^:2��:,'�(��#�;8��'n�	:�N�! g-^{���Ŋ����F] ����vl���F�����5��q0�G��cv�����لN"����٪; 	��,ZZ�Z��Ǎ:ڨaM��Q�Ak��@D����>O�� /^�����/�&m��q,:ԉ�Z Z7�)R&:�Rhܳ�E4\�����&#�n���ׂ2�_��UOSR}B��M@EP��=���[�鈢F�amΌr�!�c*a��6
�Y+�f��M��b�����f���78&�9	�# x��Q�(�j�b/���	���'3��%�O �Txb�n9W���{f��1�<�)�b�@�1Q�������a��u��<���3ifǔ�f/\?m�5� Q�B��t	�� ~1 ��2}��jp��=K�NE@O��:1���ӑ]�����l/�xT2�Z���ڧ�NJ�&���݃���:�
�V����=0�ތQ��e�Z�Aq�cmAdc���=�:�&6푳��A�bM�u��G���C�*z��O&�ۨ�B�^���Ă���Y�u6�F�|��k�٘�Su�?�V���<��.uۊe�c���ye�?�?�[D�t��
␵;C�Εs��+��vՒ.v4�5  �s���2O���\A���5��;��i�cq�N��NvF*���{6�}�0K��a�:sh�&3�v�L�꘠���׍����Y�-�Y�}lg���Z0��QAЇ�7����_@�;YL�.*�+��A�B_[���{�S`|�獚)=N�P�VN���-�!���ou>(�����������{-� �Pw~�i>,��F�������Oo�����p}����y�/�	�8�<��c.�
�n�V��:p��o���Gy��f�D�أ�葏hv|%�z-�+a�`{֨cE�����Y�{<�V�ӹ]�zĞ��6��R��X�N��go�S�Am�(J*�`���s䗐���gM��⎽�d#X��"WvN�Q�$|�Bo�"В�3�lGeu�T�M���Y6 5�|��.&����B13���*���O��I������t���_���� UtDPG��	���c�Y����k�<��Y��I����bO�5�9S!�:e}Č����R��v�ӈ��Ud�b�Q }����޼�Y���彦�β?q}ag)��~f�K���FJH>�$Eto��l���z�] ,+ۮ)Y�|�xd��F�UcQH�6Z[��,��[vg�&��9b7EC�b:��%c�U�~S�lM�5r��Xģ߶���b���]��8�ٝ�Hǂ"��vF��a�,����������qer������,8��|�(@_��z8f�G�S��n{�X�~i-A�^���G�'� ���Pה|�6_$��L�ct=����E�R%�a)x�7��� ���:��O��h%����x���Q���w�Ty8���.�{,�Q֙�&[&+��ϻdwE�zw|�:�X.�,V� k�-{�8G��8{Ꙇs�^"��p_z?�o�-G�Ԁێ �Ou���W�I9G��9$#�	?)�CQZk�_=�X�f�+�o>8�>���./������2���u�6����6�d?lvi�5����K������~oJ��ŉ LYdҋ���+Ҳ�P��T�I�)&%BY��rWցY�z4sC��l%�h��T~cC�c6G��֯�y�"��b�ݜ��5�+�`�W֦���:���UZ�އ���G
��Q��I�p�RU������m�g���D�0�֛�9���n�^ nJV���YS�&ݭ�
jhs�v��:��\cQ���7�L��B����L�N/�с����?,1w@{l����K02~`�K
�n��;� �m��,�e�`&�X����p�;_�PnÞo*�����������r+�w+uZ�*���4�޲'
J*�Z��s�19x�o1X�s-G�VH��^�0Ԣf��9]�|��+ڞ����/g8�kТd���72P2L������UmF'o޼�o^���u=B� ����#�:w�����/� �sq�$۟�����yv�5��3 yu����}v�`���v��W�-�v4Ga��Օ,�=�)c>�}�|��n��S�f��duX��ȹ�t�� �n�ю��T#[S�yݺ�jʌA1��G����?�,�'�?��Zbmv�����N�!�Y!���j���A>^��۟?���?���U�(��v�A?���=�2�u'+��d��-�!��<��ɠ���kv�Q߿ޛ(��w:��>����2��ف.�����c��r����<I�k)?��#�-�
֨�_�6s��{��ϯ���F����Q�]}���I��֥�+�{�1�[n��
U�nO�5�Sj_�N��5��;�g���~�{�]Q�+�O��l�W�~����������Q�� ���^�(T̒g���L,�S��;�$��CjLn�f+��OvU)5���5�&�:�9�U 3�2���]�u��L�.z��F�pG.��e��f��'�.
+�*X���&е�X6�;�c
*�t�"�����A�\=�WS���;��c�T���H8p�9���q��� �������OG�CT~����m߄*��Զ���ىC�n~ύ�d|�݊*Zm���`���fۆ¨��_A�"���dk�`p��f7 dZ�C�SL���^P��{Y�ο/��;�h:��1�zF�p��k77���HD���y�bE�!�G��;��@�Fw��>"��a��>�����9�G:*J�r���G��F��Ɣ����Ь�F-���=�
�~Zh�$P���S
�Ƽɇ�*�+����6?Y�nT���<P���{d]�����{��/ H|�}�D�	N]�����c>�o�m�y��f)��I!��x�^����qԮA�Cj"i��M�;�K�3s�v��'6&�_8�������бh�u����8��%�@�ֆ����;�VBr+���z��r�/�Ru�Z�w���[5$�6�c�̦5Z��L�՛7���~'�~�;y�����9�\��M�tќ� #�Q��R$�-ȆO�n[�0�w����:��"m_�\2�l��=�X���j
�܉oO��W3s83j�:�PBl��9'?��CQ���7@C��ޜ?���>��e�f[UcB�溨RY��"?$�y������)��h*�UV/�J� �}A$h�{],-ˊ�\��x�
�m9����ɫ>S卾A��|�j:Ν7nE���{��՟,���bUJp(ؠ⸤�1�~X�ڱ�FF5SmA���1���H�T�5���}����ؘehppE�X��@?<���W�q��װn�-@m+�p*�Қ�F��)�FPC{��F��K���~��Zc�w��Y�9h�G�h��auy����1���}�W���]���i���K~��r�왂�+������0�߼����?�����:���s�@�H���GV"+��v�ڰ�3z��?� �@aE��w�>�����( K
�{�ޅo t�����7[��7�B��D|܁�]|��l�F��N��JA���ѹ[�}`�27(�����~��s���B�QdbQ2 �'36�+�[���ύ�@:(�Ldu��'+=�GT22���,���5�����:a��G3���M�vv ���t4��GׂT]d��D6Q���Ú*�.�@��3�w`'dUu�빬�����%����DK��3$�� ��v�+yo>��dPO�8_1�`f�b1�d�w&wuuM�I9�ڲU_�~%''fM��~r�s�i��Z��(��R���5S���$H�!��9Q�C��r���Ɉa42d�w�_�`.��d�����C&��}I�{Z�5`O�+cʉ��Ԗ���F��~Y{�弛@ebũ1�a�;K�x=�X!�m��rYpdCV,J�g�k�0	e �*�Lc3�\��=�d=�dJ�����RƈJmwK��1�ON&.�zF�f(�ڒՃYKK;v��a��j�!��ۊ�LY}�jA��a&, y'�|���m� U>1@�Ե31�&%�����g�Ao/� ����B]A�.�����Q���t��ې�T�6��s(�q'��-�NF?AmBtOAIB]�~��}~"���L��ɚ�f'u� �{z3w�j�� { T'��S��6sD��b�*�a�(@�ֲŸ��N���C�C*��r�^~ US��{�ʢ�;DsNQץ��H�i���c�@��J%�@���*�N��FG� ���p���g�63˥ǅ�N�L�k��<��D��`�/��PBB�:r #:�`��d�HS��M5�%����SU������{�X����)?a^�p'|�y/�,Eէ`�l|��w��	2��P���g�����f��d��S�رa����U>�
�� ����G��H�J7L��!��2#!�D��?�ƀl(k�`V��=���F����X�B_��ǫ���{yv�����:6]mIc�K�+ 'cn�:�Pm���~gY]8�P"C/���(��/�$4��K����=�
)�h.���@渦`
�q�� �9�X��O/���7��W�7_�N�ϞN��.��\??�{2�B3#�7���P�#�Ia+�~V�N6�^�Q:���^}�-6�I��'���PTL�uH���)����G3^f���&ܔR'�����Ux��5�D��4$*E��$�ToP�:b��L���@qϬvc_��ܟ�7�eM�u���8)QK�F:s�c��\�I�C�}��i��`�@ў���l3˾MY{#,�fM*)��ʐ�����V�sTʺM������z��K�qD��|ff�U'�,���cZMOe�8�(Rע~�^V�9�
:Q[R45�A��z����߭tm.��~�,¶���k=X7{
���2��Fb셨�ڠ�7�ܑ���v$�7m<S��o�[s?7��ڨ�hF�U�~�"�M��y��M�^J�/��?.���7rz^���O����869���$w��<�����L��T
�fd��j�v��o�����rr�V>|x+�߿�s�݁6ӟI���ٻw���?�$W
|����^�B�������������f%�1��(�8�Y� �k[�k�����0�Cp�ǿ�]������g8��v��z�u�5V���^��fB�eB021��펙ί
j�F�E����{��_�.����|��+�NΌ�f���s�-�:Ai�Mf�Ԝd���,XK����j���ro��rEG��\u���O���_�yf�;�S�m���n��`��c�rJiW�#a��^a0 >�����l	0���7�}=7���h�"×B�^�
���?�R��������/��� h���O
�R����;h�ӵD�݊�l�槷�'����:A����냿cA�\2�����X6U��2!���(g"T��.���_�\�Hi��8-���|�=*Vmm�2�jc�UL�ೂ�8�C5�b��d���`�~�٫�7�>�+�ѫj��;�x��!콩'n���Z���:��O��ؗ���HOU{�m��ŲmkEŔYV�f�)�(�}|B�#���q1y\�pEAO��Ȼt�r�;��m����+6�����濇2K��({A�����j`$���'T�z�0�O@i��+n�0��e��r*�N�R��43�	����S9��٬��5́�GO��}��UDy�p�:v4 5-���xPQ'�c����!"�� d��@j��j�vpv��¸t���dzP&u�`~�v��d�xd?zsz8לk�S��h����z<�s4D��Yo�\�#�UY���)$X;�Ao�C����4��3�3fpb���"C�Hbn�1�E�z��c�;��F�����9̬������9�.�,B3q��������22Y���9Rt�{�|R�UѾ3�sT[!����w�Z���ɝ>�;?��`��>Wj�W�௎&���D�{(��]1$�?W!����GA��[���O�']������)��Mp||$/_��'"�2�1C��N�^q�q��2������a���'2����������څvĨG��R��YT��Xe�8���'qY�lx����HmgIS��0�8��)&�lU�ށ�;�����c+
7����B ul�,C#�T$�k�����Y��}db����j+�XЁ�@��� A7���FS�{�`i��{��>�/�i�iɂ���O�U���B��-��N�X7�k��,��\]?��j�:��uF�E?'[#+Lg��)�lÑ�DC���ę%Cso���)�����m
!�bE�Oآ`=�b���E	�9��on����'��񽂬+����vhQ;�������e����Ǻ&�����t�F�����N�?�3�t{s'��_	��զQQQP'�sk�5�������5.,����l�eژ[��0X��F[/�`![��������lۄce���3A
�]�����]p�̔d�"��s��]_��u� �˥<;�Շ�<���;:�''����|��]eԵ�δ��w�U�u��X�@�2kю��`��S@�K^+D��'Z6�=�v��Sj��x��"��ڵ��,Lب�{���Q���9�.���Aإs��/c`Q,����Z�I5W�����]}�Y��o�^��,4�.�f�y�eb8���~�JP��u������r���&&��J^+$C�|�;�eI��5=�����A�0Fe�d����=��JdK��;��Q�,R�'��k���Tn�)J�<�߲y�(,J$7��Q�:9>���F�hr��嘑"5��0*P� �9B5�0�l���SF�F���������f� �#�m��cJ��N��G���8�9��gS��Ig_V�T�C��]�)uZ�֎�ї$��_�o1*b����ǂB�É*4]�d?�s�8?V��T��9�vQ:*��b�sO���Eo�)�ڻ!��P�?sc�Y9ec~<�z
��B�b',NgJ�y��TgF(x�ub�{�@j}T�'J��P�ٴ�T��v����n���SIk� �\$��Rj)zR<t�J�a���@�B��6� ������*�x��ڼ	��OL�Ȟ��I��=cd�/� R�(�������j5��f��O�1/��qX�����aFռ�T&�w���!P�Z���{<_�Bg�B�]�����3���J�����3h�f�\{o�t!0@�����?��< A'���|R<z�l쏕��l�H��e����z��y.�'��*o0�5G��Zӹ��Sy����x�J�Oό[roFKL%���<G7᳓�Ӏ��Ho�mGGx���2*@埯��d͍8Y-Y� ��i�����(�=�iP��XR�*�UrZ��������֜��\ٞӗY5��m��y��;oUE�0G�f5����S:<wD�:���t�P7�g�.Y��b�Ǎ�~�/|��g��� AD]K�e0����1*�y,���� ׷��)��'kI��*��\qP��j@��Y_,q��_�#���P{L'ګS�!y}|Lq
.�|R�kd n�ۖ@J��0Q�9bua^3j�~���7�,�.���w�P�C{������WUims�;�{}�������۝�)����[�С�M�Q&P1klnH?�����Cr�umV�4�j�:[W�����j;���Rʟ�S)1��L��	І���l>���'��;i�;���������|��=���D�T<D��F:땙C�&�~�c�NoeV㵺�	��V�<���g,�r�4j[��J�dL�����S+1_�y��FA��<�Ǭ���Jk		�]�A���f@�'J
&m��8֠~#��Nnt޼�i��������{�������5��t��ŧ������|�,#&2^��|��) +h�n	F.M��}3��J�d8�!��w^{%v>��c�v ��,�xb,0H�H�w�N0K� Pg����+� �ѷ�E�b�J&+2Uv�y �F���d�ƹscݿ��<��xo�J�@�mt��R��6H�Fv��⬲���~�F�=hĊ֪��39N��1��}D��i���'<Z � &�B��=�sj�E�_C���>D�?�8D��W�B��v�����_����H�v�ĸ!�F�4�?�(w�2��<�F�L��Ky��R^>?��g�QPC�^=(���{3�Gt��cr�tgr�8_DTB~�h3we6������sF`Q��"�K
M�*��r�{�6{�O;9�e�S#GN�$6�1���F�N����
�ɀ\�Z�vos*k����"],�Zh��"W40���~�⦌�z11��p��Y!A�h��e�'o�g���q����*�$�:�(�?��9ԸF��'/k ��ѭÏ�'c�&�h��<����R�\ylD���(�8�6�W����2�it(N�eޗ���ʚї�ā�룟N�v�6ꘊ�1u&���9_y�cSg�@E8�qoz�P��`<���7�&[ ���Q�pH-؅���b.'��|)��-�ļ��BW*u~	`�#P���Oaz��d^���gU���5g�#oז��'ҹ��t����ζ���t�^E6Ν_��`���j~M ��'*qu��0G<8d�,�2�)�4	 a�����hӝ����銵G�ASm��%�6ǘa�-�H'5��M:|#�+sK��6�Olߧ����B%ˢq�|r݀%�����k��w�{��]��ku�����^�[�ɂ���ł��F;o(lf�l;���֪T&!MUQ�{hJ���`~@�J���h���\�Wl6�*&q�o��X��.W+�I h��%�U��ĩ&��"8,����&Ң�e��M��N,c��:؛Iσڱ��;��P�N7e��*2��ʢ��@�� �G�sԟ�� ����W��[�xjHJB�1Z�P�̚�5hE�a�
���RT��8���!�0���XV �Y��u�(L�Z2�H��ؒDV�h��k���ƚ�r�d�;g �ֈ�Of�w:^�-��T�\Ȳ�6^�gC�MeZ�:$)�p}T�����[���񄴸�
��,`�D6q���dM�֚��:�>"���&5CS�wײ�>H���NA�Շw:��	ꋝ� Dq��{U�����ܶ��M�9(���� d�+��6ՠ��)Ab��÷�8��� .\6>K�����^|'�d�샯�A5��N�Ć+�Z���j�2�Z���k���+����`��n �e��P[=�i�� g&�Y�K�'BJ�Τ�͙j�X j���w�YW#$l��s�HLdJl���6��gQD�!�.��g��O��F9���)�@��H9�ݨ[��� ��D���߽:[d��C�Q�e�W��[�3���0FN�nU�nf,�6��|*'�
�./���sy��>d�8Sp��fV�>1�f�ƪL]�d�ے��m�N��E$��"��gO�P�"=���)ŴӉ�ӎ`�W պ�<_:s$��@�^zݠd#�z�@�gM� ��Sٝ��$��v��YsKI�n�x�Q��hR[�7_��[6��(�ܡ��d�_?���Lrr㈉��9.�u��?`�/K�L��D� r���UF��b�c��a�?��嫟B��s}q���o�1�r�z��xr�t�W��a��&�6�^�?T_�8�Ӆj�v�r*N�s������)�A4
�D�{��{m� $��#kI�ȊX����o�`x8��a�0Phۢ�p�d��F�	dݡ��3�q�;����7r�N��ٹ���q'9/�F�Jf��k��0�����v5��~0�F(V�?0��"�10]+҄k��u������S�7�=� �^�Rm��D��}o4���.�B��� +�Kq�\�Y�(�:3���bCҜ'��`��y���K�V��qC��V&�K�Dv� ��ug�HR9�k���Zg�ڹ'iCsL�������څ��`BMYz����Hu���5��}/���\�n��f�:��nF!�^|z�Mx+k"�}uh�R\�R���/�_s?&����33"z�������٩<�x��$��g۔)��@��S�5���
zjOH�Ē6���ɦ����nvE�A�*�u	��s��a�.�"��C����h$ h[�`�?C� ��l~�������r͊�BK�о��z�5�4��a}�. �HQ�L��g�S�z�{��}��yd��l�Y��X��g��I�?����@��`B��b`���)��N.�SoIc�2X ��<�~���m�^��QX2��)�ǉ��NP4	��a��;�c~��V<h�%@���d��zݔ�gS�����bf�<K���X��X"���Y��[m���= �V���5�:e�2x�x�����ń�K�^����u���B�t������ +9['��-�	dz�'?��$�}F�(���T��R
⛌r�#�*j��%c���m�{����d�rA�1}n���0�`�al��m�-�pv�#�J2�r,|g+A��9��pP[�{�uq&(, �r݄Q��֋F_�z,�&���dbH�G�����5��O�"�NC��2ZC�Tq��\���p^�/y�������(h�c���7��� B�\y4���r���~ɤ�A��ڙ�E߭%`�FK @�(e���~)5R�sS�Bϗfjz*�5+58�����+�����ͥ�z�L�_��Ѣ6.j�30�@�ʞT��4��"TCAUA��zo��w���x��[L ��B��T;m)�=��و�k����
Z�?������������=���W�t��rw����n������,��[���"�`���H�D8�U��ފOA��2Oe�kK뛃]2[9��yt��ԯQ�>�0l2Dh�؍L�`�"C����_�ȣ5p`2m���K����2X�(�jVl�T-E�s�^d�7u��1IO7���gL����cgѤ!��͛7�6^���m�@���t��~��c�vs������nd{l3l��ʌ2C�XF��jYp*v Zj��1Z��>�)\��Ӳ3���ŉ��g2eVc�"L��X_8
�1�*��6U��˜{\�:�9�-&��\7��Dm"��_��ǐ�q��D�٩95��rΆd<��خSZ��ܛ:�	\@���S���vԛX�~突�����wlO����)*S���(߻�)���@�%鋖�a�kD��dmrA�E'�L=H=&�n	{���]�<IQ������<Ƶ� Ou�f��{�z�
[��b�� h:��j-�7;y\"��ń�$}8�������C�+����;�(AC(���T�e��@ ����2�S�q���5��:�'3*l`.%��P��׆��`�@����ޟh{3��np�IQw+�0�`�N�|\B�tkv8��	�}KY�-?���)�H-��!Qz�F&���'�Ί��Ђ@I4C����=2�[�ǝ�{w�:�T��!����4
JD������A�5Pptg��4�� ����A/�o��Z�������K����!�=�VT�<�����0�=���P$��� [L�X�z�b�u6�Dj�i\R�=�ؤ���o�BR���)�b�Of��Y��8��;~���k�w;S�e[�ɬ􌥤�������΁����,)�������~g>&=���d���]m���Z��[\�VSP�Vp�Z#G���q`Բl�8������)�<�"�Uz�7��Y.�v�Qط�+�ѝ��}��_� �Hd�a��X�[g�����Ye�-wVP�$�zok�r�d�t,� X��vR�ٹ7lpʬ>��1�0�C_��M�i��7)k
������F��dFr�0R�a�2!�:,��R�	��Z��8@i8>f�Q�Ψ&���~2���z3�t�q����hY+���'��Ɐ1�6��z�@c�$�K 7{��<{��Xk���S��=�$2Wh�V�<�5uU�	�&�>nGs9>=���S�|�L^������������Ζ������WflG�.Ԑ����������t"��eX�}���P�Z/�s� ����d�ک��Ŏ�0�6�-$b�Rd�h�������:���S}��>^�����������{y��&X���[����EVѤ�'����5�S���U��ϖE0.�-�쑭�?����__�����������j����{��'t���|x�\V�6%�`P`�x~���̏e��s�s`kT,f#hLk��o_�Eiѕ����6*{
��9W!���_�w�}'_������_*��� ��rY�{NA���A�#Г��}P�2 j|��(ًŬ��)�P�kRoզ.�2o2|C��ğ����͑�+ȺԵqL[ ^{a�I���32XA%��M�M6�'7{�D�.6nryw������ �_1&��Q��RP-���0>�`����y_�}��Ӣ�A݋���֧�7L��p�F�p�[o�s_
��7׮&'p
�@4ή�(:w+�,��R�U�}r�{��izF��5F[4)�$G�a|����9i��v���=$��, ��2�&���v�l������J�˲R���1�mj*嵽:���_D�� �i��f�'��v���`+l|�"d+Wv�mN��L ��n`��C}頝�<F��b���5����"ej��ԇ��2���6��<[v�+�Yo��$���8ǡ���H�mK�r�̄yK��U-��yCt���&�ߥP�B8%X���{P�@�7g!���b'�_<��ť�~�(K��`� K���2+�
~Vbh�=s�{6=F�2^���Wۖ�,z�}��o����^^\���Q��]��C�~>?��T�]�M��f��4V���L��'(6C�B7����F�k�j�h�p���p��ɳFֺF*��Wm>kH}�zޢ��5�&Y�ɥ�;��%8Z֞6�2�m��������4s�Kȸ#���k� �� 6�y�W`�۬t?]�5*vC��Y;Kۯê>n�r��n���\e7y�� ��O�K R<����@����u�yZ�{�� -����$#*�AI�Ƴ��c1��;JM����=C�B�6E-��tn��� ��i�9�zk��X��iwIF�j(�F� gI�ގ��쓰��	�9^.�LG��,�}�P���d�"�z��P�h�'r�fz���a�^�z��\��8�e|����^T�խq����'�b��U��wiR�7�Ɣ��;?��Ǝ�1AdԴ�j�&�eve�]s��w+�۲�0j����kI��g	�ŝXy���DE � ��]�`]�������XNO� ��D�1�(�b���=Z�ǽHn4!��L�n�+k�k@��K��y�^dJ�����1[�I=ؐ�PUj�7Ɵo{S���
GAch��,�nL:��Of�\-���fǼ�����B�B�� ��޵��ot�7�4�<��Μ,-q����~jTxr����a6�Z2�6W�
	�����_c*����3h��?�G���W�Gp�H�%���Xt��ɟ~}�P)�)����H��-�LA��A�����n���R?�*���g��	�.zs�h���6F��o�PO���ꫯ��=�̾4�ޑn�G�/�1��Ӹ�ml�ݎt�	!z^�Ōv6~9�(�Bv�9����W{�%���=�@�e��Jag����q����� �!8*�B��4pt������&���"A��@uY5zXE�3iX��^�Q΢��
WCo<�� 2�5.㜝�Og�v0���11z��\���-ֲ$��,�h�D���,�eMĥ���<�P��Z	q�S���ԧ)Sh�ޒE� ���E�#-�cR�����zd	�Y7w8��sd����0��ڴ�����zP���u����1r����怽q,�l^�*�<���'�G�?Q3�Y��z#�-E�O���f��P�5yo��>�	�Ud��h��&Ԧ�s����3l��Wy ;����S�}� $O�1Z�e�6(���{�K�+�I���2K*�ܒN��qN�O^�\�d�6���D��g�@���n)��*�\9j�'ڞ?�;��k�S����9�{a�e��������Q;������A ��d/k=�>��^��7�+̧�d0QHm��QP%K�]�����W��{��'�@�fK����B����k\����XR�#�Ƽ��X_˸���� 86��̖-����~�vC�5gb� ��l���>֔۷��TD�
b)A����}Q�w�\�1!��Q#�a�ٛ|Qp�ׁURT?c>FK�U�N���E���+��Fq���w�k4�.ZA*y6q��eV�S�'�
�WS9��c��3V��:�&�D����ёay�(����&8�48��h�i���d�� ��ܭi���9d!�y~��|��Z���䄀jqdM�֫�dp�^�x�����a�SA*��U�=BalP sO� �=@�p�^��Z��=*�ҋO�V���S�t���{��A���"�w�@�k��B/���f�d1��Ts>���'�\��W�.���K5�Gl@wt4#�yF�@z+�4("x����:f$d��(�'<�;O��#�-NK�]t�"��?��y�@�!=qo}(��3���.��)r�Z��bX�
Q%Dd���N�r~:�T�^���P!᜚3c��q5�Ĭ��:�]i��hNޣMSP<v�"Υ��y�1Ǹa�C�_(��L`���R:D���)�gr��J���?h�bDu����If�q�Q�_8�/���������{ �(�GT���
�0���ȶW.6`kջ��sP(��� �<b�N�=Dao.//����!DCN���b1���|��˿�����=���T�&ժ䓻�*gSQ��཮�r8v��������W�=g�	g!�n{�g����)%xt���/O������O30����/�Дcr�к�Ao=є�Rr5"��ʵۜ�l|��b׫<�CA	p!�<�M�eHg�����,d������嫫P�uF�;��o�қu��~,�j����	�R��舱�>+�Yf1*�U�$%g1�z4�b`�rY��Z���DFO�Hr�{o(�ZM)�VG�CQPo�j��ۻ� Z�]����S��4p.�Cx�!��R睉 �i=�S=&s�ΡŜ��"`rߡ���>��{��aB��A��m�1�!��KF6E?��Ё٣��s�C�S�{�|���Y��#m��}"��Iu��P���:hGK�ز�q��8��gTM����.k��\ ������s�3��~+���k��%�3h��CD$��%�(��^ d�(K�v���ĸ5#� �;jL̂0�XQY�Ek4��[��u�h��-hL3�l|�IC���
��Z:�FJ&�er���>�ln���.Ȇ�UOќd�2,؍L9�_,�hx�=����Ֆ����9l����t���i_]y�t��q�/�d��QuoT7�p�n>�f���BP��M�V3��,���Ϭ�6�[<�5���ux2����!���ߐ�oĩ�&F��1���fk�>��V�DhUcO��Z�_���13lmc�� �⁒V�B���*���
�r_ф�i8%������ش�o�TeB���X���r̽����x�X(x~��o����^~��+y��� ���E������0��9����/�	�,|�}����8��UR�W���������*Ǹ�W����F���h�&n�������pL.�mT�/~n�,�5AlR��$zb�/G#G
�������K��z}� �RAl�1�3�kQ��i�K��f5�T4&�%��"E���8�p��@g�'1B&�u�^9}��L�R�o˾V�3ņ����� ����@�o�<���":��d��9�R���B�)�\>���#��;�s��0�F}���^�vB*�,J�2L��{mR-���<�WpJ���RVt����&��xf4_/i�����_��t|ί�3@Ir؉<L��H�\���Ύ(��"Bj�A뫽W�Q@"c5P#(�$�(�y*r�~f#� B��;xτ�3����x?���<��T3�"8lY��� }
El����R�����~��)��* �e%���@�I;fq�6����%jZ@F}f��:�|v{^����¢_r�G �7�x5����8Ŀ�G�_�9p�^M>/<CTU�O8)+��|��{�:�J�}tj}_�O���Tl�k?�ʝ^;�{�֓����ǹ���q=ք=�j�G[8`@Q\��3����c�k�(1 �61��&�e`ҩb��;]��<�������� kX�=� H��T�����L��Nq+7w[�x����=배Gt���2���+����)Qƺ��{�+�����K�"�i ����QgǠ��k�I���j��m��Ojy�+(�ݐ�h�j������8!�(�-��!}�Z-�W�WN���K�Y��r��3<X�15�{P��Hk��FM&��K��De�t���,�MK�
��x�XCF�_��J_/(��x!���;�A��:j=S��]�Z �)�4R`uЈ@�sՂ%`3�y0�6\����[�������kvݕS�S
�K)�mLl��0l�T�L�)W�ͱ{a3?���׃U��������=M���.�n��A�z��Ei4䙎%z�e��7�� %3N�h̍���\nv4�5 C����	���b����څT���l�p�LJ�BL�/�%(����n8���fZ��a6u��]�I�d�Q�5�fq>
bJŇj�x�xO��}�
�J��C�AO�ڼ�vM�������Q{���s�'�\Q��]��i �)�K�uJ"}��gA��s:H�Ή�q�
mi f�#y��|��o������V���1)�(����b��J(�pv~�Ƹ�p֧5=�z�L	z:PТ�>0�3R���C�c�cT`j��,%aw:���Lf	�z:���["��a������'Ql���m��DQ�>��}��7�Y�E\,*5��Z�G�Re�(F����[
`��O���X�x�B���|�����%�ƱN��JՐ����F�D���>U`�^�����Z��!1�Mk�{믑<R��ߞ7S�������gl�g��He-���e�FϑvAť�Z�f�('EPP��]v4�8N]�9��P���^7���.�}��5���)V��,����h/��'��N�����/�3�N'��{��E���*��&�@����*�Nݜ�D�,S��@R�*X�ٸ�h;�GEP�g�"���Yէ�~�;�~�jd4R6ޯѱ��J�ZN}1:�s���4٨��e�(��QE�D_9�ö�X�h��@�%͟�o]�-Kp�ms�恹� BvEɚ���7!g�@m�Z�׍Z����S�F�;����qa{�Im��p^�z,�ҙ��%�l�:gK���=k*~-���B��(���_0C��%�O6B/Cg�x�i���B-��"u���Ok�m\K��`��J�P�ˬ�B�z��i���t��e�s��fI��j+��T:d�����a/'^g�Z�c
���WR�kG���ܻ=��a#m[��0��عxĚ�w��N�;r�"�������k���57��Mڼ�ё@�m�K��=�DX�7Y{}8���;d*�;|H?�y��tZd������z����^X'�^�PP�u��cO�֋�unR~��T�v��a|�`fT6�	��������٣tG(k��w���Bx���2}�C6�D��I��q�T��C���	���[����(���z��bq!�f�,�nov�㻝���ɝ�˭�]��y+�L�:+*�� � ��_G���BO5��`M'uM�M��a�̶��S{�#�LxO�9��}�`f��Ǉ5i�WP��	)`���-�hg�x�]�3�T�MIx��Q	���R��:O��l)w�
�օ�����y���9��� o���_C�`π���)�y�7��9�����kA�){aJ:����+f�����wo"�=��{/j{/��C -{NO�..��;Oh�`�t�����Q�m���M�=T4��U�ǼY��?Zb~�KS�������wP���Y����f
��)�[�1Mi����Շ��x#�
����u��Α�H��6�3�̙ ��Dk�	�����癢�}e���S.��7[�M�"К���ն���Tl�V�	�S�h�
�U��#4{k"��Iۑ�|� <_G?Q����#fې�k ��M�`G�j�S�FMkK�*����:����>l���\�k,} �q���s�M�,d�f��],��V�A�ւ�p�Q/���~5�0�� �mG���*�s�}[�mD�30E�b�s�{�����[
V�Pů��h��}���F ��Db���R�=|��5�k�y"p��lq��^690��q4<���t���'�:�OJ�>��A!�*78�T[A=������ȿ�ۿ����
����FH01�����Y�AHi���}##���,聣�N�������fHu&?�X��p<%6��������6�֣�HGz�a�~Y���Bb�]�7H�8x�7��0I��E�������卂-]��-��/)���������J3hn�0N�.�χ%;����d`T�/�XH>m;����r��n+e�l5'}o5�~� ��R�ɮ1��0��8QA��t>[ AY
E� ��Ӄ�5�V�z=>��fw�N�178��k��hO��/�l{Z{J���c�o���f�xO�l���9�enl���=;�~b��"�X �+U��e^����FY������8���N�����A�;�VC�}tM�F�{�N"8�>�A�Fp){�h��~�
�^/�a4�f�o���� uP �~�Ѐ�uww+���rrz�����@�܍�9�T}��2�ޟ�y�iq�}��b�ʜ)D���H��8�)� �]P� �P�@��հwt�Lb"ш������emw%=|��G5�i��z���_K9�R"W��X���B�n���#�WILz�9�ܠ���,�p`��}�+F��Y<B��䔲����8>�=m�B�����*�聞�+ �60G7�:yw�׶ٻ��}�K-��l�x�������ŉg���;�V�6���ۏ�pvˢ��0s߳$%	�dx�?�H�����#�6p�ՠ+u�^ɺ��欗��N��������:��m�5 �>�_�2&������C�@������a����-����Q��#sn�fv���>������xG��g�B��x!���N�c�3 ���/2뫕��1�e�.��$(�^��vg}Jf��?ko��H�$	��; �W\�Y���N�������0��U�W�<@pw[UsgdVU�~���d� �n�����(� J{��Be��&E��`�i��@�z�M>ߔ��Z��f&څ�c�޺ ��Y��)UQn��.l�k�Y(������Fr�͡�$�ڎ�~@2@�x-D�����f��30�P(D�������^ �@�[��������s��7h�����X^��/�K)ͽ�UL\�f�A�K�K�2�5��f?{�ˉ���=(o���XWK?����BbE� F�@��i����`����]يZ�e7���m(��VV8�w�8U��w�a-Rzl7�g~^W����
ۉ2 ��(!т�<���#�x�p�R�� b�|�c;<8&h�����U�M?��c�l���Z�n|r�Mu���5�n��(0�U{�A�s�W����v$@p���L���|�3����_b5��K�������6��`@��fގ�S��ZK�G��i@9	��ݷ�ٟ��*�"���N(kE�q(A��g���px�I�D4� �Q8?[������������֦L��T|7�����Yp�k�P"�C3�����(M�۴A�TS̃2�g'\=+@�=yrn�'l�G� ����B`b�Pix[��/ �h�T-"*����HQ�EB�)x���J���R��O�]G��x!aJ��=GJ1ZS[✆\�[���46o�-�8j�nnnY���;�`�l൬V]ٸ�<��m�7���Fs�
	g�-A� d�-��4H�J�@�jK��H���-�<����w�uU͝'�.��7�^_��6��:�zg�e���nr����7wG�Ȃ�T�_����Q/�{K��Wiګ3g����!���ݍ䒋SB�pR=��=�����,(:5�t� ,��E�=�1������vv^n�`9X�(g!��sm�f"��'͵�j� �I�#mԪ�Hۨ�)#ޭ��Fe*$��&��C�b���I�詊G�^}�U��aZO^c;VZ���/.6���٣��lbs�����w��{��&
�׉�N����^g!�Ng�wت�"�(R (��G���а����N��<;b���Ș�?8�eu^�ߞ��f��j���kF�!�}{sm�W��sO .���z�*t̄�j\�x�L�X��A�F2㌨�R<D�zo�$�Q�36��b���_���LϏ���p���b���j=�|�?��,��-Z���-������v}�a8� X��:xZhȌ5NK[�+~K:�Uëj��
��H4�>I$	��6̗�k�����{�-��R��q����f����o����@=�4�O-W-�<�j^X���a�#\�������!H���œ'2��ˌʍ�D��¥�׫Z�W���D�W�s<���{�����l�l����;{��--�����Y 2�����괰����s�Ө��vP���|(��fJ�}�����&Z�9I_�Z ��f��t���tY��\ǆBF;f�v����"UY�g�����#k�s=��|��
ڵb����_h��?@ufY����
��@��i�@z~�<� UZ�"P��Ulb�,�`�n2����/�!�Gk"��ֳl��n��V����lpMkt�"��D-�	�$~r�2�ծU�<��D�s����
��{\����5P}���̀��vY�~}}Wƽw@�x��.�&���)�_�0z�\�~$*g�͂�a���#c�kC�`{����I��sC��'UR���O� <R ,�H1tcY�ɣ
M:��Y��v��w������Eqz�����Y�����P�� %2�L76d4�T���T,��c&�R�2��&�����|�f��i{�M�&�Ҳ��:�Q(�:c�	h�a�u
�8W_`�RP"���9���|����c{��ܞ���&i�@a�~wg���E9������ȼ|����{�Ĺ^n�P!��hMm2����r�G��a�����,�7�\6��J3�Q�x�@��[�^��3�2��4[*���)y8���wtzك�:(�{n��vG����2(<���Ég=X/'Z�0�$N�(E�e���[��X뎄;1_9��߉��l5��+b�+���s��b�#���0��;��:�4et�b�ړ�Z*N�������~Ĳ����@�z:Y�JLNt�NO�@�:C��(kH�na͌%���Xv�ӏ^k�&�Y�S#n�ͺ���j������+�{}��>~�`Ϟ?�gO����"{1��:��r>�~L
o��`2q[4*���'i���!*ۨ!x�����@B��};���[�m�>(`t-!���a�co������袏C�գ�Ms�w�mfVE�+E{��j��/�������Ri�[y�[㸡_Ϯ�L?�(�F���>5_<ynO���ӳ��P�����ߣ�3?cq@��3 qó}J�.������������/l]}�X��'[�ݖ��*R����I�d$h-�B�6NOi����<�ݚ��DӺQ���Ȫ��05 b����Y߿�d}*ʮ���b� d�����UX����*N��Y�vD�l��-5"P��T�NM���r��6ov�M�8��}���k.��%����0(w_ ѡ"�pj��{��) ����!���O�5����H!���l�΢W��B�^�X#���E�-�A��s`�6�W��G����=~Hm:U�����Ÿb\�4��o��*�ߺ���?�Ͽ���~���}�Pl����A�0��� d)��������2��*���o�l��|Χ���/?�/�����NG�����EǌU,�{,8���א�G}؆A�Č�8sB�s�[0��ځ�
(�[dJ�L���T��Ӑ�̪�%�Y���� �-�a(Q�8)�������!t�Y��-�FqM⼄)����#K>I�l��P�����8z���>O�ϙ_;�3_�uEDe���:- 봀-H�/�;�ڹ�BC��8���Y V�� Y��!����aK�RF{t/�sa�%������Xp%ʼ0�=0x�0/��`�hĢ�;��yՈ��}[~�kt�v�H�|�շ�'U3WJ+�j�@�!Q牡K��������1����4�t��݂O_6���1r���<0K�ȡ&��by��M*HkB�!E�g�*�wG#:dW��YU����>h������ �	@5��	di��$B����,6NPds��\�wOS��<AE�@�:=A��R���i�����ȳoe�$���Hj2F{�W��gd�s���!vFidf���j#xǃ��39�E#�Q���M#E�Dհ��[W�����g!��B�ԁuv=��w�f��Ȳ:t��[D�*������fӲ�&~Q �����H��fd��f�m:��霈�����5Q��IT�����4��+Kkk�7Z�#�̦�(w��DC_��u]�x�_=�?�ƪ���*�I�=����x��ִ�o���Zi�d����Ve_�H����ý�Iu�Lɷ�o��eNwqW��c��s��!**��s5P���s[W尺g�Y����<­@�����&kv��#)�b��l|a��(#��J4��X�]�`@�zJ5�H�Z�����bc�W�����n����B��A��ض".>v����ү��U��W�	hW��f�;��a]�7������=\�����[��4��" �FV��*�gAv9�Ϟ<��/^�7/��Ͽ���3�k���2���k��)�?�]Sq����ഫ#�?>���/P���}.��Çwp�����m�o����%[���M`�ؒ�^˃(|B���6�7�Y_[:#/u�;�� Z�|�o;ӿ1�>?���)Ş֩6�.&/���*��DV�8������Kd��v���/�&��"�o� ����c������T:�Q�2�qvF��a����<$G�FwF��I�����A k}Z:D&�@/�[P�V�۠RM��:V+ 5�Z9XU=��;f�$T��ڕjF�-��[ڬ����r⅝_\�m���ϗ�Ŀ}����Ȩ��cM�-s�@�rF܉d�`9�$�Y��|���T����՗��>ڛw��4��p0��x
�3�Pm�ZȦ�}A�۩=.�J{<�vW���w;���؟�t^���d�	��,��r}t�N�s�.b�TEՃ�L}/�d�a�ŀh������^|��N�d�3,��T5�iK�E��a�1��g?K"��%�"���Q{�����8?!��Y�HL��\�l$�����)���/��n�[�k��?)j��+��%`{�Q�Y��=�[B���}0n�t��}`)������ٹSx����������Z6�N
 {���R=���@���5�dr���M�����w��ly���5ۥХ�y��x��3߲j��<2��P�{HA�ՑA�@�o��(��%�!m�kPK�'���W���|*���Q7����Z�jĦ�F��Ii�jT69ؒ�hn��qʩ���׃�ajD\3v3�4ٯ�"�@���Ӕ�E���������8d�,�f6��+@�ķ�6�^��f���h��%�V�@���`���6/�u����s������pѝ�l��C�z�;(�y�Q��GI�e8�x�~T4��~Bo@M
���Y�Fo�W��f�jM8＿~�Z������2�Mj�`��H&Xo���f���1��@<"^��N��`�����:E��su>�����C������A�nΉ03[QV;��:Kq�%/��W�zn<iV����Rp =J�������b�~�LӿF��E_?\U������xD�x2,�?�}�}�R5\����U�1�ìoͶR벃��師|v���5C\�x�P�P����8�TC+d��N�^1�蹂5�P-�Q��|��q�|�˄%w08'�M<�Gg(KEɱ�v�ݖ8j�5$%�}W�h�cZ�AX?]��/��w#��8m�>=8���=��[nK]Z:2a>���n��E@��湀���}�5pY��T�d�0DG!���=}�<}^~��x�����N,}x���GK�3@_=���)`�WC��G�ٷ�?�g�_\���ݐFxE*����p���Rs�*�V<�������v���YX��4���NN�o�#K�4u��g	x�{tPJ�)/���Uk�*���͎��_n��{��.!�5��Al�&(�`�Q�4���:F��~'{�z���s=-���jlF��Y�s�1G �Β�����9%�����}�^S��/_��������ʀj]㙙e���R9$��vD����#�t��{�c��-�����s���������=��vrT���)�����޽}�L��?7��1�!
YUq�2�ȋu$J�@U�'P!�1,��PK��=k�n�X�6�.6����f�j]p:��w��m
vDH�{���;�Ug����޾}k�߼�?|{nϟ]賲�� ���X�3e�:g��)EY'ґ�W�{���_��W�SrM��6���S���gg*�؃4c��3�&�GU�@V쬺e��p�+P1?,�^Ma��@8k M��z1J�����w)��E�������k��d}G��{�S��VK�\5m�-�\��X��8<� �Z8��~������"�M�^�1���3U���ey�z�)~�,�\�8EYL��ϙ����=亟$W߸/2�d�l�WZ��G�����p^�s�Q��f�-=��[sA��Mnlռ�����������Ϭ���qrz�%$���%2��]��M�lѸ$��S""Vu��)���2��A�D��p�v�W?�Q��\�T��8�z��"�6(���Q�F�c�����d�~(Q4j�Bμ��ES �,����e͛�����	-�� ��R3>Po�A:�]��G��=�Lc�%uqgĹ�^�W�_��%�L�IIJg;�Ħ׹׵�x��igY��T����Q/��UT��(��(M��墍֭"S#�*�.W�_��r)���#���Y�肭+��	3�`PXm��N����Ѥ�F��~D�������\te8�xd��A����гWU\�ѓ���t��Z��gl��_=&��!��k�Ș���V�&���Ĳ߮F$��#�Ը���a�BXƬf�߯ֈj�+����꫆��}��8<:b!.F=�n��Y8���?k�C�7�A!	 �  s��j;��u;[�ذQN��a&���>_�����!���?ޒe��q��V?���[π��G�ۺ��9���?�l��y�Fj��t��	�f������d��:w4SG���HP��b�b����{�������Y���EZ{H���� ���p�ͭ�^�W�5��$9;TC-c���,�r��vsxlGG�t} ����;:mm���:��g^dޮQ����r>^G丼�QY/;����\��:�qM1�Z?_�������ǯ�&�]�ֈ�׍Gv���?\ۧˏ���s*wv{�)�®|?���f�m�s��^�j[�M�ST�A�a��M�n(�2S084�'�j4��8̢TA��/w::�1~Q/A��/��/ol�&���~�����/���[�]�1X;I�e�W���Ds�>�I(��O�Eq�N�Ȯ_�\�1�e@��NO����L�B���v�ǔ��qd�uQ?~$l����w�Ȋ�����+!�(����Y{�)׵w ��ױGT9��l�ckV��vk�E�Og�b����.	Z��xi��׫��HZ.h��������5�z6 �]�.Z�=���}D؋��.ݳɊ#��9����w�v�Ȉ	ug��I�u�}Q�zڢ8wG�� r�_H��.�?��uָ/�=@Oq�$���uM��u�wſA[���JUTmR�������o��#;�l�(�9���A� K�L�g׾Xo
���@6��/�.�r\�� <�� >�� ڨ�1Ȅ�;���S|�|�<�*XCW�����俟J6��a7���,�K�S�q�'
3�;~�_�`���Q��"0TY�踢�2(J�a�C����Trʩ^~~}}m���ŀ\�۷���Sa|c/_�,��E���䣅��/��P�n<S���I�4����ੈl>��(��@k�gg�������-��  ��IDATن�N�7�%?��q\ üw'3��Y+OsGCJ>^�JE����N��I1�����.��(����yd�tR#��T��Yn]�]�����Y��ӑ#�s4�78u�j����;�N1�8��N���D��d�׉XHd�����V��<�����kAg�Q����(�NJr���,�  ��?���#�=�'-dp��c"�z�,�'f#��jV� @�8��]�-��ot������5�S�6�*�sd�`�7����8H�s�KR�`����4�)�����<0&��=����~f,�{���fA�S�}RK�ov�BɁLv
k?=E�<�&A����~z�NTDi���ňrb���Q�w�pO���<T�P��"���C0�C�$*)I�q�H�Mi:�飂��ѣh�˖<S][j�|��Ȟ�հ���X���~uc�_��m��w�3"����ow<���^?���C�9���5�h�3�� �LMN��&�=�@'2M���V�S�k��:�	RP���<,��������dA�b��(fg�{+:N��M �0��!��5e;&$�Y��/2��ST�2�l�~G��+P��i!��� �Y,�F-�8^�K�#]��謌Eq@��X�I��c݀:�<05CI���=@+T��c�Q���� ��.`곽{��޼}ko�}�O��է;��B��(׾C���O�l�=RY��P	
Pύ�X�a�Pٍ)�Su�ӋX������Z���Q=�����K��޼}g�����!�^���/?����#�Y�1c��j�S�m.�E��*T�q�؇�8��@���T]�1�u{s[ �'���(���������y�'l5�A��ةo^�F�^u�府mW���;�K�֊;��F5��O~���<F�Z� ��7{T����}$�V�@��=��(��u\!�L���-̮��}��C�Y�cٶ�N��V���~Z�l��Nʞ:?=�C�sI�����'����jA�52W-?�_�>�DP2X��g&��ND����J۪��ln��R���C�y�'�Y�J�����-�Y,ή�B5�M�}�cxPe&,�<��z��)��2�����ƃÍ���>mi���޹�mxx���#���VNr�s*�w�H�rɒ��r��=�qP��k6��1�E�+�����g�L%~ό��rew��z�R�ErQ� ��,��d�3윲U�3"�k�-K�U.3A3�P|l�^ ��c'��i���8�AF -����a�@���td'��!�=�L��Q2_���o�����8������D��(,W�t�!Ít-h3w�"B'�)b�v��H�if((g��e/)�R	#3?=~����G�����4�)z̍�'�E�G��h��aZ��h�ֳhgq'�eۗTsY��%��ϟhA�"	*���s��c{�\�����Ɲ�l�yZl��.��K��7��C�p;2��Pn��mT=����c��,P���d�_���є��|$5&;�K�JϨى�{�?s�YQcI�vrL {�B���;��B�׊�^���ih4����a�.���4*F�6��RmP�����ܸa1�3V9F����1]���Ӛ����$Rw�h���&�"%���]�Cjd	��3�U�	���#&�����d@�F�3^T
I]��Dh!۴v=��?���R4z�Z �i������ak�j`Q�9��g�M�/��G5��"2Ĳx��JBU[_-"�leR:d_#ԇB�d%M�1��&y�J�j朐�mj��s5x�xmD4�;��՘��`1R�� ��Ԅ�A���5\7�w���[����V@���r�F����s����+���1s���n�V��2� @uelFo:	I�+C��QȪw�|���A�j�V ���[N`Ȑ}|�셽�������vr��ش�*Z��Ӝ����oK�P�Yv�����{
���p��,*�.j't�b����0��{����X�RQ [u[����{\��iq2O�_i��N|v�}�V�vG�sJo�h�ߩ�?��;������EZ�������~��^�~eo_������g6k�k	rɐ�+`0�3P����� d�˾@6�
���}��|^��!�x#�
~�z9p(���ZfO:9��������Ȃx����YK���{��ǟ���^�B]sZ^�t���C�b\p!��jd\��j���^��ؖ�����uxؗ�~��٨�.����s���C��j�� ��6�sf��MA�ƴ��c��ټӎg!���@y.���� �6�^����x�!28zQ�R�P5eدN5U�w�`��U�=�Ծ{�� �S[��7�M=����iy�mͲ�Y�j�;��Ծ��c�B�d���썳T`k�2�ۇ���J��}oJ�������Cv�;f��S� �����,�����.ɼ�ٙ�,����c`�M5MȂ���`
2�G���כg���lV�*=
Y|�c�d�Vm�#�k��['���i�P�Q����E�`�X�:���X�-�#���L��2�\�(05��@�-{p��̶��^[����!�&�����ƿ�^�#1��S�V �ᭃ�ks/I!kR8h�>P&�,(�1Rh}T����(э>�P���㏅�4!������V�(��=|�s#��Ae�h�H��*�7��h�{Ñ��fl*��Ǎg�׸<Oo���;)O�C�<\�G�q��ʣH,x߹*I�H_e��B�U�)��w�� |�gO���gO�:��i�k���Q0 4��B]�t`���^-�4t���0��f�0�_�~�u���/���R�=���^_7��T{���rlկU?��,�z�@K�Գy��):�H`#��L�s�	{x,E;X���}��{䭼h�3LEW@Xo��_����4���Z�6ƀ��T��@ktJ�#����a�R�6��b�[����2�0��s��n��fT1+ȳ��S։k-���_�k��^�7�N�Q�Eu�����M{b����S049��g�4��4���l�	�j�7nX1o��}Fh�hh�4N���~�%R�.F�����{j��A)FǷ�C�9(�=��|t�u/#����.dg���)yѬK�GP*9�m�Q� �kѦ�i9�Q����7��س�-�l��D��� �bAO��qk?���~��G��o�����j|3P[��+G����V�_����k���dKe3F/���=��-6j�(�4r�/�ZFe@���T��1I�4`���]\؋o^��w��ol�wd���8�hD���ty�<zT�"�l�o�n��~��S2�ɮۄ�/�% �*g���U�7�we���8��]���2�
�lяgT?����������u�>'W}��3�K��@YzN@7@�#7�?|d����t� �!Btk�?�����۷�������d��u#��$�U�A�V���<TЏZE06�N��]/�5������h8F޹|~��"��.��?T���"�FY$��p/�?]���}x�6��>����8[+I�3C���i����,¤�|x(*��	UR�@pgŠ����^BL��պ�*�-Q���o�^O�xZ����e��Kڰ(����l�ϗQ��Q�:8fծB���e�w_ب������w��
�C��I��D�y�CR ��d����Y�{zd���Ջ�l(����Q��H~��[;+~2:=�v��k��I���e� Ɩ5��!8܋߱d��� 1�Dm�2Y�'�3��\���R�!�E�`a���� �G?k��ym�,m�$����=z���23� �ԧf҇���K�b���<{��lAӘ�ݗ��3(<kbD���c q���x�3���YF{����:[� 7���<�1yRK_��-Z�Lg4�Rd~1��Q�\��* �DOP`�NvO6֛g����j	�Y3�'�of|�ZH � a�h�B����.u���@2#A�.���P?�4�����}8��GP��߳��'|\(��(.�R˸������R��;fPc�M1?������������O�@<�A1g]@(;���=�@�A�܆j����wr���̬��.E��W%{���� CS�����tL�	�^�`�*�N��6z6`2�;�;M(e�pO�2j�c��&��)�m[�v��#ݣ�[Iݫ�S�@�M��!y��V�o����Ҟ�۳�3{r
�R�RJ��po��-�	W�\$;B�,����lS�+PE�Ӹ*�}\�c˞,�@��QƁ�Nʲ�vDp�����'i��Q>CW���H�P< ���F;(�oN�(�$�4Z ��V\�46^�,g<u��4K� +
�*�*�c�0DB���/�_���ɡ-����۳� �%
��@�=�6����/#j�'��:��?PC��k[��
-G[�Pk��E��e������L� @~��Ɗ!��.�2�Zk��YM1���j��h�V�:)Z��oD�7C[)4 l�_�ܹ� 杸bvu�	���f�2)�J��������(�n�����H��~���\�0] d/�T��9��Q��:�ܳ
��je�KI}�ާ�w.�$
����_��.��;��X�k��>��Q����lp����r_rg�.��
�.=���0}�lqf-�^������2ZWO��A��]~�{f����Z6"�Z�7�}x�����/��'ggR�G��px��#2ۆ��j&AR'P�O����]U�
g*��G�[��L�����{�}�ꢌj�>���a@
x�s͖����HA�u��������������ٟl��ت�jCb�M
�~�g�|R����/&2���拎�8Q�gB�{�0����G�vQ �}gc;���b?6�d�	�.��:|�L���l^Y*��EYH''��M(����$a��6{�N���<k���c������	�ݪ�����C�*��T���Go�|��~����_�7��ا�;[o��vdcY��bgo�q��%����m?��. \rx�2v �}R��	^�."��H���U�J���`�=y��ƒM^w��(2Y�r�ޜ��k��}��v]��Ns�;T�j٭�ǘ��T��\�bgl��@�l�^���:l��$6���d� �pQ;x���Gv~^��n�
��^�/�i�Z�r� jg�gŖ��#e_����R�I'�����u�F���"���hw����A��nC�H��~�Ζ{j���!�������#�C���l���FH�/��ŷ ��ߣ�q�c��4��m�\�F���P��dĖ�<��Szd��{�Z���Y9ǋyX+P�}C����kY �_�7A�5yV�*�&X��U�a�xŞ��b�c����Qm� ]��CG �\ � y@�$���g�|�n��3,���HQ�5���� W��������b�qG�#�A=��ݗ��=�^'�U�mP�i������`(�)`�C�&M�+��a4�Zta�	邋��^+�9�Y��7�S��]زD����� �t!%H�P
�K��7/���Ӷ%�?�*�)�Є��ф;;:��[٩�9N�IQ���i��%W̜;쮦�Q �|��7��ݹSǛ�!Y,D.����FO����	�r5�^͆E۟��z�x������P>�"gg'��s�B	 �����������C4�Y:k
�?����7yt�N���O
���5�U��LL$O���*��9������g��,L���)���8<��4:�[�ʆ+����9G\���)�Iէ�ye!D�LS6�W�cH:|���o�m�)ÊHS�\������y��=@��F�ۙE���(��Wr�a�d!��k����^a�q�A�y�|$�bT4�Dz�s O���ne{���7|]�B���R�k�Ғ��3�tP�3��4 �r�  �]P����A##mf]B6��:i	�G8�8P�F$oi��
�m�x�;�ʙ]����x[X,�i�Ǿʳ=��ٔͳ��5�g����-2�UD�� ^��� /�q�k�h�����n���a��NC���ŋ�ݷ�����|> ��2��a��{ō�u{O�h��4Mu�s�*���?��~4r��Ơ�+�(��$j����G�4�G<@P�A,��8??��ھ}��}��wv������G�m��h�t�7��j�,��!��cY�l��G��ܦy�Қ�X��$ŉ�AaFe%Y:�^]~�/W_l�2U�k]����R��G��O˽>{��]\<��rf�Q�^o��vv���$��"����,P��g��@,�A��b�����)!��_(�~���y�R����7�:�Ἱ�b�߿-��%�DP���ڑS�ۺ�T{�}�R(���S՚2���HJN�m��=j�{�5� �B>|m?������?؏?�*g�'�����ub�n�}��}D�6��3ڧ��P��g)�Q��|�6��dK���� !U�>YQ��nG�k%��� ;�T:v��͠�����\[�&�/��R(�m��WPo�vVS��|���g�i�?�	�@y{(��̠�^��3j$^\<)�����->����==	���E(D��x�J9u&�#V�(������l
���.�칽�!���;知 r������@3�1�j��Qu�u(�8Q�BvA{`������h}�I��:c�rjw���yVF�a�c��a{��,Z���A=2�^������ �h/;µ�Ju8���V�l[��A������W�ѧe�$C�~����R�{���i[����ȿ��,J1�%k��(6�� �Nf5ٴ�	�mVǄ��L�X�S�R~��ɏ�Đ�E��a����C��������J �Sm��65�� >��D��[C��a&�x���Y̉p,�.̄yr��N5YsGĿ��d-�K��S�_�0�]PΪ��e^������ʢ*���9Ⱥ[�1S���H�i�g����0�I���,��\]^���}E>�oO�<q�/��ۛ�}Yh��K��"��<�.9|
� �Mj:���?T�o��q[p�%�`n���8E�q$�1L�#���̹��kF*�����/N'8�PBm���A1���~Ǿ, �w�Y覭�l�$�s�{��w,���`�#��)?[� �q�	ZF���w΁�37�d�	��4>-�Hzì���㙙ȯ����/�J��*��|,��|��''Vف8�[f �^��%�b��	��]o�n���Cd"���ѧ�9�k����	�������E!���΄�/&ﵒz�7�2:����4PJ�B��^BF){�hf��n��=Tu{���wx��Q*��Y���"������!�� RV�����j���kN�W'o\��PڒQ���T�yis����y-��r;F��-"Ţa@��O�>�Z�y���E���@R�hc:�Z� YS�a�{�~�y��F0��X��Y���rH� �]`�ŗL����- ��/o��?����=�����h!ۜ&�W����um������s�DGI�����9�8�#r�M� �'���
��re����|I��\��9^��AIi6\���b�g����o^~[��Y���{��^DG�o���������|��֚z���`������8߷vw}e�����bs^�cγ�c(�U�_�,X�v^�:����}�f�s�@O�4Vw�{i�g��Z[/���涊��b?��F��
�����=�~�����������~��}Xwv���c� ��N`	���KT���6YB
\uކ��ƙ��i��JM�YD����1w���8-���]��Mݧ0�R#՞�az�}�a�	!�r�u��+�r�?v�>}V �{um�C�y���sz�f�O�����#���N��������;�u4���\xeGg_fG�R/3I�C�q'�bd�s�lsߓ�4fe�K��^�w�!�"�n3Jq-5A�_�͛k��A�� �}��oR�Fo�n�	8WHm���5P��)�:����9�d`V������b-� 0������z-x_X����*X��p����4%��F�T1;�b���� k��$3� ���'h�#�������ۖ�!7�YM���wam��ӄ�[���Tk��y�=?V��(7�x�r#�LV��c(f���h�T)�\�� hV�bj��:�nk���f>�|�O�\�����󨟘8us����k�����IeC�v[�2Ыby����]8��7�ɜ]�;�������Xp�#��N�e#�P��Z�(���f�@V���1���l9�#߫w�f �e'�&���n�X���5��jp���Z�h��u��f��h����o>�W�O�D�_B���z����!���P<���gei�\�(�O��3:F- �J�u��[��Rnf�ʸ���6�@E��X�8�o=32Ff���R�̞!J6-(8(HO�6��M�qlaE3��<7�����Jʟ'�i� �Pʿ��j�nȲ���]��C��f�@�F��Le&�Ff����͏smr9�T�q��b���n��m���'?��1�3�JCh<J�	n*TK}���uy
\�b�7k�"� +���<�R,��.��ll�xX���R�f��k"��O�-�5��w��`�Sf*n[��՟����qjn"hR�\�O��+��&�8#?�4ٮ��eQ�5Eۂ����6����:"�>V��(Y-y�X��1M�}��_����J��EI�OI7�w��v�G/�D_ldo�?������h�|�������
�t!��GQ�QFd�������*�f��ˎ�q���L��
4��F�G�����#���IC�f��^�H�޼���Fx;��B��qt{���>�>(%d�O����^~�{��%U�J��^��T'�Ҵ�x��l#$�;���z>=��ی���ջ���Iq���k�.Dx�7^�0e5��-$�m�2���k?+v��d,�,N�!E~@1�@blc�>��� 4���6Ω?M�ę[\ܢ	[���<���n�ݻW���/����������+�aݰ�۶o��4�����]8&PYR1�8ݖ���A������B:s�3��ZJUq��>�����_�z�o�!�ɦ����6{q]N�(��Yؕ���̓mP[�J�l��|����oL�gu�;�n�Г+�Z��u�v�{�<yʨ:�7���k8�+����8V@%���}+q�V�g�s�:�~���#���ur�;��b�p�Z�feҽH=�έg(T�p�ނM�#&!���,Lv����\;vtT5�!pr���Gl�=�[߳i-j�@ido/��К��ᒨ�۠Ə&�U=�\�k�v	���asg�q������-�fwY��j�5H��"[v�z/�;����Z��:�J�Mm��.ZQSY��F�#@�{�*�=��6�i;?s���ؔlh* S=�=<-�ypb���uMs�3:�JcQ���ls�p�gv��-J�"�}y#\�R���1�x��b97�=|"87ѓ��9i2�2�ϥ�VI�����4��FO^�B���y�mrS� j%��T;H�9��f�<�l�GU�PNQ`/p&��:- Q�Ѹc�&���� ��8\���P��Kvy����R��EF�h�<�د=..�>��_����W_9���4��6X�h.�F?�x�d�RЊ4:�rIψ�G���Ԏ���عս#3�1{(�j��?,����EcW��cn��spJ�x�*lW���lV�.EN�b���V٪{���]�n8��٫V.���z��Q��;n��F���6��k�c�=�΋�uvA?9Mʾ�B��Ǟ���C�LE�P+�F��XDfA�Uu��$WC2<yV���7�I�چ˟�4�Iƕ sT3�����tD�v-	��g��N?��H͡�Ө����V6����Wd������^�%���P>�P�[�
M*ڨ��&�ا�T�}�LgtKg��#c���S7I��dw||�y�AR� ��؍��<\�Z,�?��|��
Խ�݁����*��<�F1j�1x�U�=6e�F��ym�O�U4"t)M?�:���Y������6� ��������H$��A+S,!�����y��g{z��N���6P
`�W�X7Sp��@���'�A�O�bo5+o�h8���Q �Ӣ����eA�����w���O���[^��r��7���9�Pr_vX������o�����ٳo����%�Oza�j�y���*d����/=�����q<HN��O.s`�����Ϯ�
P��B���3
~r�3�����A���o�|�(#�IA�r蟜n��肵ip\�^��ш;�f�h���Sq��u�1�R��v������<���P��������ؿ���`}�˫��5qc^r�07R�-gh�Y��V��_.����8v8K�m`�ˠf�
L��"L�1�oD��0�xK�#8�����:�3�V�?�����uh:�` ,Z����J�=�F|f�^�:��8@	�\��с�x�ܾ��=yza�{���0���?茲���Z�ܿy��ӧ�T�E�R�s-�LB����,Đ����pD��[�@�
 g|��q �|ouĚ"��n�4@�h��L[�\��	���n��;��v�L� !j�F�;	eJ�g?/�B�$� ���@��R������݇�������7<��L��MP������?��<B ~ ���#H��B��YS|d� W4��z���� ��;P��e>�w�<c�r�+6�����>g4F�=�{�7&��!�^z�$��QB��k}LWg����?TJb�A����2�J/@�ϳo^K��%�C� 6o��*`�jp �ɡb�3	����\H�a&FC��2�+pw5�e9�/^���<��9���PP��k�+������3e_��X���>�0�c�a�T�9�䈯{$�;{�௒�J�;�7n�dx� �-��4^�"�e��r���r"���e퍵E+u|n�h0NeB��g�^�@,n�E�v�6�9�2Zy��J��G�����<~M�-�T�*(v���P�Uax`�Cs�ٗ�-P5G�C�L� s
!E/��x���NOY8�Y���H���,�D\
ih#z�F��o}q��z���a��i�W�Q�,8�Z���-G �-aT}�EW�P~(���gG�Co�="�� #eNQ�����I�Bi0��;�	IhR��m6G��=����6�pC�(�������ĔF!��O*~U�L�a�Z��&���]��֛E�(`���7��s�����+d��m����4}��.��9�����87�f��cW��E9 �xb�E"r�ό�%�ɉ�VA�lX�y���Ճ���:��.�:��юզ����-'8HӷN�͡~Zi��^O�*��P�m]?�Y��˫+6�<<:�-B�x_� ̒�zf�<�.�E����)0���:ɽ�{rꃚ=�^ x՗=�����(�����e���w:�X-)����rug?���؈�����9(t����ȑL]S&AǓ+BUpY1j�%�"J�}�[W��,�� ���� �S��A�ݚj���ho^��8�?�������=�����]�Kp��8��^G�{���<�T���:�F�f�E�7��H�qЧ��9x��4���Ζ��V9��+�Y-�K
�::~b��g�^����p^���0��6TR����@��'!`�~p��{;+?G�t��{E��B&�8F�ѢY)G�q59��8͑� :/ь]T��{������������?�'��uq|�r}��Vl�-)W�c��g�?'��e���p�@�c�e/��|b�;��J��}�����&����Wi��e��iKEǑ��%؁��s;�H���V�T5�}9���pJ�p�+Ky߅��j�쐪w'T���o���}���vq~��+΄g��7�*& )l����'v\ V�?�܃���g�aA0[������O)�t�g�̉m� у�9�sS�4��˕�@�zݝi����8��{���H�#��H_N���'`]gʏ�Ǔ����h�gƮ��n�����@�v� ���nm//��\�~��2.{���<�!���|ֆ���
i�d�X�~[�O�\����h���Z)k9u��!��Z)i`0o��6�۰���3*g�강�Av|t�^�Nv+K lo��]����ŏ�_�Tv��i��Ɍg����%	�%����q��F�y'��H��zL������@ ꛏ�����p���q�o�-R@k_��0i�ɕ��Y>)U��+�5x��M�8W�߹�A1��1ƚ�G�<{��}~����(S�bW��o�};:Q��5�r�E.����Drw\Тs��若�U�b�u5.8��s���E�,F��4)�!j��":�>����i�M���p�7���|L�Y
GؿFS��'m=M=�����k-�HAm&:z�q�Ɵ����0m��wA{�(��{�N8*���p�6;�25ۈϼbi���"�cl6�w8��#�B�ϬR�`��;�u��r�&���͆Y�q[^W@W�{ftɉ�*C5-0DH-�Cmy�y5s�0��0ʱ̤bk]0k7�� )�;�4\�����׸�H㙬E�H),���>�P����H��RX�����7	�ǘ2ۋf�Y]٥:����6lnl��6�P���� +S��uY��t��F�X�ѯ"�-)=3ŉ��4d�!L� )|��w�:� e���lj�Z��y�*43}��ɹ&/���d��Y6z�/�3՛l������ ��a�b�=Hn�54��1�� �f[�D�)�'r�O�>+��;(�����,E�ōOR}q{#�vs�����L@S�����ÆEml��̻���6r�K�9VtD�^6�5$^S�!y��o>�C�}��������3hV��LC��*��%�m�w�k�0*��+��J�Ͱ�>�{(���z��޽��~����׿�����E8P|��7��SمU��'�v~񼀲',��el)UŤ�Up��}|��������C���c�s�C���T_�X�aX���g�w�����HP��5�r�:�ץzeϾ������=���>�K{{���\p��,u:]7����Ϙ4W���صZ�8_ ���ӥ�y��~����ǟ�~���?�}t_�jf����17�}>�u�d�W �����a�e۹2���̨�-_삄(��;�6��̐E� Y���N����G �WML�~��m��RM�ӓ�᝗�ӳ{R�����T�>+ ��Bz���Ӹ�
B�V"W)�̇��z���?�\���#|���+�7D5�>`�{�e��랳�_0��)��NڶR�0h�)�����׉�H~����ħ��������"�S�Yr0��xQq�6 ��/7��/�����I�m]|����aC��l`� ���Yʆ�U�(���!��<Q��5).��!���r�O����b��@�fV(M߫�<�����x�M�PA� ���b^�Z��3a��TV\�a�s�"L��DX�51/�Pm_��S�!�E�1?��ኴB=�&{��?�K��G����1�鹝���"`����K�\T�h�1#5�^Wگ'2s>w� ��h�<�G�W�~m߳�ǯ����"U�3�2���ģ�,JԼ��su�jݔ#Su`�: �&�B���[��*����gԷ�̨����p���L�YM �۝g����5E��ʯA����`HS49��>��yf0(M�W�e��j��	�ՕUu9S���Ǵ���N�Q��Z�X�B��L�Q���������],����yF��w�X�׈%��;.���ž2�~�2���D�1��d���l Le���{v��
o�a�,xآ��ݶ*��,��e�	b�u*`F�fl���PS�Ց��F/���؋󝼁7�ư�ik�����D�@-����pȷ�Ln��8�~%���'VF40"8�	U��1V�@+�}&7��6�T�"�;d�����Wř"�Bam_�u��8#��AԘ%:/u}����N�! ��Q��t��|��eߟ���;Ags����~�Cc�s�yF7�P��<�~'��82@�=���Ɏ8=��a�=h�9<���"�
��������MY_ʓj���E�*~�J;�c��G���L�s��〞�d����6�B�@�.�����%����XעL��,6%��WH�\���`��vrp���o�۳�OHQb�)f�4�����+�rq�*і��Ziͥx���&��QL.�`O�n3<0{w�,��`�{��_�~����6d'{
��߄b�ԥ:�I@������?6	]�N����8��&���Q�]���)����鰯t�dU9ϼ�)��`���Ξ�����O���Y�fe�7p_ýB;d�������*3�%NR$վ��{�Gv�9���c*�l�n��@j;������um&S�������Njgpb��v��K���/o�ܽ�ׯ������>�xC=5����iOG'z�,r���?��eAܱw"�q�,��7ʆ��Qk�=�Deт�ڭ׃�pףb}�4k�����´5�jf���1ih��A���QU��J �2���/�O��=,��O�(���/YWEb���'�UȰ�Ai�r��q�,$��%e>WS�f�n�%Q����+��;���ٲ�t0R�ވ����ΠP�@�fB|,g��F`3z͜�ɳ߫ڱ�j{�x3���f��P>{��<�U�/�������1�9�8���`nG��H �5��5���$;WmI���M��T|aw���]�ud��*clc_`t�DI~�������$�u�z���p�9���O�F��l*g�����P�M�P;��5QW�:�����G_s���5�q���L�K-ٓ�I <��!+Č�d�A�3^�'�P���,���S�ɡ�=�≁*�����;��m��yf���ĭ���*�E�����^DLn��_�"��h	d-���� ��Pka����߹�fT#���K��y��N4::�m[3@�P�����d�o"�c�m�N����/G�um��?���u������B�� h�G���jYq�9���=�*�Z�&�=�	�
:1��참��r�J�Qŵ�����k���h�S�7%R��'O���Ϧ8o*�[��-�0�_�����v ��E�;8x��� 6�8�ᱫL%��"�թ$Q�'*I9X�"[nJ`��a�4��_� �]½��΢J�8�c�G���<F70�	��I>�Ѡ6ꦘ�tǚ�-���i����P��Y'tyw���E��\)��'��ِ���Î� U���nK�,8C�P�aO�\��=�JFm���BL#ϝS�s�SM���qGd
��,V -��jъTh�(�K�I%j��)#A�Y&��9��,9 ��g�ٽ��.�� KR��K�&���9�Ƴ���SDu�%�*E`f�oEz�X���Lt�Q4�e�Q[�5�@�
-	��Fs��pp�.�0@h�ۇ5)^l�q��8l꒠�6�hт6�ý�ݖzPI�dz����}k|����e�������T��j�7��f��o(�rx���bSx�X�(a��YJy�=���yx�h�))�p45 ��,πTg������4�z�ǹP1s���2(۰`�j�����N��~S�:��@�|C�1���A]��T�|�%vU@���5A���s	ʆ���s|e3�����S�`�-� ���Zn�!@F�wo?T}|_�_���e�a�٢�Y8���o���tSY��Z!Fi	�:��[���5��Nٳ��=�.�b����f�ևl�r�v��ӨT����(X#?G�!;��O��4������q1���j�y�;��-����˿������_���gvv|jG�9�X����i�)` 
3k�������5p<�P�s@��aK�iO^�9_�\�k9`c���W���l��hN<����M���R��.��J�yP~Lu<8�$J�A�l5�� j��,�p
��2�4`K)�R������r/O/���tL��%����ؗ
�����߉��I���	�6�Ԥ���8��X�$E�ӊmn � @� �Jo����k��)�^�Ǡ\�����%�cH�o�,A�Ze1��QC���gw
�o�?�T�i�P�bL,ȳs��fY�G��>�TT�,{ے��A�Bf�O!��,�}��u�:����`���b�(QR�`��.���k��v>J�~�rO�4�����&�Ī���ۚ�x�*Ț��X����	�6�qg~�I����Z��y���(w��G�ٍ$���N�"7����G�(^�j�'>�8@_<a��{{V�ItmU7�+�ő7�@���Y�M��������W�{��e�r5��N��`�D��9�6շ�oL��\��yt�Ύ�Yz�f�|& ah:���%�1����/SG�V�0	8�v�T�~Ÿ�3���� ᣎF���д��g�:+q�� ��R)OP��T���V��K.A�0X��p���*/��Q�''���
T���f����'���04<nz?��f��"�U#@F�#+c�@>Ei��C�kŧ&$tE/�� �=n�g/,�Υp%��u]Q>����|%����mևFz�e.��m��V����5{�")]�D�� 壝�(������j�0]�����y^3����Ʀg�4�S�m̳Ϫ��p���-%�ю��E�vtH�ǜ����� q��L�I�^��Uv��̃0��k
�4B�N��p��2��8��-�������6���Ͽ����:�{���Ğ��z�� 
��0��:�=N_�lyԐ�/����hf�p�����&�[_*��/�Q��޽�Ѯ�|��D���#4B_��N�z���ꢰ���Dߙ���N���j&��I��!�S���i���z|t��3��x���<����Xk&;��"8�h�
[z�^IG\gh�=xsz�=��м޺�c��7%�c$x��8fF[�������iI><,`� -d����ʳ��={iU[��P��z9�]]})���]޽�X��'���l���[A�t���w0w��
�nT#v4�D��n9�O�/`��� ��[�xϴ&M���:.�oT��3�M���	���F�~x��"��0r(�|�����"KȬ�܁��9��Θ�������_���jO���>d����a���Ng9 ֧O����L|b]"|��͈7N�.{xkg �tؑ�</{d��,��u[ j�;�9|��-w��k+����2W@3�b-A�bf����Z�2����?��i���H晬�2 �{���8f����s�Job&2|`S���7b�:,�ϙV��5fQ��y�F"l ʴ��a�t �j� �Ã2�`[��_��G,�+�lPɷIdX�q?��g�[�a_3���P�T833]D�������|�v�~������2�f^��k�Z����/�6|�<L�5���Q'�惺k�k���dej��`C��P4?�i����B�,սl�it7�]X[g�������v6J�`����������$s�U�4�ޙͯګs��x&J�w���S-/֋�,558�''gvtxB:��z�Ft�(�׶�t�;pACG!�N ";��n�{����C����)4��)�/ X��죧�)j��u���
QV�n��uy��P�*5#�@�T+�$Y[d^Ɩ�9�;}K~��1� �0�j�m���f.m��M���E�������:[oS�(�?#�����f��4�i\���bT��Mq`���s�}��~N�JJ)�a��˞�2w^�Q���&�I�*th���)�~��@ϽÅ�;$
j #�d�Iz��=��qG�wXct�x�9
�q�k���c�n�1ͨ�6�To$�M�X4�ふ-�8mq$�ŸGr5�r/QH`;x��8�m��y@�el�X�F��o�Q3D�
�)�.��@�k��}�#i�I��Y|g�<��$ygsQ����yW�몼�e��5�},�Δ�(�����#3�N�@d<�k�����|���"(���>u.+c �CH�')!+P��rkAM`sb����%�A�d�W�}FʃM�mr�������{�P$���h��E��]#j)֍2�[�N#r:�t���)B�@H�+/R���؇RDE���u�M�Y$�ث��N e��s�UC2���4D���M��<�pP0���p_W��"1P0r��Xd:�J8��]Yð��sgc(Ԧ�x{��|�ܶ#Z <)o��쉥-�!*�gjv�1�z%+?��M�i�ç�L�&�$�6��k���`W�?������W��û���tV���u<SD����W�����{������vx|dmqp��kWIHS hP���i!G+@~�lo����<�C��qFUK�c��z鷲�؛m�g�~�h6@�����L6.�+�w�����)�ݙ@�AЙ+���{)��<����N����~�R��g�у�c�,�i�QC��gP
F-
8�6m���<�u���WP��. �mq�/�㾶����e���=����swU�DG���)�z�F�b�+ KH��r衈���[9oQ9:������1.��50|��
����΄L����6z\C-6��zq�bV#h��=3��W�K��?}�G����_��_�/�}4��l� ��~|Y�^�Čӫ_~����_�B�y��s��i�e^���X�/'|O���e��ľ����-������_��>��/�mݣ��������X�>_�'k(�Ul�e��x���{ C���8�
d��wY�m��}Y��wf�oD�\0]�k��jc���5�c�L��澜�T	\�ն��E�r��?��{*���������ɳZ)���/�v�J`�����>9�?~��}��;9�gF���Ž�D���1��?�����W�P矇��/e�������|s�&�8,���?{N�VWE� z�%0~����y�Ɔ�7�u�)�`o�g�H�t��H�8����5�
�U�9yi�����l��TDn(�#Ptq�&p�J�o���z�%o&?l&( C�� �r�/�m��2�+x��b=�c~[�9��]"]���`}]1�\�\۪�R����p0e�,��&l�Tc�*CA���Ju�l�����,�I= 4�9yQ*_�
��������j�q�@��T�6k\:�u�Ɩ���!���999��ϟ�_����_�b/�yIP��.����G%�=����4�0���|�y��f�Y����-�T��0 �ׁ�G��f8�)���/�Lq��C:?�g�u5�R�q������şe��@���A���u1 ����O$Yxw`���+�wV9*	j�-�U1$�\ۺ
��!D��Z�<j�j�EˢLd�vu-��t!�ov��'PW����Ŧ��  c��AdH���C�;PcDE������#��#�/W���jc�ē��\�qǆa�*�ߌ�S��2��LX5�\0`�eM���/��3�8�kb�N�jP�,Y�9(����i<"7��"��+˙�����$���[��\/�8 � ����,{�T��;i��{�l�Hn��#��Q���p��Vi��@�+E�B�^�er�m]J6E�#��˲�g/V��ֵ��i��h�v�h"B�&�h`�U�-L.��ȱ#@��WF=�jyf�T^诋ڜINI� et�.��E���+����q�Ü�\Ch@��4��{������]g������`A=�v��y�N��̺L�<F/�����m��ތ�����i�,�q$h�Y����.��p�����+#��Cr@� ؍~g�y���j���I`F8ْ]���2�p�CMM�*�O%8�T����v[����O�/��Ц��oُ�EH�gr�Q�7�R"U����'�&�fV�	b��A��y1��dfC�s���e���{Eb�A���lq-fRN�H�X����Ѥ��V�0�m(PR�������P�:��^�wd"�k%�����{-�FJ�ӮnKP��#���1�����޾�T��{{��ܻh>>���y]�k��z	���8t��8%��Lte�x�

�B�9w���jy2 �U�w�uQ�q{7���R��;1)j�3ұ����Ei��	�r=D�=��`�q�W��RZF�z������W���c�۾�ց����v��RػL? �Jp��������}���g����,���|����7o4H���+�XKW%����u	���������c���?�z�>�^�	j�D�~��SU��^_�=�����]�g��Ӥv"����r�=����eѪѿ�:;�_lC)�i\�W���/6�\�JR�f���3�!@wVl�l�˚�@f~�9���{�:���H�����k��_�����������r�.������H�����ÇO��:��/��}kߖ$��b�Y[L� z�t{g?�}g?�Xl^�;�k_�$�/��7�|���:O�3�紐7������?������'��M�4�B�$�}m+FG"Lj���_�<2�Isu������-ڒ������Ka/#���x�á�F��49 ��o��شsE��m�{�T�4t����b{p�A{��-i)T�ԱQ��ʰ�v|y^��% ��"I�}>aq�ې��KX�laZ�v��-�T/`k����b�VN%�d�
ڏV�̧J��S<�qJz��K���+���#_�J�_|���������_�_��w���"l0��E��6��M��AG�B�Hfe#����r��p�p�^�����?�9����ǫ*��J5�lK~36�z� hpx(�]Y�w%�z�duR�3(ں,o���/ɔ��-���f����L5�a�|>D���:�#ɂ������b��i(�4J�'�sW����]H%J�M�|ù���,��(F��ࡥ�oKQ*[�� �}���l�����ɦz!&&W�0(�5�e�l1�t������lt��[`Y�ާ$'��'h��D�7�"��}VhOB�"ј"��K�Rxc���#�T��T��T�������)n��+���>��@z�:A��.k�Qm̚�1N���P'UN�c�&���Ƨ�!kMN�VlO� I0B�0�9Y�g�Jr͡�/��r�<oq�ϩ�tYlӹ�!���;!�*~����,���4���Jn���(�A��=�f5%84��ա���*�Qoz%Ul8/��������ݝ=�o�����7o^Q:���Y�oM�4�ٳ��x>��G�Ul����={�v�3��g�"8����G;��:�J0���x���9�*��hsK�<�_2��J�WM�"c�|�ƩtP�dc�t¡��x�����5Z\�S���C!�x]�_T@��tp��xo??�H�Q�s����FT%�W)OVXi.w��YQ�dW|��:+��]R?���rl��|��;��T��a{���������چ�\sЌ�h��u8ND�Մ����X�4�9�u# �dP{�{��$��������؂���=8�֫]�@0R��\W={Vz&ZMV���x6ח��$�>�*z1꼾��9hQo C#q?���{���z�#���J���G�0x�J���nP�92��n��ܿ{��>~�H���{ݝ�Za�Ƹ��)p���o�|,����v�1��K<�;;C2T�/^ٳ��v����vT�#=4��֒�bh^Z/N���u�S��[XY�!�Cߪ�ۑ`;ŗƣ��$���w��q�8�m��*��P���>���W/�7�YiZ�6���wϟ]��gWv}ya��������A��OY{�:��U9���6�}�勒\������U��]����)Ƒ����$Z_;�H:�q,���/���,�5N�P��L���>}�a�XCW%�yU��/���./.w�����]�8/I�{��Y>���w��?����'uqX�`��я֦�WK����;��N!�lF��۴�C0��D�)�}�($�.�k�y�8޷o��7��yسH�[KD+�N�b����R���s ��{��@��Ɏ�ۮRk�֘��b����4�3,��`��6
"�o�������}�f�}��.�W�����S���|�������Sy���H��4�"��$KA������9���,�����7����b���/�ׯ��}1g���ǽ���(�I_��d�}ˀo�7��-Yܜ�w�]��}�ga�;�%�Y��MM|g,"Ӭ�L��*�"�fd�P�@�{���=ޕ �|%eT�:"m�kh��E��
��Sr������5�g��S�Z�w3H�����bMҥ�	 ϵe|J��BAɡt�l��J�qNךO�����B��s��F�@G��|�r�ðRo�䌃3s��5�|r/S���U�{��c����!):<�A=Y֌$�i����g�y:_�u�{4Ҋ�vZ�b�ŔlL� �5<ȱ�NX��fx*�-i��A��dsY��ɑd�5Fw�
�OU�b��bo|�W�u>ߍ��5�A��4,����R}/�������CT�8́-k
켴/f��ǧ�i:�eqXd�]ƹ�z�y�}�]Ea�T�1N�i>�H���:�=�A?�~�%`�H;�-$��:��{��XPC�u��cB����w��!邤��W/��Kя�.�Tv��'�A�i3)�SS�5Ռ��%y�Ǉ�Tݕ��m�Iw�yϾ�4jt ���V�K���8��4W�؋PC�K�U�aw���JфQsΚ�������s��׸/=0��ќ����Y;4fKJ `�c�T�dr@�\�i�7��]/;��_x������\<+B��pYw=z�=�*��k��ɲ#�J�E�)+�U��Ц:���D_ktV�����GOZ�7\�Wk��-����6��Ȓ�F���@{�@������A:�Up{X�[bS�С'�I�Z����6��k�x+�Q˄2ư�u���&Ő��I l�3�Aa��z����ުL�z�!�w�wD�on>����E���#}<�p*gb' �.o�+	��@vW���KVw��v�
<@"P� R_]�����Tyn�������c&�<QP#C§�m�,#������IJ���d�R�L��+))���b$LĀ�����J��$�_}�I�*G���/�__R.�͛�%Ayn7��m���`�1{<!�y}	�3���S_b϶��g��/�����}��m�D����ˋ�6�UI����kG=V���ϻ�|�D���E�����$`���o���Q��rm�7�א))<R�<���y~a�O��m��
�7�e��㶘̂F�f׫K�'�W��FL��:/m�����Q����m;�5�84ۤ(b�Ҋ��Ǐ�X5������VG�X��(rM��9J���� �"]�q�B]�w�ӬT=�<���K?�C�������#�7�sh��U���L���桮��
D�r��*,,)���ԓg�͒��#XL6�!4L+)����t����п��_�����d_�1�����x��}R+6���4������)��c,��j`���O� �����\t�����E
�k`Y���kN�*͟�OQ#�~Du&�K�����D�v;p�rm��d!��m�H����eeu?��D H����+�m�6Tf��V��<S�sZ %��GU<瓳��|E(�/D�B�sE����39�Mg1�[����'JC(�H����朐��_x�R°9��ۙ��^��t�71Q�&�xjR}�=Iф-it6Kz��tU-QNL��Zx�Y=QّB"9���/��+�2���#��+w�`��BNZ��@�Z��i�_�� �"�m�xN��õ.�tnѐ������.�?
Z�`�ڭړΫI���1UE�yV\�̉��7>��f����y�z2|j$Yp��o����a(�ׯ���A�:N�>j�H�#��]F��2­'YN�׊����g�6h�N�=����Ɗ0�J<�@%��._Q� h�kW6xmj{j�h�)u}���?���%�z����7�_���H��Y�Pו��H	D�d��2؛��(�rmQ��>(�BE�?l�O�kr�j}ԀW2�\��nNJU2�٫�LS����s�>`�9Yc3P�Te֟�?������(��"b����_�@ ��m��
{Y�
����>�h���T�ڋD�Bэ��HZA.��5�L�b@b|�~̬�`���T~�{���v(�ck�>>�$�h�]S��Fc�	�0�\K�#�q�s� �*X�h����v�R�&�v̶BE	<D=�VZP�.	����SV�ň �?�gE_����ږ ~`�T���^��#�\����Y��Ľ��.��zH�7��v[���N	m��QF�LP��l=<>h<Nε�3����=-�+@ԡ,�T�D1�&pw�=�*�/����|��[d�Y��'E"�J��;�F_6y5�ڤ'��, ����FI���\��tɪv�E����#�1�d�X�
)��.z���k?�;�!�)��Y��T���l�1�M����uc�^���zUl����"s�*���!A/�����|~��K{��\�؃��R�e�F)��n�9�4���6�]�6�ݞ�k�m��V��)R���m���b�^������5�}�w1�a�S�m8���ʸC���>��E�=��Z�͐��WVa����\��	�
P�N�<*�����G�X�wk�)�r�����>II�wޫ�A�X�>�Z��sa����/����9U��磏s��q?�D?��oh*�{���� \�2���5�����
��2�y	t-����s�C��>.���$�A���e���h�E�5�j&��P'�^���H]K9�1�}H~���H�>�gi�} ���`��AJ���P-�Ct|��hr�����1�ƹ�"s�`>��ԇ�)�I>!=IJD�.�
�.$YؼX Hv(���/͎.�f�~\9����MMx�3}BYO�#Z�Zo@�3���$h�J����bO7�SH0h�m����U0�n`��5�HT�t�CI��[p�18�H�D�UU!^�fE�LЏP-���P:����E��<��_�P�V�{�]͋���9%��	CrNl�7������p��d��ڌ���`Adk>(�3�����b���_~.��e��b��@�iE�-��*8�5�Uh��II�Bռv����r(?�4˾G�h���«�@��xߕLBhr4C�o�ᗷlF&-�)'U�L�"L\K:9rGtN3��3�r��ƚ�ӨX��s�t!ҳ\(��9�uN]Zu�����b�ڗ���e��݇{���(��uI�^�xn��v�H8�2���a_��VL�@B�$*0@��#��B�P���8�!�q��1��C?FseN��Α��L��=lg�����'&%fD��%Y�_
_pʎX�>�5���Ҹ��f�a����UU<�T��TJ�,@v|�^�́}r`�D��>�V}�j�l2�NW�1o�=�tj��>�<�������̞�+V�O9�*����K��L	�9��[�b�,�)��sg�)H�|�>�wo��j{:��G����5 ��T9k{���[y�s%I�f	��:�{�@Q<<�
ź�a���j.?[w>ǭe�	���n�$���S�I�@���J}OA�?���Z�
�'�g�扉��~�k�i��]��������}��r�@�+Yn��f��XE�ZIG_��>� `F��S�ɜ}d�	��7Jtɞɲ!�-e� \	�X�b`�D���B�:��b�6牽V�le"�����-jB�J�rϲ��s�b��4�zT�M�jg��U9tT��0w���"�5(  ��j�!�ױ��7�������j��+,���S���d��+=�$�J#j�T�������3��H��,c`�Ѫj��(=��-��<��Lʑ �G�⌒�˫�
<D�5:%�w5���Ƚ,�}�j����
�b�x��q�+ioT�?�ǦS��̌��K�7V�sL�x���s�Z���m�N(b��|rU�0r���w
X�x�p#�����z�ǅ�t�hJ[-�c�AA)���WvU.>�$4z
z ����R�}/���lL�	�E9s�8��0��h�����k���=��X�~�Ͼ�<8e~A��b���ԡX'�F��͘۩�ß�zuB���fBӱ���D�}���^����㠜.��Cg;:����͝/@cu������Z�gϐ^��CRw�2w	��s#,�m�Q��e��v�`@�ٓ)yo��pJW�2��d.�*���X���}�0��dMD<[�5� U�5�H�t�f�%_�3�1/7'w���/=[�l�i���z�z"ae�A}-Yi�wSe���Rg��d�v&4�O�z*���<�⽈M�C�Q ST�~nAk���L�"���Y�!�3���y˜|� K�Y*\N��`A������E?�^��.�$��>$7�ϘYk�{O_׊c͞ǇGr�� c�g}F�X�N����������S:ۂ�?����3Xq��5�1�a�z&1&tTVJ��|(s��V��xzI5��z�dw��%���w�?���+��Ϯ�)7�^	<Wp�P�$̂�u�Y��d��(�9��3��Ȳ;|%X�A�#N<�ʺƓ�CP�ܹ�+��E��Չ���g!j��-��{z�[Lh�,���� ����A�V{cs�ոOȩ��x�.��P	���4w�4L�͞s�bhy[�ѱܮ}ɒ����ۻ����h�nvv���Cy��%ۖ���!�٫�Q�G����RP���ʮ�f�����ӫoʴXI� �lu3"`�U����@���1&��S��9`��E�DET-�9	�
ɡ����,��8yTQQ�0���j-Zo?���ݶ<wd� G��b��*T�"�V�7Uf(ZquI�ľm��zvZ�����p�*hxҎ�����R����}�޶O�o��#B6�i}-�5�k ~[���I�@�fԟ3V�(9�"�#<��8��"y
5Į�q$\S�����z0�֠>[�9����P�u�1)H^�}\� (sV��Y[���)���y�<A̵���/�������/������ߙ(��=� p�w���=��W%�{f�e����nZn��ٞ =_��|����+WWW��w��{ZI�a�ۻ���������m���ߗc+ɋ!>�t �$HJ�'dɩ�c��dM����|����yr�����6��V�2V��_�?��:<<{P̙�
Q�f0^�4��3���Bܿ�t��ڬ�[�B��?8S$D��_�����[�K&I-x�I�o#�YwCpJr'o9�R{�R5�~��V8�&��>_ W�i4ohH��Y�䡨*P������>TsY���+��/�9X�5P�,�~����'{zP���
�W�7A�o���N/j$��iy�e�#����u���L�8r�C��'@i��Wj�1#t�V�ߍ[��P�Qu η	5�ƃO�ZG�(�L	�+�h`��F�4�U�Pjik#=&U��Wl���᰹):QS��%��9jC��Z�Z�D{UCyWD�h�VJ�hnJ�y��(�	�+�h����//�����P�Lp�G4pA�A]��4xڶۡ�%�z *qdU+�Jd}�;�
��"�r�¸���m����s��i�NE�9-s���ρz��8Eo�S��!�-��H����UP$i�0�@��a�j�g����3{�d���4��O0�F��H�-�S�P�؋$a˚�^���P��I�cA_0��Y���h!���q��vH�v���+�[6�f{��G�1����9Ӹ,G�ݨ���DЁ�\t鳯9���&:P�(v�3dt]�9!�[���go��ԩsu�_�9o^���>9}������>���y_C��LI�����A�*��-� �Z}f6U�T��4г�9+��Dob)0��J��4�=Q�G��"xA�o����3��tN�j_�_�%������(� [x{�?_&^��c��M΍���[�;PUܕ7WB����i�i�@��$�$��+��#f�T���T,��=�@��ng77�om��P�$+�#��N�Ց����=�{Zl�ٯZ1%x�`���o��跈S�Yp$|8�5��ht*�D��p=�B��
��6���.������/��";�1ɴt�M����Ԥ8�!���J�P��q$�G�E!�����ݸ����X� u����'�*�	V<@��]��Jlt~>̓W�(P(�����ފ�LG�X���޽[����[̘�S�I�.��w<C�Cٮ�~I+���#�/Oζ*�	�G���XU����uwJLuL��J#S:��+��P����F&��䊩
Z>�xQ'ˇ�?�-9��<<���=�E��5��V����_ �;�R�����vG%?>�?���?��ٺě�DEk�I�$��a@��|��ۛ{�m�ނ��-]�e9֎�,����@E�ۻ{����ǭ��!|���˲W�{��k���=|�no���7������?��?�$�w��v׫rB+-Y��·��iܺ��R�%�p#ɚ�S��>�Q� (�����qLӸ]#� kP��h�'1���T-�q����h�x.Q}ӚW� �	��1�r�4���ȿ�"BYT���k9��m�X��&��˂B��ndꖨ�\����ճgvqy�����A��0B[�c�M�9b׆"�J��0"R:�_�~���_�5)��&O+%h����w��7���}������gW��7��˒h�kbIv��ټ@%��5�u�\V/��;�!w��������S_;����e)�iF��8.,����!��� 1�f�)� PuASn�e�ת���+�(�O$mT)�B��[+��|@06h�1T��6$���^jQT�����uħJQ����T/���y.u#e��ͅ=�z�����hI�@3X�"!U6�u(���:�}:��į=�k�˨�Ugp���,ɇ�Q�B���N��m=��O,M�=
�͊}�W1�Z�]t"źNf��
Q\��� ��0���:�����MQY$w�T�^�r_���E��<����QF�ؤ�� m��"�P�r�J$Zu��!l�T�=���	U�^A�b"�W�B�_�����
\asb�%��:
�6���{�t���#�	�T6�M�쪊S�+�SՅS��X�ð�� ]��0)�c�'��T)��@#S�y�O�AI���@��e	����Y�ݕ�sa�7o�G�P08�$YϮ6%x\��kE��n$��ʜ�U�����7I ��q��������|�^��,!�f���X9� �CD��0�����z��U���G "ڬ��γMX1B�E�ۚu�P�n�����4L�E �h�sZ��R$�#�Jl,��9���@�iߖ �g@x��+�Uo�e��Ŧ��UyO���=������Gv�h������vk%WY`��e��w ��ze���k@�5&Y��O+���3�d/G8�u��Ril�_��V��XM����&�M���A&W�X�Nր.�����,�l=�>/6i���G&X��F"L��	��&���&D]d�R�>+�������n+��۫�J
l�{�ۧ���w;���M� �t]4��}��x���/�uM���A�J��b>R�+��
VL��	�6�M�{}X%��wicG���*��|��E�PH���� ���̌]����'{�ᓽ�xc7���t�̭��+Qܚ�.����I����h�����S<g�Գ+ Kڬ;(?��`?���=����oH�~���cI꾼}a�g��r���P�+�����������ĳ_~Yb�{�VԾԉ��������?�?��`����)&���6J�{�+DŃ
����+�!ƍ�����3��er ��6���8�$9ɋ�!�;���LiĞ�Z��r$p9���N��)����G��1�hG�5��-cV�\���A�z) e�"�Il3W�'p��������~ޢ�s=E���L��������(�pv�U�����rT���G�lc1u(4*h�~���
^���/8���S6s6d~���n�����%��#�_��[.�c�K�]��j�h�Ŝ�$2Y;͛~&0����S,��B��N�s��w�w?��{_�M:>� ��Bua Q����#�.��uQ�Ҝ�\�sسӪQvIT�p ����n\�K����A�A�����S�
�}OZ_vIqI��N���<b�IE�jUI,����-�캬���8��J�s����s���i���H��f��%�������<Hb��̫<�s5�+�
����J��ɋE�iH���P���h�W����C5�n�iei�~?M���G���:���ߴ��_�ڞ,5���\�s�&ҫ���c
�>w��狅PG�>M};Ic�=���X�Ó���Q���Tq���q)Ho��HaЇ��;w��]?{a�%�����'��k`�'��6�<�{�u��d��Y��b�;�X�H�%0pF��!�Bꝑ�o�A$�m�]��g�!!E�*?�U�͑�[{ڨ�L��׷/_W�*tOg]�%0�q�.ig�$�bn����ޣ�����Z?F���1��2&����F��$4�J1~���1p��[;y��Λŝ���:�l�%h��?��p{_�TT�6?�l�-~��^��P��TY �=-��(��W�@�B�� 0�w���#a��Y�B����!�P�ê���=@D	���
V� ��l� a;2�RҤ$+�G*ub0�N�]�sU-S��0z��4W2�]��B�D
a+Y�5���H`���ֳG�ߟ ���_�k�N�
T�K:�|�T��!�5\P�Ӽ"�IAՄ�U$س��8�b�0���"�����C�{̞����zx�� h��|��0V0[J��c�W��{L�u���}�_�5�����@�G^O�����#���N3¢�"�$T���˅$uɽ�#�ڴl3��&_ۤ%�}a����J���k3is�`o"��� ���h01Xp Գ�7w��ۏ���O�⪵��{�QICRÙn�>���ǒԜ��� �&$�It<�X��Yqm���׿����my�g��9��LRߗ�}_�������P����߽/��'{��3%Y�Σr�
ֻ����{����7o^ٷ���^�|M|d���n��{��},���}Y3�;&�+��2tS+є�ḡْ��j����q]��p����§�%Ks�t��F�W��Պ}o4>֧��Eg9�+O��uJJ�7��c�0y_�>���A	�^�{
)2���*-������z��&�bv��	-*k�]���xѦ�t1niY�\�uY�kf�O(��ް��UD7V����E��ɛ��l4�[=LD0!�
�����ꬼ��]]^��.��a�`���-�H�����_�uy~,��|���_Ѹz�f3�/dGw1|�rzG��f!0��r�����'=���*�����܉z���R����8�&M�;5tͪ$)�D(�i���h1��ԋӤ^T$8
����M�ͦ\����bHR	Q�z������ ���V0X�ZJb#�>_��'HTdbeR�������_O�=���I��\0"��b��3	���ԛu&�[@�ҕuF����R�s���ٮ80��^\��W/^���35�&%ssoU�xE+��$�X��}��������n��+��P���k�4��#�A�^X@��gս(����Y	(פR��@JCM;���^���fN��2�I皽�j����3��=���Ҟ@�(褔D�X�v"��M�Ӹ���c&T�Pm)Ze�p�"�z=���HZkge��=wA��k3�Ř����}(���m����@�1`,ǋ`ώz�5f�A�򿛖_��Ć�}�h��>�����bn�s=F�E5��؏�6]��J�P��2g�I�kO���?�_~i/0+���Z/�3JgO��Ӯ6`���g�q�7��5�JP�5Q��OgYh�D�3KN�����<�E�6���.d��'��e5�s�U��:���e�
R�
LI= &�Ȭ�#�#�m	��&��I'{�<ۛ��Oӎ��5P�h�o�O���~]8�+j�IK{�=ĹE#P̑ 	@���@�e�a�
����Sqp�O�v���j#����m�nۦ촥e��;�-ؽt����4�u&_�r+$���ԦM
���|���k��Gp���=�D	m˪*�fR9�_E����@���n�a�xKd�@�uThͰ�����C���cI��%��m��(l�S���rm���	�ֲB�*w���T.�qz ���56���8U��F���+���� �6�J���z;�?
���o�U[��;/��Y����������ǚD�؏>�8K4�TpM]���L�ő{䘕�I9�qPE��MY�w�Ͽ��r,��������z���C�k���'Q܏S�G�>E�MJn�}|���������I�g�]�Y�Cyi7ڍ]<S�cT1��V��%�9�MM�G�L���A��35o*Qp�(T��,D����Ѥ�fC�3�aC����;�h bX���mGUC�;^�HYGO�5����'{�߾����د������3���v?ڧےh����ͧ[�eגh���,�{�-c@��A ��p��?�Ὕ�[��9*�w%�ٕ��2��y�>�����ݑ�3bVK�I@m+6��� ��'�H����o��h�JC��l��)rq'���xƊ?�Pq13Qe%���Ϛ�F��W��q��D������C˭�p�(ێUjީ�� ������%��}��\�{� "Q̾��ڷ�H̱:?�L���`^�yc�roY�4�9,�h�J��fu��(�4ξ����%�d��ӳ�.U�M�9��0x[��8�r����Pދ��9x��|�x�{�t�&[�hƆ�ųf����ؓ��S�D�	s�j�,\Ļ'H��~�����r���j�\�s���x�V��
�c���b8���Z��Q��_ͧ��5����H��ԁ���\U�N;iN>·�F#�TǙO��X�+Έ�����¥#�U�ȗ��KM�=LҠs�Z��x�J������f��@���jt�F(��Ђ�V�4�nI�Z��U�9�GU������3Pi��zf�̠�U��M�Iz�ʪ6J���-|�클���QwG׹�a��V5"�_\���Sݨ���bqmf)�6�`Ԇ�X�0o��״����u� �8�.Z��5��V�M� �jX|}-�荎qM�vV�n��Rԉ����9�ܧX����,��!����J� 0��� 4*��F �+�<Sb��u��y��vȞ�I����g(a��`P!k�ʮ%G�f�{\��.�<���no�YT���)@�k��}�TɉD��{_3�� !�)ze�\bn5E��X�y=3���e��$���ߡ�e]~�u�����#����Q��4�֮.�Hz�ɚ 7�ހ*��1%M��q�4���BeM:��fZ�K{cF�S9�[N{k��2����C�k$��uZ|�|$�ه��K�O�ѻAX.��>�Og)�\#=����>��}c�p%���^��o'�AA��@l��t������r�w����z �CI���$�k:?ht��M	��G�2u`-W�8Zp������i��d�$��@.�g,�xSC�*\�6��Q�4�p��ٌ3=y��'	��\��I�*����'Η��ʢo#$�}?���HC�[Y��(E��������~�C���ߗ`�g%��Ą0�9f��_���D� Xߓ_f�
�W�Φצ)��%�~� ������Vϋ���6��#]�.ꓒ��LV�EF�C{��$I�K�u��Yr�h����T��]�nv�8Ġ&�2_���8b �������CID��g��H�F�������('+1)�Q��vg�U���jP���P����[��0�����Re��}�ߔX�`1Il@�; g���˖��
p����qxm���$�����jI�o�3�܏����7��}]�/���Y����ا�ظ ����#u�Ŏ�1��SK^�ef��cV��o�9c5ݫq&�+╶i�����q{��,��kz��Yu�G�qD����;��l��I�y�/�ym��	f�Bu=}M9�{�È���,�uSPE��߫��_���
/�03���YM�q�#ъ�R��Q_�f�I*C�ʅ�Ñ�(��M�����7����?ۻ���vG#��y�u5ˀ6y�9;�S�6����j���#K����E ��q��L���:�YZ�j�Cc�xf6s�"������gV�������p���+wrS�a���]\��-���g,�F�&G��l�T2e���&@0��v`@��s~~i��T]�t��A`̃@/��E�)�� �Y��B1�m���}tn��J�x���5�<�j��h�O.��4Lx�FϔU�п�6S��H�9��g^Mf!�t2I�&O�\�̓ٚ�EP�@��n;y����<E��ԣ�tJt����J��h�Ϧz�*��`u��T��]O�����;=�4"��(���9U�$:N-���X	@�K7�ιVe9�����7���Y�n��;M���e����嚞� Μ��z'5�UѺ��=���^��s���!��7��U�/^�7�9;�=������xF���1���Sɑ,��d���YM㬪�i��\?�)�w�y��T�`gx��V����\����d����{I��ػ(��S�N�A�9�1�1��l3�fV�H�g}�.+�u���m�{7��%4.7�5�ƞ�]�/��<A���$@[!����7�jR�s�k8>�I�����N�@O4�������������\�Q��A�?q��V=Y�E�p%Y瘏��:�b�{��GV/ʽ*f�i�K�5��.�򀤵�쁊�נ�	VR�����5C�]N����5�B�2�G}cc���ێ��U�*:{5�Pg� �˯}=����$�>�c�7�kB��n�i������<	(��H�e춗�b��5����&�Ydy����8�~c��_� ��~�W3��p�_�&u��ҶB�G�� ����UYPT���W}CP��r������5Ջ2��Pl��%դL��E�*8����/��j����$f0y�W��� ��Xb�Uy=ڭ0�zeV�FңWI�@�>�A���N�NTGQ�V�~� ��r<�^���bu.�]&��\�F8�r��i�Y��)r��m��B��p퇱
&���*'�s"*[oT$C�.$�1�m~r�.��{+�3�����9����~Y�sܿ|��:�YV�A�}U�̵�E�w��x��M
���豦�ʳH�2�K�A�˩-���z�^}�~�h��D�瘍�

��Z>onU�q�]8�ѝ?(X�U�6��ۑz �0
�����\� ���e�y�܂�ո�*�E	ābbQn��D�����������?��nn�e�(j ynj\�O���X^�j�"0�`8���<�7�7���Y�<->/R΋�>7>2P����t�]��&?�]Y��`,�J�t�V���7���^����7�}I�(�ɏ9�=��8��3���c�jz�^����3�|�L�8�R��U��p�k��r��S�JV<���Qe�x��Q}ZV�.Εd�\��M�X�&^�i�)�r��ǯ�ʹ��l�e��v�<�i���[7�bx5!g5;N�R�s�|��W9�\������<VJg6�έ-Ϧ;+F�D�-����)�
Fe�^̓�x��GJ�w
�5�	�e���?^�|�</���I��e�B�a�d��w�w)v�����-[�i���+��6E=���=1�u�[Tskp�	mT|lMrH��*���}%�9�4�e��d_~�ey~Q�ҵ�WTo(��+�I�W�68��n?����st���=���p��k�����x}�M�HB\����73��޺����}�ّ�Ɲz;��)A9�8�v����v{ovqі���������)�6;�P��'�ɃU3l����I��
X����Z�D��K��PاQ��4j����ρ����Tf7Q/��_��\}N����Ɏ��d�zM�v�������$ԩ��=gZc
�(�3H���j��R��+ORA��� ASB�@�6Q�Ǧ|&�V~���H� g=LRl��H�Ӛ��R���f �Y����NŋA�����a�@cG\���=
 +���$����v��׸-V�dU F_!����R��\�m���8��J��nc�J0�n�4����6I";i��W����[4\����!�хq�E��Ȩr#PSs��&��_T[���8Ԫy�#(�$򘏓�:l%�;b��Ĝ��s�3#�տ�������_'�����`�hf�Rv)/�!��k�j��A|s*#7�lr�>��Y⒲"/JV����^?���󕝕u�A��A�X��$] u3��`�#���=�ĵL�u-[�+���#�U�O�f��x�qCd�� �FL�D�ԓ{�^��+29�73_/�����1�jխlY�Z��{���D�������/_O|8��y����Q���mT�4�N�&G1`N��Y��L�B!5x�������^7�N���)���H�,\�w6��#�E����q�K"��x�55���>��x�D��B�J`���H�������pV�2���?�{��<u��p���g*8���\�^�u�ux�Ç��g�ށ�!�����T�{� |.?�T�O��e�k��lqq?W�K�h����Yq����������v[��	�S����:��,�3}��B(�H��TR�,�L.�q8X�H"*�2H����(IŜ�Mc�^��i뉍�O���Q�����ɍ=��bI΃�	|Ŭ��M4j`�Qʖ��׶C�J�~0����q���'�D8����h�(��)��a!S4*0��p��(�
[o�־P��o%X�P�I*KU�[<��� U�ܑ1���!ʄd����MwQ~�/�R���	 ��&EZ�6V�ղ\���D��588îc��Y]Y�����u%�J���k��cB�a>�Tۯl�"�2G��3o���M��/@��wU�;�R՜樕}�����,:1�Ċ��������4�̓�&M�U����Ы
�/ߏTm��FU�ZW Ȫ�'YQ�i���|�D���x:9r��x��s��B96�؊���U��	U�����E��!q���b:I<�A��~]�Y1�\�Z^���$���V�Gۜ5%�Zsp��gk{�lU���I�Ht�/@��o�Jx@4'NI��J8�c�������i��=������Oc���s�[��5�"qת�{Ī���T��?�����t� D�_�N��8MU&�_C/�����UK�pΙZ�����@ *V#+���c��a[8�<T�C���v�}��C��j�a��)�/���좊e�D7��RV�j���)� �T���m�ʬ�ͼާ���0﹪�6�W�'9(��cd��yo
���wX\v�r��.�4zrP✨�$)�(��(Z��j�ZT�1��&Z�O��&! G"F
���Qb�F�y�q85
��Ǖ$��P��NX��B��#��Mv6)�jҞp��lS��d����E����R���dSl0�n%rš���95FdOE��]ISd�$)Q�c���8B�c�#���� �2ډ.�EA)�ұ��l/��ٷ_���-6�$Z��v+z/7k{~ynW�p�'�
Ed�ˏ�U�!��>+>oC�4��`������cP/Y�N�z_u���jN��c4Y�A6��b�
��NL���)�s\�H =NYq����W�C�f2�� �ǈ�Lyͤ]�V���y2�?��f�����-�@��&Gm�4�_S0Q��*�y��ì�Bx���4	�yuk�	����M�7UZ#??S.z��S�~��0��_E�uB韃ﱎk���r\$������8��q�b�d������pcIߡk���e(��Y�g9R�p���gW��_�7_˯ϟ�`U�$W�y��<<��}���no>QA��]�ɔ����8��9�����̩�g�e����%X��r�&��A&�9Y��Pa���~��8�lG�%�>�:i�ա��/��7��Q��F2$�"�=tN5�k��P%0y?���ʚx$�j/�2P>pߚ���5`r��ZD�Jq���I�x�3I��E��u�p�E)Zb������4��H�p&���v�0���|6�ϖ�[�N#{9���c�q�{PaC5i�o��,�[�	����Jq�͹�=%�cu��c�/<)�aP�ZD��b����*Y�KK���>�0Go���ᐬ6M��j��5�=�2F�����٦$Yg/lu��ߣ7�4ˬF��)"R�rU��b�̕�Y$;�#nxV�3ٜE3^�֝Gג>��|�UU�A��g�'49Җ��?�w�{���H2XTX$�Չ]lZ >���� f\ê�w�I͂7�ȕF�T�MZ^�]4_V�ܚйV�e6��=�#-�#?���`b�i>��^�#		�@���!�f� g�y d67BO��k�8E�չ�G5� ��׮8�u�G��b��}����ʞoK����..6�Eƌ<T�2�3 P�}�3F����?.\S����Z�� g�'����$Z�vv~mW��n�#�� �`�uqA�zU<q�����sR�yShD��s������߅�������=<�1@��#��[�RX���;��hJ�㠹A��0�b�x���H�~vh����H��I�BC�o<"�j��$	���}��F�dOn���O�j�v�M�_�^>��Dple�ެ;/���='�ö{��b.�t��?q���Y0$lGN.��b�@͚3�`O�b���  ���t'��Ddn�ʡ'# 2�w�=ˢ�b�A=���{e�U��.ضs�_��`�@�z{��?��u��k�h��ׯ_3����n>}*k�A�*@%J+M��a�sB?:�Vv�\.^=����R�eeh8��&�.����\�9g�z�����Sh�g��T D���b�f,�}�����k��|m_�~n_|��dN(D�j���u��M���Nvy,�&,X[I���FO�_׊Z?�O�mra�#�| ���|� W�l,�K4Z0\�(�p��z��r�[�G1Ɖ;B�vOT�}�=C����89� m�SEI��^�����G�ۚA-b�������ʒ����β'�����<' )�T���k�d�ƞ�v��$�qU� NJ'~�j$�����Y�0?��ad'�V����.�r��ɼR�0��qQud�+�k�ٴIyP�~�v�W��9W�(���B�#ΰR3\F�:{�c%��p��eS|�����x_6�H����m��dh��IV�"��4Zm�g�X�,��0�3��o8�xO�P��"���\��z�0�`�����J���*n�E_LM�j�>�H�@��(%&b`i-�����o�=�r'��D`�rn�]��X�^�� ��aY���2"p� �j;�S�D,̘5��$%�y�Ì$�%�f��\���Z�wTŒ�Y�R� '�a1��wP�9�=%�>�>E<(<.�01HeCI[�J5�N�6��4�{�TS=��>ֵ*Z�f��I�h�,����U1�gdO�ɒ�G�^��J��Xe5�Oh�f0��8�6B���T�]I��t�
�Aa�'*~2'��>3���/3�����r?�)H��%�������0 .�ڄ��^�1#^���`�l�b '��)��]��#�����/_���qss� �i�fkȳ�P�cN%���	�U�#�r�|\�\��c�J:ڷ�F�U+s��𻹣��|(����-�y�W+rjF��^�UH�k��= ���DU�Z�G3)XĠӾ��P^5§}O���m����.���o����_7tJ9��@�D�o���%M�ЪJ�=�ў��n���we_*�.kZ�`VI�
Rc�y=]�3���{�z�+V3<�,R���pQ#g%��ߐ�~�C�9P]t�>�^�I�
�XׇQ#VCId'��z8�b��d�T�b��je�`�R5.X���|��4y?OC���X��lʑ`LޏmNǔ�nZ�SJz �����Z�X ���`�X7��ͼ����[�6��p�������5�h+��6�� 襜|<A�-��K'k��� qs����DY;ǸC	b�����DŅ�#�ׯ�p�g%�����C�w~���ەD�ű=��J�~ſ���o�֌��wmC?_�HM���9��Q	��)/�V~��B�>���x��&�+��*hF�s^��\��&��^D�0|,���V�'���6)*P�$�NX�H&�2�ZM^U���Ǖ�0���08��ᩭJ�tq~nis���-�K��X��r��:S��Ĥ��Zڳg�낂*�����޻��%��gc=&��ɖ)�N�Fk�(O��z��ั� �ñ��[T��;V��)��Ii^���T�]��_�� �5��i��ϔ�$�)3����6��IeExm��-����1-�\�d����=�by���Ώ%�L�R����=�(�.S�^Ʌ�w��jP@D<=�T�"U��{��^�;���ٯ7k��I���90�CI�,�/^�D�����(��-�^�u�­$��I֜c�x�$�=�j'�ƞ��D�?����H�����5�E-�jP�b���.�����z')�%
���[�L%G�`b~�f8�4��򩫵1Cv:*���0e�5~�#�z>*u��%0 1�(7�U�J�QR�=�4�}G�İk}�US7�d�s�R��Z�`�ltJQ���>�[� ���i� ���TP'sP؋u����ÖO�ZXu������4��
i$�Z/��]^��w	A�I=x)�G�N���Vy�5���8H��l^�z3xb���0��fL
$(���F��ע�֠9#����F�z�$p�II���QmJ�U�f}Q��ܶ�j8n4)�ӭaj\�s꥽U� ����Z"Jh����a�N�r`�Z�a�񡁈�j�����H��:q���PSc��8u\��7���ݽ=�=� ��=<>J��P^Z�َ�"M�Z1�L�"�X˲J/�1��6UR��Q��k��<-Z�dW�gZ� C�����+)9ܬ�?hr��U��ع���V�X��t�ChAU�-�÷S	n ��K�����3���$\g.�O�A<2��e�}�.A�㑕��d��f����Y�~�F{-h��p�p�sR�zs��+����=2����P����c����>я�*���V�F�%
!!�X�Q��SI���z�K�z�-�U5�*>v;��82�H�`��}0���qD�i�l�U���ڪ� J�Ԁ�K��㘃�	�|&H�tqNe�W�\V<�T���`��Q҆j�<9ť웥�h��G�^9�8y�[&j�VV��U� ��#��G� �
���}�v0�+6B�]����L�`�Q}&�A��>A�Ǿ��+�?�_���t��$Z�%Y~�Y >G�Da]����� ��f���{�����f^0�j�-��9�k�+{��`��O�So�*%����X6Vt����
�s�(T����k�=�!�CJ���bD�H��t ��{u�̙RP|���&zꑜ@��������1�j�.	����d�8ʄi�2��o$@����fNp��M�w=����!�S���?�Q$Y٫���O`�뗂}`5<��h����x�o���^2�q�$�r�t��'��Sw���ż�F�}�a�RX����XmJ��
����ǮLG�K6Y$e����:�����y0�� �-A���C���L����.h�i��#�� � �  &���Gu�p0��Hk���^ӢY��H��\����Q�͛y�ɫ���@��ig��ű^ISޒ7���7o��o~Q���>~x�_qSY�j�ioqSue�dM�|��!�
��~~g���<��<��On�E�5��g��[�H���)��T�E�M�!Z1�K!q<R��&Y}���64Tt
k��j04.0���u�3jٔٴ>�Q(�ʛ3p6�s�JcG:/�G�dX�䰋~�󔇹"�iD%G�}.�7���>�&���+�����	�'���i��ZP�|z�q���3�z:��j"u��B �D�ZZ�e�U��D�>s�#�<�+���d�+;�f��D�T1ȳ�Umm.%����lg��{Q�����=����/�'�����������%�ыE1S�H"]Z�u��_��c�����Ϙ'�� d�ׇA���wt�^C<&�{
�"��9���uF�b��m N>ӣ�'��/^<'2;�u
)`������a�����?��r��*��'�.�o;ՙ!'�~M]+���8`�+�Ӹ�k�(!�	��O���s��O^o� ���I��[�|}�ad@0Vw7Zh���Dj�S�:^$c4x�P�z��,A��$V�k���(�`�$��+ϕ�c���RO>�6TӴ�$ơ�Nܗw��R�=���K�F�Q��E�埜�	9��߿�'��c�������6��ugw�����c	�o	*^���s�ZB �j�P���X��0��r�%ɺߖD�f�$ι:�!-\�Ŕ�LJ�8%5�x+pcP؎5Y�~�R�"O�<�]�+�L9��z@0H��;%�JrZ���|60������1E޹5��t�BO[
���脃7ֈ����4��/M�#]�R3�6�:��%_��X ��,c��j~�C|� ��+JV��U���gʈ8�1,�!�g��:��bC����=�$����/~���{�$�NM�H`�?f_�D����ߓ�dV�2��s�^3V�ث��i��z�Ђr	{��H�ZV����F�,~�Z����-Js��UK��v�������U���mQ�w�b!x�6!3�[��յ�_]��⌉�6�oT��2�m%��fQ19�3K�O&����+�H���p�5s�Ig X��S��y�u��cG��q�C[aō�z!�l�a��K>h�M����񡽓'BK���D?R$�ɓfO�L �*��\���N$�6,ՅUA�f�[1�0
!K
Გg�H��I�ϊ�u�"�����?����at��<�)����K1d�9���l���n���v1��%J\Njh�f� xѫWF��y�����0��?S�@�k ��<2x$YOO[���#s_i������s6����PB~�;��2y�zX��[^�zS�0�SM�8�gƶ�9���$F�O���|�hE��Y�LDR������J3M|.�v�|<5k�)� ��j�Y5ҨfJ�"��w��40�k�x�B�f�����6�������W4�md���h�g���;5�s'�+����������pF�g�{�~�{]OG�Щ�JΛ��:�t�'ݳ������s�U�aƇ��?>B�y��|��B%��@���R3쇱�(i'*��5s�t�M�H�["B����W�T��V"|���$NH���+6�#Q>(��+���8�}H���������_�ʿ�p��/��\<�%�i�S�H��C -qbQ�["]��kp�اJ�t_�4{֌�y�	�-&�M����%�����e��K	W���b�Pɺ��"==XgǕ�6��P!E�*�{`�y˦�-FuZ+K����N���b5Q�N
��	<�WX�������K ���6�he����O�Tuo�� d��V�$Փ+qŐo�@�'�g�I,��!tP�[J�c�ñ$Y ��2{�B�+�/6vu��ͪe@�YOL�6k�33ӈ� {�u��m	N.J�|�ެ�ؚ�k �S����\*<����b2��?}��Y+���u�/�mҧ���GQyx�>��hk/E� f��<m�����0��ӓ(�H��5�CȂb%�;���>d�/㬩,�E�3�}���[�mM�D7���OE�@��G���U�U&m�՚������ ���T�Hh��=�6�Ώk����4���*q�N�k;W'"���S9�����z���J�B��b��x�����k��_'9��i�Z�=���#�m�;诺,�@�ׯ^��7/9������[�{��{���<$e�Ϯ��>��*���g�G��'��u�G��<�*��i�H�d���k|���������y�Ǆ��sP� �%���I�Jk��!EbtMWT���y}��)]�D�x? ���v�$� %�42.T��h�R�l� 	@bV#m�94�`it��뼔�_��bdm�IM��|�&9=ܯ=(�c ������^�
*-/�0��T�0�]U[�GG�� �����yq�hR�5'2�)����~?*��'|M}������r���|����R\��,c����f�=�gv9��xm�Y��~��xa�W��2��:!��愋��n��2�'tlz�����D:��-	e���iVFme�f���L� o:l�79��	%y��<�=�?���u��H�n������P"���_}Y��%(���h�/J�]+��L�yI,n��Y<nd���$�)�}U�uocK�-�*��]�`�T+l��*߸G��wj�G5Ys���_��L��~��0Q������+?[��ʣ:{�z���tnIX2�T� !�$�{;�>��⴯��F���I�B3�4���ڣ�SSw%E�V�=H�`����c��5���A���#m=;B}�|��n(��\��U���n  ���RL3j���yk EzO�$k4��Ve��lU�u���Zh*�Ȇ}9�����������]�u�T����{�/����>|z��{��/I�.�����2H�u��Qť�P`p�A{ b�l�ΦA�m��/�*��<6h��l��}�|P��)~		��� �6�q��j�K��N���GS�d$�=e��N��]qR�Pa�a���J�s� =U�t�ܡ*d5������=��L�>�=$vs`#�C�����)�ή����ި�zp*K�y(oƵU����%A�Hz@��L��ޥ�M{S��eYG�fA�Zs0P}���7vw��|>(�O.�5�Ep�'4�8��cr�G��
*�;DgR�'JT��M�f!zC��U�R :����$��k *p�h�B��2��I����
��� �^k*Z�wDy
�gJ�RPSE�Dg�JV���J��XN�6y_M%�� MلwiO��leW�%h�:#]Փ�s���DU������.Re��d���ʱ�-ǵ������^�Y�ť*��Z��$0άJ��WPp�V%�$�k�3bI�~�MO�^d�8�h��g�~o7�����޾�D�����Æs�XQ/��aa���Th����Y�x����b��g��}߸z�D+h�a�(��yЊ��!�y�(b㪦J��c�k��.����QxdI �Vt�>��Q�IT9R���1B��yyi���oʞ�\/��!%�E@�+�LtQ$/��T �6�����uyn4��Q�$���M����l7�ʞd\�F��\g�����{�D���GrUޫk�! ��\��Ij_��H�������P�g��%�(�7%�zc�^~�$�u��Q�J���?�ճL̞�|�jaG��g�+,P�&N#R���Ŷ\O�Wi�Ť�0b��{��f}F�%.hx]I��.�Hy����%�: z�Ʋ�'X(�A׀��1���¹P��Wn�-�;&A�S��ց5l%b�Q�-A�Q[t��'� �)�dmg��U����?DÎ���w�{�o����R�XC���d��a���_h���b9&�[�$G�fb$J��,�ţػ� �I�X-=�F h�����\��F�UYˈ���ѫ;S��~��K�S��`[b��r^O��@5lOM�5Ɋ���D<bf{H]X�Ka��d�nF	��b�����)�:X?�M��QY��9�#k�=�(UH?o�UU��l�6WJ}���� �׶�EB?�����T��9�\�/1uog`�$�NW�-k�&��C� 	2Ÿ�Һ�;�%D�y�ՓY���0�x0e�Hİ0a (���%��HА�V�hdY�4�oQ
|����=E9x	3��٬��� �WP "K|1~m��6�Ϳճ�Z��?_�gv�@R��� �XX��/�Q+�F3�`b(���pP9���Po�����2��1�����}	�MF9���F�7-Мg��y�J��	�d��Xц��O�_�s�Ƥ)�\@�v%}�h��D�H�d�g6dU����M�ڸ�QTW����R�,^�)�|(��	־%���l|���;��-[W��h]��d��]1p�G�tw����=n�0~���7B��Q��qt^詚i׼gc�m,�Z!�5���90\�,*9Ut2g:�p���<g@b%�Nmq���.-�Kb�8��Ԩ*��I��Ps��c{Nj��{@]��%_�Ag��Q	Z�HK[qb��'%���j�@��G6��q�Z���d�}��@����=x��v:�	L+;����*-
��v��|6�1;(1� �/����^�ib.�	IľB�9�\�S�UF�OQEa�Ͽ16�.���wamb��_.<�j��i6W����S0y��q,�ۂ�(=��"WU��p���:j>3����HO��;��9f�K�_�� ��Lj/*7 �`[.1�ƕ�Pт:>��$�!,C�S���9&��]�΄�Nޙ����M̫�9�ꂑ����_,���b;�P٨�j�05?�;��z��G����Ƿ���7�=f�(=��ơru�c%��đ?����ڠz��#�$�:ۊ�!k�U�ݑ�<ߋ��k���t�Fw�k�L���䪧Gk��R���cXQèҞԟѱ�j�cP0����9����{�ȑdI�@
jVuW�u��}{���̾�3ӣZw)�$3��03� ��gϲ'�,2�����\�/�����&
:�8�N�G�S�^�}�g���'��G��*�-R[��CN�|��}?NE���#�h�f����y��c��z`�v�G���y�g/���?��/_�/$�>��y��k��@�w��A�7�|C��ӯ��Q��e����q[�C��(.�0gc����@��MQG�s�[);e �N?T'��1G��������	x�N�V���y��Ǖg�&�����;�2#�-K�+���jթ�[��
�)Qe�6a-PH�@��k `��r����5���u 2�
� .�S����'ZaJR�,G��ǣ�y9�E 	{��,z�"� ��,��I�1��,p��������A���/�~�wp��^4N҆9yYB$1�n���y�I�R�6i� �{���!o�%�	�s��E?Jl��Is��H�aN�c��糤m���}j{q>S#8:�,ξd��ZO��0����z�� ��Dj�| C����P"���S�PӾ��{D��q�EmN��O�תY�������u�:Q(v=?[���9#���w&��Ņ�%�n���?*�F/(	��Z#�80�˱ZS�J~�O_Q�Ҍ�����Wѻ�$]�,eJ���x��Mtx٣g���hM��<9<�RNU!1%v�B��6w����vy��=���)��m�>�?��`� %XP�����:�A��� ��!�k�*��������|�)�ytІ�mra���^�*�i�H��z�t�Ǻ>�v\������_����~����� d�m[�_��t^�b���hwh}x<�g��#�?��t�k����?���iN�@d�_>����ش���V&ֱˡR�.�#�ЗQQN���]Q�2X�3��}	9W�Fk�&�e�=�z���A-]�	��ER���!/���� �ж����X�t\�T�,P����f08�8�g��x��������.�a�\O����,�q�&"{-dzdM�=�̗����mH;Yy7�hr��P]`���b���>u�c�~싒b�����th�P��k������pN)��@�J��џ�M])���d
�P8�_��/;� �5�+�`�b'�a�8� @�bZ���9 ���-��������E��G���,�,`p��;b�vl�G��><��&���n_�:m|�-m�7/��vPf" ���:�$���`[�`��X���9�:��u��(X���az"����������|k�}�����-)�����#��L$�$̪�V��E!�x�q0"��y�u5����u����</��N��+g5�-F�,���JC6X=�|8Z�R��<{����91+r�XȞe�jSZ\6p���Qm?ʬ���ܹ�7�>�BQ��>R���u:K/,��~ó�x���
��N�[԰h+��/g;�}�� ���é�#��DlL_kc0��'�a��V��㏢^_]���� ����o9��;�P���Q�V����6�&����ڻ�'?��FVhH `���h:K�ʔW�������#��H��w)��3�8��^�땉��S�_�L�P��q�l��cO��f-�{��'���pW��Ș-�	������ k�H,H*�y�D�3a-V%��
�p�R��k�UǞX���:R��(�^�gt	0f�=�[���
�JL�8������A`�=2�GMo�-t��N"P�T��-h)��e��{\��X���q�=4v��'"E�n��L��lW0\ȹ�$�)�FР*:#3���X���b :C�����acۮ�]wb���[�'�h|^����::R��59����W��wzm�Je����y��<|E��y�lQ���lnFdy#1x-�q���xD'�D�q�����=�zPCߔ�_ܲX7C�S=Ϊ����߯l[w���_c�\|ضVH��A�3Y�x������D�Nj#�(��L�����l����Jrw�����@	Ϻa+�AǙ�Ӭ�X"0�d��J"sb��E&���:gvu�B�Mu�� g��\Yó:�+/�W�Sdo}f��Ac��<wrpdFԛ��>J�P���Pg�>޿Gu�2s�S8I��P���└�	��;�����{�����z�,����q��H���7�>��\�� ~W((6;HH?��N�< FG�D�p��3��x�. 0֏�)���L���]�>�[I�¢���"N@���~��f��6ƒ�F��#GR�@s7�#`cM���Eq�a��k.1M��'�ſ����x�4���}�nM��k.��Ȥ5 k��z>P[؃��yD�T"��ش
��V۩L���1�Q#S���k��<WQ�j���1e6w0�n%j�r��Ң���.�7�x���ܥ$w�X~[�m=o��Ɂrd�X3�@ک�*e��͑���5��P�����1����-���r�7��M���������#ꅽ�A}����+TQF���:/ê��jW�7���a.!jS��S��
����Ƚ���R�,Tj�B"^U��I��0�3c�c���T}�ǶvA?�z�p��~��;��o�ڷ���:�?ػ�(���,%F8�P�&Iգ��� ��D�!֕��{e�x��� ���5d��z�p[��*W�#�Q ��n�ˣ9�ʔ�^�k��9�J���+:�E5�,gbψp���8�Q�� ��q�@I'�tD�1^� ��A���g]l/*��3�
���F�w��	��#���T���1ꘊox�c���/ڞ�~H��,��(�Y:��"@��/��}���ֿHr����?��*��p�~���.��P��G2Zp����(�]�m?ӎf��R�	��+��N�=�K%b�O�h)<�x����I����w�&��T�Kz���T�<�^*y��E��*�xwg��{[����^�ֵt�����}�g��
F�;{��j�^��A�{t*q��� ��o��ds�>y0��)�U�R�'W9����Y��9�������U�O�s+��m顶:&��Igt��OI�{��w�)۫f�#�:RGf��!�`�00� �#z���8z�z�s-�%J[���k�g/A�����T]P�W��LX~�k���b$'�D�r�d!�`�?9c~�'�/��Kw%�;W�iރ5[�&�
uaZQX#�=�F�b��"�x��>I����4r��:���J��_��tnQ��%��f����|M�sO��K��������u4ޅ2����׆H������͟�k�6��f�"/�b8�X�1������.%��������h��i2�>V��C��	:t�N0��BՇN�܀��}�&�I���	�#��>T���4�u���>֔5]������[$.��ʃs�D������)�4�G���Ϥ����r�1;-D��ȑ�Ʉ�Ի1d�;U�ծ�N�;�B;����ݱ>����T����_ޠ����@���� ����,P�z�H�CJ�0��� j���s�8��P�H���s|���\H��U �o��8�����{Z�A�1�rP�:7l(N��,Ce$�Yi CJ����{�K�0���6�I�`iFJ����]�ߒ6|����� �å�����Q������­`5�m��'�붙��;5��J� ���Q���wT���}�||PB
�9�%v��j�9"�Ǳe�� aNy^^��r��mk����X��ř��Y>rY������7T9��(�Ny�>U
.,�)�I��.f6��T�TDL3�P�S�
�;.ګPf�Q��e���z7�Q����H��bO�l���ڋbw��
�w���d/���n^����K��֐R(U1�����`���KZ>�ؓ�w�Gm������?��?�������_��W��?�I����Q���68�#���d֕A2ֵe���&������{��to�g�B������1����M�M(!6B�CV6�p�NWd�=����I|�՞��Z�!��v���KP�t��Y��Cj~�0K�*��� 0=x���z���l�1�n�޴/̙���ո�䈂��y���m��U��v4���������>@0���j������ATH�����v{s[A����� k_�d���+��^���֞��&kʠS��&��19	-�O+��V�tD f�>�3XC�8�N�R ��L%e�/�g	�p=Իl����Uy��y� R�a|�w ��ٛ���8��{��I)����~��*w�F��*ɤ!�߉%��F[7��KZ����Sv��2g%P�Ne�h@^
}��e?��:�O�^���u����x��H�ĹI&�#�^W�	5��T�s'6�h�AMԃ��*���T�gZ����t�:7uBE4�?���;P~_*|q.�(0���Z���C�Z 8!f'>�ir�����J���3�@#x�3�#�p��Bai,�Pq{��K�N}a� +�(c��h@}E��Q�E��m���max�kv\� ks����~6��ۍݾ@?��`:|�:g*��۟N'�4|��?� @i�����]<��(e	����h���==F��yv�i4d�@pe{���:����C� �Y콼���,OU�r�����#��z['�|�!� ��lʃ��f��M�ұֵF\<��0Nx�h064��A�#@��|MJ�f�8�O�i���08U����Ƅ�y��(��T�V�=U�$Äz���z����'DP��Y�Q)��s��1χ�چ���,Fg�4ydCJ�"�+�R�`��# F�k�e��
���+$ o�e5x֖.C��.wl[P��H���8�a��;�!��^Y��k���8��+���˃�[9/��;'@�������J�ЅhF3�NIi
E��tՌ�!�[��/v�H�>6Q�s�G}��s#�H8�cO��3�w�.����{cMYb�	�E�=-Ԋ�F?�}-a�w��W��(f^\���m8ԋ,��S�u��`>z��q���� �^)'�3��Cę�H��\ҧ0.�Xd�ln�j�6 �~ꮅZ~��:�:��S�&�*��3�ڇ����qy�{[�ŀ�g��V�lw��}x8T�����HN�������\__9u�7'�^��(���#T��(���4<(D=���=���3Z������?�Ο��QⲔ�Ы�����7T�)�B��:��z���υ��}�(��i^r8>!b������E�Ȩ���a���Y�u'Wq��w��g)d(�'sa.lo�}-`2[X�m���t�ȡ�}��s�f����!������E(�_�:����5��x'f���s�$p�PAYߖD2M�V#��Vi��|�T����� @g�Ƴ�
QS�җ��8?g#]8w��`�b��-���Ai�̅R����FA���%�cm�#�Ի�K5X��^����E}ĸ�+O2[�F��Ȗ������M�����88b?M%�sMc]=?�����*�� ����*	RMb�A�]����W�o�Igų�%�Z�<�����KJ�	L�-��4Q�Is��s�T�@�S	t���ߌ����͗��ī&��}@�up���Ț7�o�^��$��`U'���HG68g�܁��� 5�G�u���j�)�t�����(�$���S��&j�f�lGP<����7�7�m�ƒ�m���.X���o���1E����;|�%+�o~{@�~}z�5�]� )P�{��8�k�Ω*�#	���kyt�?}ɡ�%2\���J���o�(N�|������{�{���^�O�խiC�9{X'4
a�&�E�s	z��rBfV�5��y�T�]b+�o��:��/����{�`:1ߦH��p]�i��i�(CV]Uز���p����A]�����Æ*@�gv}���+��H�h1��MF:�N2g-��i��8�2�f`r�!+.��z�'�Z�i,(Z�HdϬ�)�h��C��� y��"�zT(��45FF���uXPמʚ�2O�K> �)��h(�wF�
��8��<��Y���
��
2�*�� �4�~��-��X��h-����,�X%�7a.S�i�1L>o�|�v(d���j_8�y��E�Ii�7�kq ����%���%��/��>)�:=�����Ȅ���X�1R� �d9L}P[8��܍={T9(ˤ-�M�X���ߠ�Urʂ��g�`�*|/^/���͈��<"<�a#��� ���]�����P�|�dы���fl<�:�`����b���@A:��Y���}�	p�`���v��tə���ǯ�ޏR�INH웈�R�i��� ���>��h�];��,�Q*�o�+�z� ho�_^�3�nV���^\]?�����l���Ȱ�J�T?�}� ^�SS?��3����`?����y�`���ZG�GzY:f�rRmU�Y��E0%�Tu�(X�;����
�3�������hw���gm�W<�Bgi�\`�X�3^MŊ�o����#�*�O�&њH���:jf��S�P�4�a��<X����Q��e.VT������?�^���k�����6��"R��g�!�X(B���ym�s�|�䎲7ԆC��ϫ��zV_1����[��vd�����ͭ������wl�Φ�!0q؏���]��T�@����if��8�j��Σ�m:s���e����Z�N��(t�PD4v����QBb����2;��� RGR��AA?�r�({�z{1a���UG�	p
i�U��M���fmW+�������:D���h�Sh`���ʨj�R���ˊ+�!1�I���ͣ�Wֹ�)��ɛ�gǺԀ��I�}*�]˪X)'���EW�lS������X����.|ΤzG�桔 e:dA�
O��R\NC�R��/��c���R�ز���*	E�~��PA�qRfUBk��&��9P�A4����Y�[ ̧�	�e�,N�v��x��5�������1yb�_�|?��_��
�!��R:��tV/Y����  Q;�tz�,����ݶ��r�θ�����I)Q�#=�Y �6-
�A��-WHwN�`��"ʒ�>����)t�T(�tl�
��� D����%
�N��?�}�����%�K�b�G��������� �2$8'<֊����;��G32�N4�T��z���{=0�5�m5�8XQ<�Z-Pd�#Be��̩f�}�oʙ6H�����5���ӻ�U�O�'�qr��=�9�$Ox����F��;�.�KL'���NB�Y튑�z?�{4�0`�(2Y���J��\xx-t�I�.X(�>�ы>"!��A	�_+
�M��ŗ�ظ
dk��螱�	s٫�\X��B
�<nCnB�h�Gsr��X�� ���t�0'����T�Q�+ҶȤ�Pc���R�&}��,��9:�����j��q��h+*��>+1��@�c:�,�c޶���~�u�Ad�d��;���.X�{G]����]^^گ@�Ț�IA����*|��,#k%��4�L�8ˑJ�׋J(y���`^G�}%�5��g"��yM����2���� X����ܤ񶔼֨x�I�&�����Ί�8�6.�:��N�L�Ank�����{��#�gu�tf�9����5�h�ժ��K��5/wtnQ{��v��V��2��A���|A�@�B�.�?|����~� ʁ��s��y���أ�q;YJ�O�F�WD�J�zY���,m[�"�e^��A	�����<߹�`�@G	Я�cJԜv�����ŉ�_�<l�W%+�!���_C��rP�M*dw�u�ʹ�(pތ�����f�{d,�|t�zխ�%��% ����=�h��2:��k�����5,�渻�1�t ��I���@RV|�5"ť��&�hɢ^.�P�һ�� !�/����@�ݽ'�z���%2XW`������?XB�u�P�.����9����?�����S�b�M�z@qے>��+�4M�I�4�+P������cggkR	�H��lv�5�1�70f��(:T8�S֎{;�G���`l/��V�������Y�mn��������Ϭ۬��s@�ݣ�:�N����
��a;�sL�	5I��s���8zVG=���	:�6���h�.��٩5��z�~���~�J;�l�+�[�9�~\�g����OV�r�:6+��0o�1_��m _��z��
�����;,��˯T��c`H��w���{?��Gj�u�\?�a��_�s ��i�xU�۷H_vA?+�� �R�����kɸ[�&�Y���g?���~��ꘃ��V�f�8l������~ �����2�V��qO�3�:�:D/QgD��N4]�<Ç�Y"�9��Hc�p��?�Hm`����(Y�V�q�������Z�w��a�T�ܠ�P�Y�by$�/��M�q%�U�r�X���D��>��I>q �	�.
�+kv=����y�hEg>{�$�kv/�����l��~�g��*z�C)�8����)�߉s	S4߽���c{a�ދũ�A)է�F�x�����y�{��&��au�LC5��
��#ڋ��$J���5.ku�_)s@�����C� .Lj��jH�H]�k�y�c"�F�V�4��/�I�ʞ�g�T��#�D1��ܘQ�=h< Up���%���<��A-Z��!;}�h�h� ���z��"5��\uA�?����t?��3�S�JM��m1���+�]O��Զ�ɺ�4�5|�?|ۅ5Cѯe�h�)��
�r���z4F�&E���Zfp�����#����=�h-�^?�!h;�͚�6y�D�_�|a/n_��	�e�Zu.�zbb��CJ��j�N���k��ʝG3U��=��ن%Zp���������H�k4~`j��6��s̳Ys�)���UHW�p���ǁ�5*�}�=�Ӝ{����]�3Ǐl1)�����NL6���Yzd��(z%������Ov��"'��vκ����Xo����=�W�N�8���Ǉ�����W{��]�����_�㍽}sG@7"S����{m$kC�2�4�.5�m���`��4���i��h��9+[�Ϩ��7E?��*|e�0O��e�ݮX���{�̩X�u79�����z�ǵjv�@ո���A{�Ƥ��!�qžc��{��q���n�Yt8�k̏��P<�:���u��c�6
5�nl$���%T
9�^�I�Y�t�����:@&����^��54��b�X���i�w>�Cؕ�������?p�!����:-����8�=�_}i�_�F���`�ԍb~_V�t[���Mu �q�Zd��$�|8�t�<��iGS�ef�4�o�(*&�zgda7�#k�>?=��K�q -XG[�_��y"�:	��SU�<�Z}ꢺ�n�ɥO .��;y������}VA'������/h�T찬�Ӱ��H,����T�:\Q�y*�uՀ UX9�B������!ұ���`�����E�o')BX?�5E��������.L4�&�x��+�䄢v��lm09�6�%K��d�1��hA���kA_> \P���.��/(�����Z&�7�	[��|Wk���3�k���I!���dL6�j�TFo�������Z�1��{
�I�+ڑ�
�X;��܅Gg&���`��S;_sk�lb��s�>����~� �x=Ԉ��S�>(���N��@�*�����f���Zr˞U�OR������i�
��0�!����l����m}�ȚgU:W�46yJ2��+���E�/�OG�xl��ӯ��¿����3��0��o�L-"H�s"jPz:�}��	N�(�<�TQL]�� ����9x�B�c���������{:�ח��t!�����F^i�˦"��ă��|rzD���/@X)�٢����N�ODw,r���YEA�86��&f6ʤ�P�
�\d��)g�o���w�[ׁN��ƕ�Z��|�؎��{dL��Ŧ?<�#\�='�X'�vf�<S�莝PO�N��;wz����%��G���X3ɍ�P�ͳpY.�Pr�v-eϰ5�x(I��&wV=�Q��={=�Z��\�����.�wCۇ~�i�i�|}*PP�dWZ�x��~;�nM�hs<�}�����i�����y�0�����@��Qd�u``����}��� ]
�z�L�����Fd��O�p���p�EcݯV�Դ�/�c��X~��v�Ĳ�!�Y��'H�x����@WPʲI2u��Zn�6����?�Q��h s0�0�ޘl�񙋚.F�Sq1�� ՘�����>���V���������%��6*ۏژ�]W���� ����I�~`��gڐǇG{��d�˯�ڛ���ݣ�ywo��=�ã�AR�2PA�� ��2�����,kNYL˓8�z����9�_�� Y�I! ���Ͳ<�L���t���=���Z� �B��P4S�9���c��lp?�6��O\GV��`ˬ6�[�/���06�!�4+��ﴧ��}�m�K� JG����3z>	4��l��Ǭ\G��a8#�<Q�a�}��L�ڒ��A�أ�y)Q�d!�$a�9���N(�#��Z�h(~��״+�������ի���_��_0z����ۿQE>��� `�Pl���'����M)�̞�>�����3o�^{2KU�:�Ϋ��۳sC�ʚ�Y{PI����p?#AȞr��z�U�̌g��?��m]�k���05UY��U݋��v]��z'>�*�ҙ�����cT`��J�-�uoCS���T�E5������k�����}���>���{W�B��(e�� ?F���l7{�&֕!��N�ulW�K�� ���2)�e?$yAJ\�9j����p�k��'�����{�����?���~���qow�~��ZFm}<���2q�ꁃJ�2D�-$����D��H(�#C��-�P�,ԜI6����}]d�yR��<������Zz�~�H�W�+��؟��g�TX ��@f�-��Q�$SȲ;�c�	N�D�5o��dſ�E3]8�}N����"b��vVZ&����^��p�qPm*z><�z�����?���������^��NJ���fW7�H?'�teW��^�Jy8�:��m2��t�gD���|T��qÍ��;�ӿ��F��_����N��<�g*���
*������f?4�"�֪<�3��]��a3#=]�gx�/b���h�%��^�18O�$Y��]E��������1��1�{,��~�Nēm���`�{t]D��z#rv��Ԝ0F}�b�d��5V��L�5����~��x.���'fWێ�y>����+{uemN�n
��Cp���[oJ]7���Xg(/A�w����� ��5Z�f�}v(�f?�����W��bww�U�rT�zi��Pb���ƿ>�Q�d]Ry�S��}�cvG�Qw�h��cƚ1Q�"�g	w�F�ճ���8F�Tɹ��F��,>:�	��jW�Htc�Qs������`���G�9������乹���>ze�y*H5f�	�s�FG���k���tCp��s%M^�B������or��S�����} �L�mD��u/����'i>�<���7Q6� ��yn���!�P���!����G*p�Qkx�&�`8�`
9�]�?s���<�th�-� ub(�9u%���s;{w��_�g�~-HM�AJ}w��j���P��V����p���$\��(I�:ⅉ6�s��ɋ��{��9�Z���t8��w������8ںC#�l����Ѡ���WЅ�x�������ir}�h�������rя�~�d� t�#{��龋2>U[Bm��^��6{4�+^�"#yA�r�V�[F���1���5�D�pda;�bD��=��
��*��o/� l�� Jm�\Qo���B��/�'
I�rI-B�̋joǃ��s�
��.��d�l�)���~��+�=��T&eE���NR��yo�V�� ��g �R�u�/W�v}��9����M\�Ϙ���L�2��M�� H=ltvj�Si<�ieI��|�=f�ʥ�E؛�b��*\�5�����^�������믿��*�ze�W�T����/����O?�_~I`�����Agn�L|�~�A�ы�H�ݛ�L���^�Ȝx�z��n�  3��4s5W����۫[����m�kvX;��]�k���>�pF)0Q\d4�=m~N�빑 �P����R{�>�3i�G־U���go���xl]��ǹ�5mn�g���8Q`����vOϤ�n�S��^�����&OG���N�GCo5�Q�=�j�y]����%�8?�+�H�1��뭮ɱ������� s+��́�ȴ����_d޶���+=%�0��v��ڢ:�%�4{����H?R�R�L��#������cpQ�����gվ��<W����K{y������uvk��{������ݽ��8@,�����i�
�Nt�Z&��8����H�1'�Ua����w�1�{��hMD)5ԟ�t��P#���j��̼X���5��XEy����D�T2�&_���Q��@/������Ͼ��/?���6W�x����#�f����[�ҙ:>ն%�.~`LοV=Hߎ�8��"b�NDA��J-(�E�=���&�w�@z��8�~������������ڼ���"����<�a�1��$�ы9�p�Nn������l�,K�g&7���ema�9j>o	�3�;�7ώ�Ö��i�֧TC���r'����#(Y�R����=��j lA�M|!O}~���m��C���=W��8�!��ʧjh.e~Fu*���3���N�[Og��b�s��A��Δ��:��j@�Q4xuyE^5c�Y��F4&�?$�	��e�A��0y:.:&���;�V�5���z$GO�5*ʊ߳k@z|�Co�ڪ�,�LJ
�4�[�>N�0]P�N�ƈ�D̼���'��ia�;�B
�(�۲��#���OWvjo�+��bs|���G?���b�&Ч���?yA��D�`M	p8��ָ�Q�?.�\��sԂ���SZ^Q���]l�:�ie��em4������0�?��!}Ǧݼ�zȦ1lC���t��@�{��������9��Nt��F��,���
o��d�<�����:�͖��t��)%��s9�̓��9��A�g_N>���X��;�o���+H������9�S��t����xØyeH�:Y��Gl���s���w "���:) Z���I����=*��xdO�jk��6��aD�3W̨O̬�2g�b/�q�47S�řs1d�`9���;��f;Ìt��ɦ��˹�(x.8d;GQ��ښ�m�$%:W<#p'�]M�Ao�M\;
x��]���W�P���iGq+\ "�S�6	�S�U�B��,eyB��׌Z��.{��ގNw�5��65��9x;�����-ȳX]�K����� Y�-5�țϕ�u�CI�F(���=�\T���?���Ud�^��_�b@��￷���o������ݿ(�0��77/(UԜ�\�2:c㚂T���T�|�uq��M��ո�J6��tLC��#h�(M�&��/˱���{S�p��9�9e�,��l*,�D���A��9����ωV	�G(�>���@�t����9�B�Mc����G
@���g��Y&��!F�"�#O�27@E��d$�!~�����1�`N��A�.t�
�=6=���:�w�����p�+(U\g���g��z����_�����a������Q~v�fF,j��6;�\�[�W�O2U�V�zT2���4�'�0s�2q��}��ȞΆ�����`��-�-.��>N�k7j��PV*�
��D����ƩI�îPճ����zm�|�MR�d�<=Nd+�������c�#�#�A絆f(���' t���"��+	�%ݤ��Ο�x���j,znD��B�)c,���}�R�_UC�N��o7R�d��>$�o����� W.J��N��󍿰+�G-h@'����K��������b3}В(�+�_`#��|��FqT���y��*���6?���Z-f"�#��n��K(�I��"��ڃ���P�S~�NDVE�����#
��F��g����7k��U�a=|]PE醑D,bn����ée�SE����qx"��Z<�u��˳3x���#3�N�Z)ӎe�� �H�_d(�����? ����{O������3�KS[�vpY̧�ԪXf'ˁ�VWyY�P�Ru��vf�HE�[0���ЍT�%��������7_����(�ĸ��YjN9�ָ�F$te�ۇ����pX!�0���u�GNN���l,3[�c�'��^�.����s���ͮ��޽{�h�n�Uat-,f8`�ԅ����D/�I�+�ܱv獁�>�r�;Ϫ�R;?�������k�,i�!�߆~pz��-'���o`�?��P�>��M�uY�ȞX[�Qo5o�dK���7Dy���Ś���� M��m���1��?�����T�P�P�'�X��l�'����L�=�&���L}�`%G��1�O\�-�
����/� l����ӑ�1n#�������p���i���+Q;k��f���Tg�v�Vj +��jñ˝@h|�r���|8��5A����ݪ�\��'��GGϲH�P`.��}�F_3�ƥ�y�u���튎P߯:��#�Pa�rS����Ҝ-�D.*Η��[�Śk��>��J6�ZmZ	 �����曯x���@���~��~��'���o���{�M�^��z����L񀀋����:	6�e�H� 2���M��N3(ի�5x�=��Ǆ5�ZEM����L��1��D���m���q���N�f9 j�x�GƵ����^�>������숆�R���^��ܫ���u�+׼�
k����8�Aჰ��S���;�&=���H��@�JTY��Y�g+{��TU��������=�ƴ3� g+���\_��� v��+H�c�Y�gAV�s���A�+���	�'6����(1�X���A{{��W�;c@�����wo߰�6��k�b�L��T��tOe��lmQ L�ț/�=�J��@�|He�p���u�(��C�w��y��sۛ,�=�7:T��K~�*eR_�`.3��w�qײ���_BX������/�S@������2� ������jI��J~��j��&x�f'QX�v~�@�n>�/2�˯�쩿�p����Щe� s �q|�Ru�� Y�n��1Q�eI�)Ü���Sy6 yV���Ym�h;��4e�df�������E� Vs���Z\AʿX�T�ꬂ������t6n[�f��Q�%4<�b��F�F�u#���T?q@�z��S�=�����:kP@�DT�~�:��<��t,n�L��c�cOu�K�TC�J \3�B�o���7��}M�V��A���2��A�2���y;ؚ�N@��(5ؔ�3�i�v z��㨂��(e���=�8�e�I\�"��e4�fܣ���Ve���=� �Wsd*r��KFj^�3���\����@k�s�
<�|�~h>��＾c}�9����[�Bc�v��y�<v���;���}�_3�*-�a�p
T�P-�?�S�)p®;�W���OZT}�M5��lzڟ��#�_�����Iʆ�i,1��ciҶ=#�S.'7�b���)m �e�SjM��B��	�DDpP0Gm�%�k��Sv�S �.������Z2/�$��(��Pe0r_��XiT���u��n~���dKP�7��sv�K`���M:��ɦ�)f���`2��)����z�v���"@?N�IO.^��+���M���j�)���Z��$����nw���Cۘ�?��64=�{ `�|�3�0��l�z��MjlYN/�O�� ��R#�	m.D�F�N}���
d�&	m�F�K �PG5����3ۼY8��U��p{�s������B�,�\���jR�_��(�#j��&�4� a�U�m�*(�����tLN�E�.����L��΃�8������H����嗯�swU��
V=>�l��H �����~��5Y�o�����s޽{'I����I�!-�pZ\�"��~o��<�ػq��Mr���l4�!�j�6�͊�� s��q��e� 3�����?0C�׭L4g��<��}w�hv-q	x�8�7�D|vkW7�Y��������m{�Q?����/��9k�}�{�==�F�h�R�u��k[_��_���g��!{�I��puy�u��=�!��w�G�٦��Uw��5�g��:����`Ί=Mq�@�uy����E@��i� APjWk��Ӹ�:�k�n^���-�
�λ�m��6�`�[�hb}}}cW�q}��n�%�J�~v����K.*D������֐��P��3��C2V
���<��@vD3ݫ�uFYR�Ȃ8����j�ԟt5�2��=f^������W	�����1܋N�\���J٨���sy�⥽�:����Y� ����h��J!��s���d� e%>4��9p
�D�0
-���Ha��a:o�	dš�4��\pH��Q���_R�TE�ձ�wj���j�V�Cu�w�>ѱY�
9����S�yz� �v��/��ً�I�����Yi -�~z���'�*����s����-W0ֱN��>Fә���A�Z7sO� (JA������t@D�]s<EZ!m�2��@TA�XTs�O�I(f�u�t��jK���&q�	��5��{�����
��]G�)*��3�.�ݵݜ3* c p���\�d��Y�J'�/]yZQ-0E8T�:���+������A��X�w�?d�ң�Zx�fD�\�GȫQ  ��IDAT�U�m����)*
fm��
��x���qm��Ώ��Ӻ [8�s�>b�/?�by.|��*x-EPJ��627m���K|���>�~݁�>r8�#����N��S!����Ji5e�wP����\��D��ųw�I�M�ԝg�s��T\%�k��0��Cj�y�f�g�G �X��H�L<�WM��J.���#�U,5
�.h�$���[)��t>
�jr�̞Y|`���WV8��?S��R�iw�'}Ʊ;�~k%��&�6<\<s>�'�|�>րI[;� @�F&	�Do^0����	�R�/f����=�����ɰp��W�����"����d�W~�p��K{CkQ���uJ�A +��#}��N�+��i���:_�sd��:@���QP�*�B�/<�.�Q��ʅ�k�����+TE�4:�?z�B5OF�?�/�P��	���i��+zܡA1��М.���W�Uv�[1���;(������J �b֬c�E�;��K��Cf*� ���� a3v����Pw�3c�|��0�ב����E�A���I�鷞��|�ff��9�� +����f��������D\]_�zAgx�'�z��W�\�+$�1�o޾��?�GB�,8�:#��@�%�s��a��Ѭ:��(�a�ȄPDv+�G��B$ �R�4J��Ÿ��N.T�Ybֽ����`����3s�l�1X����;�>�T����~m�3PMuF�7�� _۫/^�׿{M���B6��GR	?���]_\������>P5���T�ַ Eg���W�! ���i��Y�Sÿ����=�0 J�[����֘��4�?y�������=���T}�g�(�|���k T#Yqssc7/lU�����3{��������7��o~��
.!�t^�����_����g����r7��ͯ�5��?�k�ɷ,�����
ؾ>H�sQ�hV��Br�ɳɫ��qT�/6G#c̒��k�db(�.VS�����\{5���g�]
�N.*��P`���X#��y��czu{�q�\��\=�[&d��2��^���g�]���G�,���o��2G����90�^}t7��L[D'=����}E㫺�_�^1��:�X�0,�rvF�9S�����.�g*μx������XZ.�@���ZK}��'Οi�;ev����I~h���%m�a�-��>|y'K+̫���K}���b~8Xݠ�]	��?_�oο5)<ɰ:��N&�rR���%�l�T��g��="wu�7��}���Ohe;RcDI�
d���1K9��>� �Ų���,]J�R���ep�|�mJr���U�*�f�Y�E�Rۓ������|) 623�=
�	�(�	��K�N��:]�(�()�!��W=r����oK�ْ� �������I��E��X�]�Axע�Y��x�`8��|��I�_bJ?�Ii�FEך��3h���=x���}I/E3��S"�9o���~�t��������E\o�r�D{�Q���C�����\>֫���E�("\�����V��&hn�;��p0�����a��f':�d����W�L��z�CF ��N� Y%WBa�P�x���2k���&��<X5C�b��8'�L��xve�Ȓ���fό�)ئ��y�����g���&o�9v˟g�(a�Y�$����Sc�0+j�s�M���L�Y����iQ7��~R�
��Ȉ࿩�(D[�.;\|.�0zD�u����}��XW.46�S����)%
���Y�@�����:�WC1��q��+sI���E�b�Y�F��u�+@A��\�FO�&J���Vq��(2�3�������)���<cRfp���|z�i�H7�����\(b�V ���$ˢL��e``rr��2�iT��ُ��Mo�q�'
��O%�S@�<��=fFǛ�����}�Џ���l�d-'Ϻ[�N���;R'j?[�=hF�L:��h�
�v�?� �%�X�	2�Gd<����ٷ�{q�/Jd��U>޴xYq@����A��݇�
����Q	�EF�)�M�낚"�����R'O0�KA���#SU!Y��G��ȹ���w?�l���_�}�R��p��/*H���_b�*�����9�gk���L�B��˫��(_R�����l��݇�""g`��&<��د X��AkP���z�����w��ෂ��;�/{?�N������g�}f_~�_��
Q�������]g����k���>3���*To���`� ���������:+��cM}��k���G7�����*�������a����ٻb���@���S���nQ�ԓ��,�S} ���it� K���i��f���GI�c�!�߇/��{"�L��f��k=-�B�6ê��=$��}Pq��_^\�+�Z�o�g����u�d7(���qS����g\������z0�$�2;F�� K�ϊ�9��_'tq��6�pj�k�Ι޲��;������_~��c�h���7��.������gM��E&�qe9sͩ�$3U��i���<30���5���s�ݘ,��v}�ʮe��=و��_p1�����ģp�"
\F�L���
䎃(��ߌ�}0�`l�P@0
�A�Bʃ�!2�R�R�GU/�\>=�l� z{����.����X�a�H�����&���Z��?"�R<�.�  .��;�$�i!�׫�WP���GF'���M>����(Dl0)aI�Q
O=h(��yݼ��E�	�.{�[8��:�y��=�'JP���7�l�m��+�t�,��;��atmʍ\����Y������"������:o���e�ۿ�����s\��$QFR{�OԊ��@��ԌP���=�v>�|hH"p2��ų��6E���`�>�g�&��g'�\�\�ԗU��|1o$=9 �󹟅\¤ՕekR�:S{�C��8D����1)��qb�GF0�����ի�w�>�8�0�<�v�%�Qs3��&Wdj��^�HC�XS$ZX�%��h!���O���ۜ�^{�S�.��mR�é�_�/:Bɴ�ԀU���Lz?�뮋����$��[dƊ�nd����{qߣm5�%*b��T�|`��V�\k�J;����UO�Ea�v��Ing�|ꎻ�R�lĝek��0=kkO���w�@g8�A��:��Ӥ��S�t<�26"�ڣk�5� c~�w��x _�g����52x	Ze��ڎS$�ޛ�"j�p ��k��},��YQ��Yʼƾ��Ђ�yź�[�b]\����L�`��������=_���苅��Rezru��)��cuΑ�]�!�_/ao͜	�ʃ '٭�$ϔ{mԪ�Xb� ����v;����0�$� cc뤳Qªhr0��B����a�������5w��~� �����E�oms~&�WuG�n/���
z�^��]Rj)��'f��N�A&j���Q�v���{���`��/.�f�������A�
�6��?�{�fl�N��W/�B�{ׇXS�B���������~�_2�vy}a_��U�;���ŕ�z�+2/�j"hq`6xW�wn�@>~�P}�=?��8d��+( �t
}�I���*s��;Llv�z�=�?�>���t���sȩv��nᧂ�o{(z�E�7�C�AV{��s-y�	���[�3g�l(�cѶ�Gf{��8(�S�"������5�'���8���yH[[_��jui�����v~� �l�Q���o��r�Û���x�QN��2��4F�h����J���c�YE����x�»)�E~�־��_����?۷�^�YG��>o�e�nj;�r8-��,�2���/��O|�v�����A8�1���v�~����3r�V̠ ���FG'P���:'.Ħ�A��H�ޅ}�1��Ը��#�>��l%⤿���a��>k�NGQ��T������*�fo�W����b��7i4xLZE�)^�f��G<��:�V�^� �X=k��^��=�q������Qubl�L�_f��-%zElٜ�Yf��Y�I]J���
zQ����[�!����N����?�ę��tB s=~���	�Y��t�׶(���K?2K�[~���L�/���2oƓ���� �*�����"Ŷ�8Ӎ�ԍ�z�9j���|���,ƛ h@���ZjY;�@ȉ��+�0��3�p�Lү'�N��Sú��5�������D9p��}���9\���:��4���托<�.`&��l��G��b1/�y�DA}�gu;E����6'��<Cw���u�uj���v���e�;6�Q�����J�m+b-�Ż�/w��c�׷����@����A����2�|/�h��\�k�,�b��95[�ki�GN�m��wek2�y7 ���lkxo�{�es=z���в��_�u'kj�_cL\�M���:L�nJ`�<;ш((I)�5\��bh �ʻ��cv� �����I�^�Yτ��%��!MV�P'
�ћ�[�Jx��J�R����n���O��Ȅ\UG���}��k:�8�ޔ�>5=�X#V��a��7̄(`�s�@1{�����?��gގJ��7N��,s�!jZKҡL�k��5+?���j�I�I�= V[pa�|�y&�ȶ5
$3r�%'z��@�������ϫ�g�3K�P��Ɏ����\C�4Տ@��3{a�W۶gއT��p�W_"1p��Ძ_:^���e�ΞuRP�z������iL����`[F[ԣ�χ���H�������}w�:�k��o���_}V��3K&�JPڑ�½�����fd��h`=������F�Z��qQ��$&�S�|��j��5�3w�G�����?@gU�+W�t;@�h�Zy?4�J�;(�۽S�����0���vF`{�s��:'֘�˘���!�d�,��O����\�z�=d�w+W4�����^/���՗��⊦P^W������W���B(WQ�;�q]+� !�!6�� �ȋ;�֡D� ��*�{�w'�e�hA��i�f��>���A����
���������ۿ���������;������,(]��٢V$���wo�ǚu�V��^�=��1wp"���p��i��_���9�#��P�� ����<���M�yƶ@��� �C�H�s�����1�����CʊBNǬz%D��q?Qͯ��ۂ�}V����=�_]N���p]^<s��ںぜ���`j\O�;U��R�Q�#2Pj��cN�������)^}����0z��$f?xp�{�O�N��p #� �����L]��\�Q��*\���c�!]:m�1��kS1q�5-�U,� "i�|��lY���Xe���+���o��@�lC+�c|���e�����'{UW,�Z�ՅF�lv�S���[�1ڙ�����65���:f��*]S��� ҵ^`�>�Y�Hk"91�E24�Xc,�:�r��v�����Τ~1�-J�`1;�9��a�#�dН�L�|v ��3藓�+[����4۩��g9T���s���4��X8�9vk�� �/��N϶�}���SN_T:[�t���]�(����C*��/lu��H���@sR�M�ۜ���u^#@� �y���.z�]�:Π�f��� �b�'?r"�פ({g���8/�ח��f��[����縈��!�,����5�I_G]���;g�����7���2HW�ѷ�qD.B��t͡@e�ܗ)���U�!�]���lSb�ND̢EMl���G9*3"��t��?��;�gǎ*�Т�l�H#�k��E�ۀ���^�~EV�mvՙE���>d���Çw�����c�-���ō�W������X��Շ��X���f��ғӐ���TÞ7Ɩ'NV��U5=�.%�i�×�}�y3W�s ۅ�K�q�ݙ<���5�>F��U2��}�*�\mΘM��ϛ��u��b�T7�@s�@�a]X\���X,��C��v=�X��᪔O�3"y�V\���!D�gk�+��@8;Ә���m?�����i�6J�{��n�Qwg������ �;[k�F�ώi'mofz�p�
w�X��1�k>����c�E�]������v�L�+f��-E= �{���m�x՟ @���>�+���v��f{;/uȹ��`��>oV����L����>�/��$G���7�{9���|\��Q�
`��@�'�W$���}G=&2�����e}����X�e'�$�������J��A�Yf4����Y��4#�N�8 f�B�ΕŁ*W�*CA��ݽ�������������e���?���7��%�[q]:��^��4S��2Y�xv�=��vD�g�������8g�.扟��a����<$s�`rQ����{	Oj��!J>�Sԫ�k�"��.�*V�F�8)d�IԎ�}3�`S�$�qh�{>�O>PB�]ls��뻧� ����a��zP<�?չ|d�_��c5��Z�,���u:���EFZ��R���N46o�� {�T��G�5"|{D/C���u����|m��Q�ByEF�0�V��hݰX?K�5�{q�e��.����'�C�2.C�i���&
�Ǻ��3��n�����?�Ϝ��c�u��s��=t�[�������)�~�G��H(�G�#SS%Au�9�@����a�{�y`��r�UA����C�p�`�����Y�C���@�x����ί�75@��Jd�"��xhqK[V>�a.��q�Y>'�H�s7�	U���e��@��M��`��.���rI�.Ϭ�g��@�&�c1_� a���)��7�ש��7qMq�KV=|9����|�ӬkP����SW�	K���u˪9�Y�y�m�Kr/��9�W\�%3h����y:�O-��PI�۵D���[����Ѱ;ʅ���9H�e泼�����s(�����}��PQA:./��;o3
@d}�I��A	~��ft�rd��^ԛj�F�9��Sqg_�=)(No����fMY��'��}�M�k�ּ�
���� XN���1̚���~d�3��=��9��~�R�)��#�)���������T\�Tc'cB%����O��������s�Q./\cR~?N!���6L�=�jc�dE-%��7�E4�l}�0Ł�Ȣϙu4�Y��~Q3g^�Z�G���3L��>6���S{�g�/.o��]��%��Ա�?U��+����{�O͞��|��x 0[}�����^R�+� i����9�$��р����,?輞���̙�ԩ�6ADn���!SAR�p>���2��%�Z�2�Ǳ�-(��|
�l	�j��Y����H�p�h��5V=X<�� C���z˺��>�\u�G��d�Ba`�><>خ� '��9j�����lE�==�")����x$XIQ�}���F�B?����z�{{x�<� a�~b
J�	��]���=�W�����tm�� i�/hAQ�������K���3���!�S���5�(���)��\�N$	_h:zm@�+X�8��ar�+-Ξ�H�����M��6Ӣ�=���7]�TD�9�������h���=G*
�y�޾�����KFj6�s�d�wh�(��$o5���4R8U�S(~4Q-\�$�^�+��O�-�x�ɅJ8�ij ���XD�c�YּB|�8L�����NŎ9oI��M ���?K���+�<� 9�ڔq�`�+�̰w	 o��N8��$Qm-�b���:��?#��h�v����BO�Q�=���l7[J�tS����
��T��۠^)|C��]����ٓ����GI�����%F�/��*��rNt5��=���Sݔ��/�<h`(�D.�:X��%xa��Ҏ�K�=������9s��=Za
5�\����)px���;��0S!�d�,	�=�XƼ֊~^k�ז�D�+��?7�*��&]8���&HZ᪆Kw�e���C�/\��zcV�Y3��U�t/3��nam�`WJx��M�C�n��KG:z��iX�u(��e���.w"��Z�Y�8$���z��̼"J;T#Ki���z��� Y�e��z����0��ay`��} �O_����	���T}�gw�Rs�5�8�׍rЯE*.�wm��.�����7ާ���7���Ӟt�pee�P��]����LkQ"2)]�͞���g.ʁA|A grbT�E6,Q�N�1j]�b]�5�(QS$����T��Ia`ռ��5c��n�y�"�~�ژt"����rb蜪���j ��k�uEhU�Jk��w�� �w�<���|��,���Q0�ΐ-?�o�Ν6:�A�4�}$2���QY�Qv�裸���N���m�F��ʷ��$=��$(��bN�A;d���#p�h�a� ������(�pzo���:t+2k:"�Śܺ��`��	<)��Z/8�I������G���ƃi�m��y 32��������>�5X�Q�(�Pԛ���
���R�R�A��� 06#?'K�)+�K-8]X3�3�WU�=��#�z�I��B0�51c�,��)j��U���慿?]�M�);�59/o^U�p`m�9R�����u��{��u�Ի�YW�$��W�P_�D:�<�hS$r�� �������}T��z�S�{��j&�eɡ)�W�����f�si_�&*����+؄��{���l���t^�Bo���>�'�{��/_���[mW�K�]FO{���d���E6�:�)ؖm���k�����5N"c�2�R?F��N�A-�&���1�@�*(s���=xבŅW8���F��B)԰����S��d��#yy����q��8�+�s'�'@�+|�|�%��^�ʽ����3����_�utA���
��z��	�p6>��X)���3���,wa������ɳ�%�Ea� �5�
p�0N�b�Ա^M+�����fC�;��v�.��X*`�J�ս�'ݏ=
�\ُ�YE��d�mS(~^�U�5�#Vb�E�,�p�?!2��ak���G�#l�0<P��,��bć��Ϊ�~{�fФ�Nk�̂���I�PQ�?ԁ����O�"ÌR���f��ƿ��
�6X\��Ц�W�T�W��fd�G$�|N����K�|�ǯ�^������s����l�"���ұ�X&>��6
q!�kZ��^�R�N	���I�y�:��u�8�4��yu^܏�i���sĪ��;�s�9w�J�69o_�R_$3ϣ��G2���� MIuɮ*8����bo��k��H���?��>�I�v;��=�V���O��v�]]���Ņ6`��aw���r��̲	�B�^%��~�H�bP�f��q��A�N�䄗��\2�4���rJ�o�'K��>��������֐�n�`W�%���{�5��cp��=}�����>z�G�>��%�O�$��s׹|��~��kfQ�O�m��9�y�J��izH6�oE�T\������
�bo�ͨ�������e�67u��C�#3�̻y�"�����9��6쳻�e���Aj�@�����1�{^��\x��mg_;PK�ց�������J���j��=:�IT���pۅ��(JQ�W��xv�xY�+Y~����x���;Ԩz���%�X�,vI����	�Ȭ���|p�9g�ؐ�3�ѷҲ���	�B�}��+^��)��Rd�����n3H�z�C��9���8� Ӹ�����,"�C/��A	[��??GˀȨ�#|��E��R⡀� q=e�;��@ .�꾋D<��y�.��ѷ��7Pt�-J����9�{lԟ��6���$�#>o̓׏�����U"Ö�9F�!0'BI��l�>Q_;����?<�+�m�((�Z��<�ֵRp9��@�s�&q?�/��΀��ԘE�((RgBGzk��+�  lWa�T�����ϒrb0�M�|��Y�����h��>FN���{���P��h
�:%���� &���ɶ%IɷS�ω�����|�sh{��7o�l���û���\��߼����K��Wv~u�o��a�Y��#���q��`2�+���� �����;�*#��5x Dx 0AB���� `�����.�l%DH�T��A�����L�#�}� |2�ճ&�] kO0�H!�����Mj� <{���+.��p\u=�\�8Ӑ%B�s���ת���#87noo���ZMB�߇�����G
k��*�=�Y�>�<�^��d7��^��dAT�
EM��l<@ k%+ ;���]�\��׸����j� eP�0�R��l���20pۅ�ڊ���3W�Zh�z2�L��0;����{�ߔ�iwG�-h��`'A����R���z9g����43�u��]%��ĝ�������{$��ם:@ 3ws�f׮��4>>)��E~^3k/�}�zswK����U�]þ�si���"W�ȐcERqB��S�ր��X��)�Ĉ�lA�e��TG�M�$Tt�A��ψ(��lmo�6��B^w�#�C��Z���\{�8�r�}�w0��5_%�����ꅄ���Gl��a��v'_I|��U�-wl�G͉ӍD�r��1�*�瘍JFG�k��ёMΑ�������+8�$��1��a�У'�P�	q�ЯCVuS��dC��9�3�Λ���l�f���y�)��w�����>�V3e�A)֐Ȼ]uWܠq�#�Ri[��	�|�z�E--�$M�،5F%8�����8R@�F��9qGm�����Kɟ��p��Iiڼ�	W����z�;Ъ�H�T)��~���~�r%Id�R��S��Fם��׾~_û�;����sPT���1*�������v�}pM�-���ޓ?��+u��hD(WM��σH�̢}^܎�o�6=Ԑ�}g�g����Ժ�򛮓�L\�J�t��
�Šy6R���ƥD8\��YO���=��i&P벚�ޫ��iLhg7�t�*�gi���iSf����X��F8}���S��ӓ>��2j�����i�s }Q\�� ����-*��Ɠf��my�dl��r�9��J���^]�N��zM�â3YD��S�����^��b����N:�©8	�V ����Z��c��=Ef��Pկ/�S_
ԓ��T����K`�>uD�7��<&�Z t������P�L�LL��h����AP��TIj75H'��5�5bd9z��HURҌ���K���e*k�V�%R��9�iMN��A"2��\Ey�*3���=
u���\Y	��ɴ1��@adT���N�+�_Mo�j'�`��@��0��0Vʍ=�d��|�^[��z���ݽK�u��@m�!dM�j��2K�=ِ��{\?x�O�Ni�z�z�
X��.ҹhm�S�����ZdR�y���8�+��AK�T�>����ͻd�QG�xft_��Ԓ�t�ƪ�F������х\��=�8�?�ȧO'r��CJ����f�( Y軶Zh�YG6�ǅfƣf����	�G�p��\����l�lN��v����d|nkg�6�6
 �J�m��"p���A��`S M	Z��xuA P����Ņf�a�H��x�Tؘ.^`d\�{�e�a0���p <Ȧ޼yC���H�:mp��Ji���\��������?�@nks�b���R8d�{���t&��{:���(�em��@}K��Y�7A�3n���|� b����;$����ܥ���hʍ���D��叜��t�Ol�̒���e�X�3���_ӓS⒨jr��,-l�7������f���ށ!2����2����3YaLo,l�ٲQ�W��� ����42U{�4���Q��q�L�D��V��4�kQ�X<�4�u���aV�rҐծX�fX�h����*Zm�Z�X��i���cS@�����iA��>�v��ǿ;�4��D4*I4�2���s�[Y�'Z�c#�%�c�q���*��3O�3��y�"ԠR=" j�Ⱦ@䶳�/��}0��	#��|/��<����첕�i�//��R6h;cP�����f������t��&􀞔/x�Z�gDG�P�� 'uEY{���������7F�a�k��0ҿP�^X�t�F�f��A��RP����������]�A�����B�T�2��I
k�P��@�H�e���?��i��'~~��z�Pޗ|�8�^S&嘵ND�Iu��A��A�Z�Sm����a�s�>�f'[[�M�����$g{nS�����^l��z��i$�l�MD���؜r�����OY,�=�JG1{�ʓ�k,�?χ�	�X޾sH���\޽{+?������F�&�N�f:t=Î�?˽������r��>�G����9x�����r>e6�?�{�$c 4�<�q{�ƅ1��o��~��=y��!�1�]�J�����\]\�Pd�& �އ����Ǐ�x���)�����OK�.6����و�2ӟ��M�4��={�]���E?�R��i�>���J=�T�E4Z� �� T��l�=E����1�6��W�������|�NJ��#�?}ѩj�Q�}s�-���H�m�M���H�s��S��0�T(�HU�
�� �J�ä�6c:��w8��f�:s�����Z�@BT�+�G�88���ck�4�T��ߺ�(l
�馊C ��/�R,t�OFdhh���������,���P�VyNjR<�+��Ȃ������]\j��[��h4n$����`�O�{�t&Gt`?}�Ox6^C�y"�x#἖��ͷ{�ƱO�f�t5H�<@�����&3)���b	�A@�IZ�9��6L��2���!C�σ��;�k�����t)��3ZxN��l�>1C	ьYC=��`�jG)�`�,��N���mn*5@G�#΋��ҳ����(�{-��*}&�.��d���y�]*������V���Q#��3�R	u����R��\�����Z@Ń�eu=`X�'&�"b�"#s�������f�kn4����'hH���6%�D���+BF��P�U\��kE����N�6���Q���F��;����J/F�0�R����~�t�M����"ϑ��˼�*Y�������V_�<��qH�-Op|�]�=� ���d����;�c�-Ua�-Qb�3�H�:�pζ:&�7BΑ��^��rO��MT%H����I��}.j*�*9y��\��iGV���y�S)⑗ꄔ������w�g[���gqG�(j(Y�G���`q���t�f���Qu7G`����� �@���5+��T��"}�U�B���%���mC�A�,8fX����NT>���X�qՖy�̚��_��m�wNy�0��l�.�K:8���"���X����Yν��{{K�"�����#Z�F���A�	���yCRud�7.�N��Tӑ:�6(Ѯ�C�.VCQT�R�(�L� �H����W��U�Qv�~@�"�we=�q�-�W��ip�k�v�b������#x������Lyj�,��9��4���n���wC���r�'ĭ_�p�15��h�О�zf��.�uS�(��5V�����|�z�ra=iJ�~ ݹ�����x�|�,D��i�p}}��і�W�����Cy��K����|����;�9��+}����)k}e
bq-j~O������sw����\I�������-:�P`�?�^e���d��Ų3p�f�p�*�~�&��?����}`��V����:����Ȁ��������?�;��U�ļQ	�<�N��ҐX�Uiu�$k���� f1�Ĭ���7웲�e��X�q�e ���������XƩ�&Yn���>��N�cF��O���A~��<���Fv6�x�x�^9F�)$4��8��y��ky��{��D7�Pקc#����m��N�-d��N6o�٤���ӧ#^���#x��sfn�g���yT/]�;�sO�箲�2g&�7p
����a�.�<٠c{yy�V/}�5��Q����n��hFnG;��>=�绷��ux��޼~ÞR�YOA�����N���t�,A^S]��6����aW�Uq�W*6Z3�w�+�cz���0.ю�  _��ze7�"�J�$�m� ��T3�Y��0*Z��W%i/Ju��N)�tӨ��k�ng
o.��M7��OI�7bCٸ���\=�=�����ܻ��X	5��u��x�V�Q�zL�3�gf��3���l��͇	ֶE�hVM�LwP<$pn 8��'�T�Y^��Z��u�m�u}�i�B��'���������{c�����RTf�W/�o]@�X���U2ap��e5cDf�\��^'�y�PT��@��rU�{��sh�my����-�>�МmO������B&�#�U��� �Keq���r:>��&{�.�T��i���gk7GcW�9j�A��ft�sD���n�u
+�qT���
.DG2�^v�
��X�8J�~W��� ^C��P�ױ�����د����9��:�$-,]��c�a��R"��44tvRg�(��-*�c3�0�f���}���ɛ�-^�{�J;٨��csvzI���r�@��L{S��s��x�do�d�hIZ�*�
��ҋ���U�����UK��Ɋ!��ԟ��ҫ�:�c���4h=�zbA6��M�?]p���?��z��5%�X����{�h�ţ���hP\@@��U�Q��X�=P��Mq�(�Ƽ�5P�/耵�+�;����Bvo�	rƭe�������,+��:��nx�
a`u �'*�2���Q�]��Y��p��HD�J�*Z�r��
%s�;�'_d��Ņ�'�
0J@���x�LמF�s�()��x���'��M��F�+����A�����O�C;�h��8����Rk!�Z����mJhF�Z�{�7liG)ں^�Q*���f�*�H��)R��$V���6<�3��8��@��h{K�Y�o��ƕ��6����Ƞҗ_~)_>�Bnݺ)?��R..����.�����u��R_j5=pZo��>z�ǆ}��i �������3ж�u��}y���p��,��s�_�h\����C�}x��/�c5��`���+9>9��٣Ц���V�� c��pƑ�w�<~�H>{�T�>y�y�㞝�|?��p������w� �f�y���_���|�����\��4Uϣ�#�r�W�|��u��ֳ��Q�d��v4j���֨GY���Xv�wV��c�,@��Wo�(���ʁ;�تCd�K,���qeRĞ�ؘl˃{��ϟ�g�=����,7aJg��{�����2�?��}g�" �o��^^g@0���d0�(�A�|>�����{pW�>}"��O�3�w����:F'''<>��p ��PF�- }�7dp�b08;�����<��'y��c���w�Oک��n�s���7����0�=}��������
��5� ��G�*\���%���P����ٗ���Y����G�3j	L���Һ)qg�݊1��1i�T���ԍ�ң�HT'Xa�2��A4�	 ��3�1�72���ɲbvJ�9��i��M�x[**@K�<��X��Y��/`��"��* �ƁR�`� ��	��\Ԭ"��N�-M�Ȳ
)��x��J�}T���'��E�KP9��}���3߬6T'�T����i]��V!�E�璟W0������_�`��Zh���N��,hmZ��L8�˕�s]�-
 oFk��,�������%k�T,��� ��B�\.�`+^��U�n��}_�l7Pl��O�>+��}��~e5��̧h���nG�R d�`W��S��ڷ�`��E����O��_۫x�Z��a��کl�t�Q�m^c("���h�I��K�+��i�b��|T��@��"g�d,�1q=����lªS-���;d��S�J�`R�,�h�����p�`�{0%W	��{��e;�ғИ΂��z�����HqTN��~M��f��4���p4���E��r@U��i��X���&4#�i�SUw�������'fr��,;�dp���՝�Z��|�T��;�C�ѯ#�����k���w�i���`0��您�j�	�B�zY�:!#�̩6\�k��������I٫J�m�(��"Y�O�ͧ��vGe�>�E]� P*k��O�9��� o��~ٳ�F3������i�eg��dL\�c����fK襢���i=U �}��J12&�R�}��d+�G���M�{��Ō�(k��K6�]�:T��:�lV @⿋;b|������>�~6c�g�T:/z)�*U���q
�����w�&�`N�|�@C�����t��������K��\7~7��R�H)qi��]X;!�ޤD�!��(��@�)s��z_�
ʭW�Ƙ��qas@g��j��~p]���g�jyBI����3U{�Lփ���B��ۑ՞����>���[�R.רO��L,S 't�f:Un���nnl�������𚨆E�5���ϯ(�{�MyD�5i���3��wxx(ϟ� /|I�5�:�x>���y�d�y O���_�: Z��� �N=΃k��+������1h��	��ׯ䇗/	(.f�+��e��?o�>��!�h���{k�j��lѫ��6�U��x0.����|?{�y�O�o=�"�q��1���R淇\%�
���#���oF�{�n���׿�Uԟ�
����g�	����!��c>��s�u���^�̀�-�}tt���*�ìP�����˃�����_��+ �)��>7��a/�}xK�y��I�Ԫ�]�F3�7X秧���s�|�p&/^�$�۟�u���FY���M��'���C�/�5���������yv�d��C���Xr����j 웘��Q"}��]��G�[�~n�y�����^4"�{Ӏ�֞���*��%.�Ԙ���(��OL%��aP���!ZǸ��y��d%�S}"m[�
��>��V�#�K�*�9Gc@Y�4ɉX�(���h=�v�[ �WG�+g�_�
�
G��f�粘_�߫?��&ehз��-U}ԡΜ�@��h���"x~����YeR��d�-җ�6}%��k�����^���t�j]�K�J��G�>K��t��^E� �H��}�������M���'�_T!t������Oe=��K��?mS�M�E9����ދ�a�҈�dƕ������yf�����Bړ�� �����d���� [*)V6�6�"��4�HUF���n���S�)mSԴc����֔d@0ShtJ��
t���h�u�{�ܨ/�݇�aG�NUK,�
q�=�i^����d��~��T4���-��e�VЙp�YCh"q\�Bf�����&?t�|���`�Nű<�h��5-��
R�x�����/=�V���і���	# 85���Vd���u굹��9�$+�/��c�_v��uR���.wj����	��1na8V��0vz�-qg�U%_���-o�Q�}Ț���[{�� 1��4T��` �F҅)����8X]��I�V
�"�Ϛ/�K���eV�	%��8�pN,���d�3 ��8ώ�q��w����s�l�s���{�o�B�/л`����6��z�
��E�;�ܑ����8;� `(�mL�ިA��({�5�8�"�(ASI2\)���"e(���c���K��oR����<�99|������~t����vI��'�c�+'2�Y����}��Ȉv�a��xc��v� k�O
E8F���R=�}e�ӺDˊAc0�7J���B` T@cp><� �Y�]���3U���u�[��Y�s�k��������x4�yd�5��0[:)]�$�`�ͻ6��iT5�b�i15\�tk�W�3�Ԓ=px��ٖ[�������.N���&���/���iV';o��u���@�Ì�����P�.�zJ$�:Ɵ�!y�߾};����<�G����ƺ�y]��k\i�t��&����S�_��q�e���e�����[9���~������5XRk�zS5�3 *�:��J$��Vy�B�]�;�G��g�}ά⣇�2(�%U4��~zN��d KHQQP�kO���΍�w���6Ǟ<y(Ͼ����������\�-H�����9=��P<�h��&�w�v2���o7�ﾗ>0;`՚��4?�;���ٳ���~����G$Wo�J�{����@xf�/	���o�6S�$|](�jw���TrC�����D�-�ؖg�?�@�<�v	J6&9�xC^�˻w�^�1�rX3f�Pt�Я&(�X�5Iv�'m^�An�����"h��A����+h���c2�~�RQ����>��ZfEt�z��`��^�b}��J�VK�(�9�O(��9P2|9��{k��b{�T?�v�o�41��+d�Y���7��Su�� 4X��_�ڦ1c%�`kF[7#�!�54'��̘5�]�gॲ�}���K��&�K��nI�6��8&һ���2y��{D�N�D���b
���.���{ً����/�P0&���,����=��/2z݃��U�*��;K��]S1�m0YͦQ~鈛
%��ɕCZ|�(�0.�Ds��}��
�V����+��Qkt3���npM�᭍��* Q�-2�')�
�WA�U�Q:N�e㊚�
L��xT�}���rYd"�DY��R���������,���|P�<���Xj9���8!�b B���l�ͱF�$p
Y�0ጕf&Ti�m��پ�.���<��yM�'V��@*��w$�c���*�(굷L#�S3N�E��#6���D�k��N��Vʅ�U��f��9�,��I�&���M'���1��j�\Ң�ޔD���c�s�t(w�+(tGRꅭ}��6�ʭ����>Qe�+�ұ��+rM���B`{`��c58}q xw}y�"|�-�	�ɡ�
� �b�кfj��Z��L��T�^նlr;���<D��v��(�
L]&�dac_u���E�}޵�2w�u6�Q�yވ/�)�fg4>L~L�.g�Zd-�^@���"�6��o�|[f��V�{�2A-p�%k��4���;�LClQq�m^�&�Y��Lҵɬ.oW'��}!���P1�9ԕ&��F*x%�uN��~��6X��	2?'kҁ��ae�0�g��0y8�k�\�[��[�j�?��Ή���f��Yt	5��^dؔ-+D
�T�/�d{�c8�p����i��2�𫱊�,=��� 4`ĦJ6����MS�����ԧj[sP�x�M�9�m���=H#f�Ԓ[�:� �B{� �J	�z�J�� I #_=�Z>z$�nP����f���t�(P���Ͼ������9��2':2� ��;(zf�'_��7/yЖf�=������
`�3��g��fJ��57 ;�#�y�ɢc�P����C\�e{{�G�dg+;�4�Kfj����� ��H�
�x"}(���\j�b_��)�J�j��;���W_?�/��L�>��Y,��M�iv�?f`���ʿ3�sfl��U}`tL8�2�}����`�~>�|.�Vn��ވ��b� )�D���� �-����i"�A�w�Y���e/�п��*k��uw������W_1��~7���b���}�'�.�����.�&�A��c���Rt�Ț*�	5rcwGv�o䱈rzr.�["{��g������<~p(Of��4��lO~�����6�i:�j�Y>��9�0�ex��~��<��<�s�A����ڇX�́L�������|.�8���@oϿ��X� 2+	�*}۶�h[z�D
�Dzp�ِX��j�j�����r?K�D ���N_.l�E�L��! b��P1`��X�4S��KW�*�^��{�g�aW��C��(	�)
1��!Uz,3d�.��E-����sX�CQ�
��H� �X��+���l����� ��Q��ƕ�,WyU��b8���cpӶ�o��{H��\�#:X�9�,�,�Y��og�FyNc��[��!����gqڵ���-? Y�M����֟�cn�.��.�3��T�ه^z��Xo��>Ҥ�����3!�ꗤX�/��4���=��}Uꔬut�ǚ���(25�#(��.�'��z4ꓩ`��.\�5F�퇕���8(�Q��1��ۜ�m�a���&�=P�"9�~3i�����i�D�)���>�2qb`|e4إ��t�꧳���֋�Hǹ�֜n�3�)T�*��Q2B�Uq�����C�|�E�~Gc�M�����[)��m�t���ڱD���ѵ��/�F�iz�R��͐����B��綊�i�ȵ�W&eE�k�$���4���Ru�ʵX�"���4�x(Z��J�,���y�[`	-W������R�
�$��Z�r��,�gݛ�SjV�`ײh��7�ȸ�;�,"��𢶋�
?�+99�b����	#�0�І���B$�������-G����ƨ�R�v��F0Cc�I#F:�qv�V��`���6ø�N#w�4����!|��!�@Cx��^a8�g���z6?ro;�P���u}]ZA������]gu(�O���.�~��*t���|X{����)�^��}Xd�}�������,�`��:lI3Y&P�"g�cQBIV,��Y�`�~
����!C���)o��d�������21[3ך,��*��?�7�7 =�\����&|�����X�>XF��{Uʹ>7T�R�ad�2��{�3;(���ǽ ����N�<}���M���Ņ}:b�U������0�;��*��_�fd{�  92&����K��_^P���"�%P�A�Ǐ�7���|���O!��|҆Ľ��ӧ����C���OD�Q��`�8��+F�lb�Ԓ��N��J�r�3���Ylg�Һ��(ͨ�����Y��o�ٳ�����[~�r>�sj¯�-Qm�l�v6�m��T:������~+_}��uky��� P�l@�v��^���J+Eu���g0Z����&��[72��0�����7��.��J��`��<}�(��ۼ��R�V�)M�} �������[�/ "Ag-e������,������{9=>����ٿ�#7ol�V6� ��ڿ�A��y~gК�p�I���H9�qX6p�������B��nȃ;��g����;��:���<ov�d;�avV�&��=ʫ;j�9�>���ץ�IQ�ThEl]:�̳d��fw-8��٩
����aO:qX/�
��ig^ۈ`5^X�4�B���cR��T��lt��N���{��͠G��A��3p�
|}rZ�։��=�������\���6�����q��?8��m���M�@�h����31��02��fH�v�l���A�����=!&S
���;e�h�
�D�<P?G[0��βC}��΃1�,h�NJvQ�A>���Gh�{���ձ�YA/e�@k4@�R=�y�����pK�tY}Vl|TޞY�N��XY�@O�1�v����w�T�hͼT)u��SkB�id��T�Õ({�7�Z���.|�g]��d	�^�m�,�@-��j(�D���P��$��7�]DN�2��	��6�+΅``}p
vĶ$�<`W��y-�����T#�-�:i�.ț�L%+�c3��,�F�b��|@gi�+*u�+L�W��Q~�JF����a]��w�|!}6���B׼9��y�����G��	7j����C�%f�
���Ct�~�![��lI'a��e���B��FT4��A4:<p8�@��R��y��)O�!�	�jM��Q��:p����Quy]�%����Uc�)���;dҳY�q��A�E~F��iT���7�L/��ی��� �?c����� s�h��	�%F�V}�J����%�-��R��� �ǉ����,~��1��]^GY ,f#:@Y@�%}�
�	Ȏ�,�l���d�;��K�ʶd�?M�P��LfJg���5ht(�8�e
���B���GT��
<������$�X������;�:9�D��+f����UKe����:���@��E�I�J@PqB�Jw����.x�uE<~?�s��!�$*�_{��&M�<�,c:V[��v��"A�ja �^��!¨k4�$W���&��R�zk�$�[�+Tݩgs�{[�ݣS;�Ц�}7��&�����>�=�u�-���� ($��t���Qv�w�3��[%Sp��=��N�훇r;�����dA@ �Mv�x.dhCTDG�y=�����d[���ݝ-m<�:����w7��;/��e��ѣ����SJ����t�%��e�R.ON���{y��޿�>[X�����)�g[����;w9� V Z��i���eA��Ç��ݛW�مE�	���'���N���$�����V��zV����[~�ŋ�ى�H������1n����Y~Z���_��C��{v/���#��?�t`�ػc��|B���l)���3e�^��gh�`\��d̓'��ɿ��o䷿�F�?�����ee�[ڛX��*�gt�"���ʄ�0Ǿ����??�����싇 �Π2���ͯ�ܺX�G�FK�Jfq�)2�q/&�]�Q?�?2U���z"7�3��hd��?<�N�Rv��ѝ[r� ����F`hA��j޳0}vճ6w��y�����ܘ�4c����}q��I�֦�����[�ӟ�,���������<��������� ��2�0�n>��ގܿ����<�^���	�2���}�L|F���|�y=�wO�̀�~��6�e͐?;�����������I"�wq9�zűQ�z}b�d�F���>�8���J#�ԗ�#j}Wb�l�2hy���<��Q�\��R�U���mp갈"�S)�Zt&u�{�@:�y��S���l�<�s����J�VdqzF1���΋Q�����g�g���إ)7*����-E��a|9�&��� ���v*�Nk��/FIbm��F�+S.�8�
k8
�D�xos-B��/�(��lŽhɀ��db�A�B���f�g�VRĜJ Dt���]K(�˛�������i�B��论������L1�T�ĝ��AlfU�.Z7�8 w��+�T�� D��f�@+�T��h����FF�gQ��j��I��� �%<�e6UNP�TTj��W0�`�CW iǾx*� ���DH�q�QT��.����p�4�7O�F�?d�1��L����X���h��������/�	�O�Y�9Z��/}\ג�,���X]Y$��ٷi�i�6~2L'��<��\|q��)�/�d����#+uA?�?ȧ�O�Dn�h�
|��0k��Ǽy����>eM;�p����а@���|h_6ϴ�!�k��q�;9
 �Ψ�	��Q��}Q�X�jG^�_�_[J6����9����k�yK�{>��6�>jQ#TX:�ť�r�g<R�� ��z��� 3������璋q�amS�ƭv^7����sFz���{skJ�(M��Ĩ���9��;�e#yz6��Ѝ��U�̫��S�K���"�p�K��=�A��MJ�o�`�J����Ͽ���'[>�D85b��65ji�'���<��sN���f�<�d��i�0I���u�5���R�h��ֲJ�>O��'��^[BZtk���Lv.�C��8�E]y� ���jc]�pE�mQ�^�(%284!�*V�M�88H�@��t�&�l3҈����trz��[��5�F��b�pc���2q�̞;]L�n2�i���\CJucʯIk���T6�M5�8�_�[cM��Z��R�Gɛ7��L������xܾ��E+m{co��M��legwJ�C6��4־U���궿�Js,%���H�~������W������߽z��A��-*�u�HV�1�d���0�P���\�..9��N,x��i�����Ap�k�掍ʻ%KT]r;��}*#>|����h�n��h�q6Q�5��n� -�i��uR�1d�ng���7��~�+����r�ޝ���S�r���Qu����J ȚN�L%��y���
��7�ܿG���� x���)���`�����dJ���-�c��&��xL���4ḇ�"�����&�|�)�����^������ǿ������\+�}_"�;�����62O��B�ֵ�,�f�{��� 5�RǴ/3Ć��wz2��_�y1�2πYmÕN{�`hwx���fm�^e�O���u�L>�ź��A�tFV�\d�������LSmT�^>:��Pe@���qr�^��vU����B�Z�F�[[9=���W���K%\��T�:l1�?\uLגIceT�3j�g�8�A��X0j��K�ic�B�LZ��BJ�#8�\����k�yW��;����^h�_2ۆXv�_UѰ贈~�ձ�h�ө�l��MtFhl���ӟfԁœ$��Z<��2+��	�(w��C�R2��Y��(
�G-��}��:��۸����%1�E�ߛ�]�T�	�&��dĩ���3A<S�������NI���P�6F����S�̬cӉ�`���{�b�\!+��~���CT:g�^e�I�Ϸ���X곂��#�d��g޼N:��&��֝uFꍪ'�5��A�D��{h��D#���0Ң��(�{y���
��t�7n���#r��驔2�6G�\Y9mY ��4�v�x�`��:Ǥ +��q�x?v�!��H��\����������k�
���ʹ���]�ۢ��b�?���(��?#���t:('!�o���7��ߣ� k�d�`���FQ�:�ԛ������$b;��"���/�È���آN/Z���R�\�3����rE��ټ������.��Ů؜Z۫"�,nLY�C��rQW����מa��*fgm: ��Z�Ð��3b�����j"D��|���yCl��2��i�y�O��n�ײqz���d0k}J�>`���Jd��5�L���5��Ն�`B�@ ����{g��}�^I|��_2�B�M��n}Z�+p !CΎ��0�g(�uK�����iTQ�y
�C���L\H�a��x9��1) 0kL���T�"�G���ߔ7���1U��<M��K��&R��:El������c���Լ�@Ë��Q�N��Qp -��j>�>V�WU���5Z;ecUGK��f�aB
(���T�U�">����^~|�R޾y��=�I%|����n�f��&��޼�����x{k�Y�����zA�S���H��^5(��Ea6�q/����d�]�/��:�ݥ��_|&_}���7Q�h����*�/_�@J�<�d.�Z��V��U�Ng�n2����}��9vwU�0���[���1�ha''��%�S~?h���1h��v�r�i��kC�dvw'���#�����O\��j.����gL��<����٬��|/Gr�����'��Za���lm��ֶ6N�蓵�¨��5�%ʿ�����3־N#k ��P�T��Gݗ����<�� z`q�!#��DE0ae,!����j���A?��w�D�3�0�g����z���ָ�6�M1����.�e����h���4T��@�5�Ȅ�=�Y�b��N�髕�j����F���j����E2���˾�L�����{c5����L�jW������`����t��vH��*d��SomĲlb�%s2�nL��)x��F���B�}6�G��mִ*Rd�m�*űU�c�`?Y�o�J��Y��@�[,��>Q�-jB}��l�,VU6)��0_�Ӡ��`�)7g�ޕާ5;/G{��w�G�H9�m��,��{M��%$�g�ւ��C�=hP�<oSdf?3���g�� � ����P�W�d:6�h�؈�-"��y�6���)��H�����d�L����D?:�2n�sZ����}R�#9���J������H0�@�6*��/���>��� k)-���ځc7����J�֣�E��?[m�]t�F������D6��?|��
�����r��=������/G�G H�X�Rr��}���<���$�?����a��O|��v}&e�9���_$� �7#��cY�~������4��U(|U��J#5d�l��=����U;W�!���ΊyWL�'K�:����x^�KW�!��){�QJ-_py���*�l(�7*YW�}C$=�"�H67Z�/8Dٿa�rx�C1ώ��lN��uu���K|��H�	�fӘ2��R��h*�����@�>0*�o��y��W�o���,�'qL��R�jx&�K��e9X{Z_d5vA�v����(7c�S�o9��T0�Y�`�����˽�:=t�P5�0Xc�>?����P�uWX[���h�5�G<`��_\w�P���y{�u��FD���Ԙ�n:׌Ak����_�w���&�o��V!��P.UҸmd=(x����lӐR��y�&��)�hE�
(��슎=������GA<c+��˛W/�ӧw2�8Q�\��KU��� ��8�z0�)��Ca��N�������BU`�,Y]�g�����/�˷�k������ρb"�6M~6��}y����2�ٺ}X;�f �g��#���"�SQ J��X�r����f��N�-�PNev�nɗ�>������_=�`�f���I����e/�������� �o�s�3�LH0 �(��ҊE� ǐ�&�(*�5g��]f���轼�����~̠�2�ϊ�7oܒ�[7��M4�����nI;=�W�Y2�pz�o�䟟�1���?|���'��I���Rr@.�J�iW�o��3��o���w�*?3�%����rxx��W뀢\\������ë�L{�a�Ч��߱v�[)�S�	UF "�;�Щ��í�����16n�ٱ~�`���=�g��������~�A�d$,YHy?$U�40�EĲ�V��`���f%%�F�H���3�'S�L�����q>���# z��MhH�GcdV֢F�-;T������P0�A������L,��B�=Z77w�� ɢ���`��m��a���?�PX���ߤ_�� � ���F��"�Fc6L ��T�X�:�������Z�S��0s�I4E"{ ������vڞ��U�es���^�~X��櫕7����${������)��x��t�,4�A�^��ۦ�s7$���bAW�9;tc`A��q�_���x���XXCF��g�jE��W�S�"x&�O����jiU(���O�����'�l�zG�����{U�2�>�q~�� )��~�j�����	�6���U�߾:f���`���+�(��R��A����AB�!�w �j;�MO���Sf��^�DE3���>�rx~ [;�Lꂞ�}-�&4��D�gt� ���8-D� I�Dί�mJy���|�U���Pr�6���ǯ��}��\855r��3��G�5��Yīj=yCg]Ӓ}�B���1]��'��K+��(���|1�r!)���$��kؓ�J�,�A�ΰ���C���LF����J)��7������� ���Dc�FyQ���l��oKz����V
w���z?�����X����Q����� A�?K�C~�	3��6ӇC� � ��Cko
v���jwI^I�,�96�/��k�*?��'��jR9�^�^t4��v���"oH��ʽ�z��с�_^o@�'��Ɠ��X��� N�q� ���A|���^�FtU;
�m�%.sb(����>����������4��r~.�� "�QPbzߐ,�(��2EF-�9�1�q�󝞝�Q]Z��dQS8����Vw���	���(?�����9ڜ�s譹��s(�a��ơ�H:b�޳��"��~8h�n�P���*�x�u�Hͺ�:�w���w�}+��7�\]�Q�F�Ҹ����ev�Ƿ��y%=���3a�tr��Q�eW�`D�"�ޯ
�5��-� �|��3��?�Z~��o��g������G����������?���������Gy�g] �:2&�4�������=��]����}rE@y������༐?��O�t�{�A�O.i�N����2�ܒ����� }��q{K���
�s��l���J�/��5�d r�Z�	Ơ��9s��������{���_�<=^c:����	�Uwz� ���{��-�f��&IU-��� �؁ �&x ��Yl��
� [Ԙm�����.�����3@�� ve�d���c��m�͚���,�%�OC���	�Xy4�^\���:�g�/�зՎ�����k-� kGn�m�>swg*wH/�2'�4���g��Eg4���l��쉷i�i�#u�g��o+
t���:����
@�c�܄�
}�.��:>9��sN�L��בuͤ�T	T�����:��>����a�n������ݯ�F�@�R���UB��)[�g�\�|=Q����Wn_lߏ��j�
~i���֖�b꩔�x�ӳ>�z�!���@����BA��;�E�_�p����x?(;�\��w�>���S�=��rO���"���=mdJ��t1��6��U�ۯ5��M�h,���O6�늽C�x�6od�6M���K{��9hK*����:-���O+2�ln��f��x�@Z���<IRd�QVU�A��hא��
��G�L����U�t�L��������@A��qs����ZN&��D=7�
����*�sNJ84h���EF��<jǷ���H<
n�H�XH3�W�uͱ3��$>�l���'���sӊ]r:T�t]w {{�AU�j�D��~p,kչ�҄���"(�f�z�	,�W^S�)�`�5*�h�Vtj{C�d1�A��6�-�k�����,���wVݩ��nY�CК+�G��pI��M�P��hf)97�IRJfP!u|���Y� ��(���aCɫ���A�bI�B�i�S8k�VQ�y`��H�:}���R��}]�off������o��qM'���񨘏u�]i}�i@y�c���^��0�wȀ��sp�wf�ϻ���5Xޜ��o��ں0��@������%I�
��|B)5{xz�u-�B�S�nb�`�V:Ȳ�SX�$�lEg�,����s��f�t�-
b�G��z�~I�Dw����XS�)����x�g	���\TjG��t���gk���M~^�_גjqG��ی��&�J�ц���<?�p���SF�ji���5�=鐈���C���?�x)���GE�V#�����E>�9����٦��_f:�HbD�d"���mFy 0�����zV���³��d���1<d	�?�~N�؞�˗/ٯN�_�]�ٜ ���B� %����{oo[�����~#�������}��N:���\]t�������o�&��=�ͫפ���'�0Jo��l>+myv��x�B��yD�Bd��ϕN�15��׿|�L��z�VJ�^%�ɓӣ����6e�������;�(}��tkd%�y�w����b�/�[��&��D3��F�!��O�(zc,���޽{O���{�!��9<?���9�:�����N3x<�c�rWZ�
\4��{`&ZR	&�Z��Џ��c���&S��zG�/j�nޔ�y\�I���,�{`LlL[ʼ�Ή�:�7���sآ���fO:y��l's���#��`��n����Bwdk��;[r��}y���L ؉�Ŋ�Akx�4 ��0jI��ޡ&��վ� }7�^�T8l$���������S�������Y>�+����	�ǳ����0�f�uv��w�Ko>��ι�w�X7;����+Ɗ�j��gY֔<��켚캇�Օ�&�]�f�����"Q���#��4j�0g�ۖ��|�e�Υx�q��z�T���LiP�e(�b��6�;�&��`�����ߠ�]��7��(N������J�}�{b(cP��v����޳]����~�{g�R�H0��|6����ݔM��`'X3p�=�|���AC�	��EP\/G)��,��[K��`e)�`���8p��9����X
�x�p'��Մ��I�`ۛ���:h��<�� E/ΐ}�
$��h���S*�!����R��^6H����^����)`�͖��?��.`�/�\���ȫ����J׮��βW2�d;� ,��� ���P���W~)�̀kVïΩf���ڕ_w��	w�ڍD{�>0�ל�'C�L�S�*��j�������,��JC�e�HD\%��~�n\��N�V�*r����,�1��.���Բʛ�ղ�Ӌ��R6��0�DdP�(��YKF(�RW����Y%�\aA�BRg�U�T��4��_��_��=��_מ�������0���j?�A�����U��FҪ@���ʱ8�s����n__$b]����x�OA~�΋���6���ߪE-���B���g{âƻQ�J:覟�q^fu-���`�K�G��ˮ�t}��}fwу��ɑ @D6)�>�k���S;�Y�37tZ��|J�V8�[����`#�-���On�#������5z\!�/�Di[�<��uqq���NUb��lRj�q�A%���
t��k��S��6��ϑ,MP 	dެ�-�P�h�)
)\�v r��C��P��ۃ�#��f�3�_����/�YU�)��Q���)�wo�j��T!:W<c?� \*�r�x���>h���Md��fbo�������w`�J<���9��}��������� ���������ٱ}����цt�ޖ'���6XqF������Si�~�=E�h����#y�����C��],��� &�zPl�4{ur��](�n��Ǉ� .�BDk�S��Sy�b#��]��q��AF��Ҭ�ݻ��嗟e[|����Y��>�\���Wrx��Y^���������O��\��3cV����'*�5��[��q��7���kXr/A$�Ld��l1��<w��q�o��������"FP ͠��ݼ�zb��@�ʂ�{K�38q����b�:�+���bEZsG�i�Op*�5�A?�<~7v�2��'��k	7is��C�u��(yT נ5f[]����ZCƮ88���u�5�>��tP޼���E3˼�,3ŃP�G�sg=>c�'����n�����[[	���L(��^�2����os��Z�d���.>�������̫%1�uS��IUᴳ�����p_�pݎ���p�s��������ʱ֨��[�+N�L<�|.���d|J�T���r�漐��mn�<��Dcq�$~����pz���րT}i��=�Wk�S�]�O*�Y ��~c��4h&��-�a����0w��1�Hz�����N-v��W�Ƃ<�E����f9�(�Տ�������_�4{}~&�B��Qp�ф"��ڀ���F��e���涱�˱vfG����Q�_A���3y����F�A7���M98̆JƦ~r�b����/�~8I<�m������FdெP帍n�A��pz�#���ԫ�m5�%���]��A$��k��`<��Y2�>���I��P�H��Ah1���|�v87R)�^���F�s���ǲ��څ�����C2Z#�D6�l�7��BrU�o�),��R�[�*>"�JI�(�ދJ�Z�b�Tj�t��<H6��s=���|���3�򳏭Ƴ7�0[��y<�ދg�}TW:c,�D���@��/2�,�@�`v�L�$�_!��c�v<)�>{`-kX_��k���:7�AK�y�P����٘p!*��̻>��V�V����g!�2��΋�3��-���3k���?x�I<t�@��j������ pƴ�&��f�us?���<���x��Q?˲e.��E�@�78�0�����������6���BF�mlӳ,9��T)��Eo��M���>i/&�A��_S^�f�p��y�!�od�y�@	��ʮ9��1 V>�֤������X�Z�1�8��;����F�5k~Ȝ�ϼG��ڳQ:|�x���8��C����A��կ����=&���*� ϫ�Mu|�J���o�o$�y��`�3���[��;hCL=������(��ȇwǬ�A]�7�>|��0 �:'d.�6jG[�a 
R�hҚ}fT0aL��ޒ����W���|�p��{��*r��<ᠫ�);�Qnܐ/�|�����e�-<�_�2�ܡ� 3)��>F�b>y�(��O������˗?1�Ց*�򙣗ם;����G�s�>aN�N�����>��)�2����2��x��&���O� lǨ���9��kC @뿣�;��ew��|eP�R@�jGX3S���B���wDA�a�� ԏG�O������ɶm��9���ؐ�� [��ӏ���W�".e?5�zg�t���6͊��tX�e�Ʌ�$�ڹ�.��h�D��0� %?��� IG���ꀬ���<�!�tv*����5k9����F��V��&�mkO�X��IWUM��Ve�V=IJ2���ZP���]Ջ�VU�F˔_W�CF�|_���z��L��|�i�����{��5eQ$�XT���\������g���o���_[��;���?�8�7�ɕ��:K��g �3^��_�y�*R9C�����L�k��0��|�ξ*e�SqFH)�1A4�g>u�I��~Ncj��7�E���hݺ��XKٽ�2X�"��/o�΃��ĩA���N��d ˢe�l���W*�+�\Qf�0'�\����6t|F��+
_�x�R�/�����dmo�f#�}Yv�&�Y�z%���T���9��Mu��� ��rox�E0��0�o��;�o�M/����V ��8��AF��+x���0�}k]��7:�k�Ɠ�}v�`�ѾNW�8R���cW��4�M�,(wv<��c.����F����.U��E�-�:��^r��3A�
p��`9�L��dY,=o_��w� 7f��4T��>�C���H����io�-�%~�O�0���9�.p�jFNA���k0���(}N�����H�*�)Tc=������?Կ_�szm�Z�3��Ɂ��\,�A2�@��!��,:���)�O�o�T.��-^����)Ew�`'�s� ��x��ѼA1�A�F���̲u����z�
T6���(�&!�����ӳc�\�"X�Q�'3�R(��&d:p-�`}G��w�P�� g��S:]t�)0SIs�qmYH��u��b�s����)ݎc��V��{u�*�!%��|�[[�t	�Z!�#��H�Z�v�pW�*ม�X��N��^6���y7c�7�~�
��<f��ƪ���?�(.�]��������l�h�n��jW��7�]W�������}���xL��1�Oy����QM��-��׿|/?>Eq����AM;`,Aq7N4�F��5�7�����[r�����=�bg�H\APj���N�圠k���Mپ���}{,���ݭ�G"�(�h�߸5�#��Ŧ���ѯ;����s�'G'&ݾ���6�փڐ�ĚP�{�!������H>e�u.s��jTH�;D���%h<Gdif�W�됭�)떑%��Z�:�@q7�c�ַh��L2 ږ�h�"*��*Aj��@~��@a�X�i`�z �	Z��D�Q��-��?��,������ ͢��p����d���k�f�-������֢(`/dG�p��咪���UK�~\��w�µ�ǥ���j�����ȥΑ�g|p��U����Mj ��R�Q�>����GF��,��o�d�uʤR��5Xtd d��k-ڸ�Wp�V�c����i�ޙ�LpchOt;L���z�IHp���	�o��O%�C�~�]����~���%)ͭ�n�@���o�~�D�(x���b���� �5�Gח>����%����
jpc���P�|N�g�D*5Tb���% V	��M���oS]������V�	+~�Ʊ6Y������YfC�9�7C�U�lES�ғ+�^�� W����ٙ|:ji������Ǣj=z������a+�:>�
p��O4��ju$�(��$^K4,�)����#��.��V�[�|S�m�����/II{�z�6��s��g�V���)/;��z�^��>,�5e��Ҥ�Hna�����n_xV�Hl��Lr�E�޴X���׺~�H�@1j��t"V���oG�����΢�	��hV˜�:��gG͸���{�������Е�������w3���Gm�S8x��)(�9�w�v6W}n��#?�NF���f����C��o���N3��P����J��l�E��79k\��?v���#��U��9p`Ll�C�d�sI��u�G{<uTi[���&�hH+��I�Yj�Ud~��f�@����,Rl����k�0>i��R�(ܲ���M�ǛL6dv1�H�G�|�����Q_��\á�H2Y�����J���c�.3&� G-֧O�
�u���:��`�X  5��4uް��Hq��ʘ4�ųg�wP���<f���gg�:�5�fC���]�A�Mg�f�^���N-����}t�6i���{ਝR�QJq��8Á�D�t8�/'c���Z���ͻ��*����s
/	VѼ��.%���3!�1�`d��5Jb�+ؼA[�5c��೾!� &}���:���^dZ��ۓg�z"_}�+�{�����A[	i?����i�U=�s�[�7�JR������.� >�u��J7z!^SdM'����9m�ك�ٺW��Q� ֠{X�"u�\�Ub] ����12غ�e`�&֋j����&�UD��X�(� �,�olI+�a`+�m�:6 5�;�P>����F�.��xfbD@+|V�z1)gF�*�Ɔ�ޛ7����{��B�#N���Z���*�b 
-˼��0HYl��[k�ZNF���c�
�4C�e��L���q~�`���^1x������F^���p��,�ӥ�ה�FC��@�I}�������k�epK+*�����~&�E_��b�N*"��� [�$�u�[- W��ưB`���={�O�2��^9��[�&��t�+�"�o��{1��@��K�����9oBWKL��鍢f����&�=���v\s���\
Ļ�ߛ9vP��!�]c@*X�'�R*"d �>n	���cr@˰�hR��3����()^��91؊�W(���0YJ�#:��e����E��a��6�&
ؒ��ܿ/��==��!tQ,m�̧��Z���<����7j��	���H{�`c[q�@��]УӠ�xj[��l�=sv,���x�M�Јt��L�i���P��&7[���$���]S?����S��u>= wL h ��r��>����jE'�c�5F��J��8�^��-�m$����:�,��ل]�
~BwQh�*ZR��S)Ύe���q�Qs6}��\]���f@[t�$y3I���[��=v�4V}�x�
�,6Q2*_R�Ůb�L���$ϐe���u�D�Y-	�;��N}�c��0PVC� ��j@����2$���c�u0k�Cj,
�_Y��O)YԵ�DZA�l:QJІ�ui�{��=�Xё�0�S~N5����A���9����*곪��b�m:迕�e������a���Y�wֳW:U�"(��N��3ZЌ��'~�X�!�`�6U�0�X;�ؤ�W��F;w��b�t2�1��&҂&cu<ZspA������qvL.�b��\ �e�0�3�1ƭQu�V���N�_�E�)8ډ��x��";|�N���ֶ�0e'����W�<r����<�su��[]���O��4�}lJ�7�􂪱�ç�
�����;��������l�;��l�n�De��0:���+"�cU��;�a�x�@qbm��U]�r��O��1��W����ȸ�>�*��O'�rt
y�|�<��ɦ:͘)�9a���Alj�R�)�46�ƺ�lƍGRm�R�qڟJ�e2�š�Sg΅�\p���lj�y^A�t.g�P�[2[1"s},o߽��?�Q���ȋ�e�T�y7��e�c|�H�j�Vj1wOZi��:mx\�Ɩ���_���&z��6�:3dR@��S=n4h�
ٙ������O��|��ײ��-[S�sT�Z*��$?��:�y�6v�����k��֤ab�j�5V쭦�琈f����\v"	�^��v��`L~��U��ʓ����Y�	c8� �g'r�8�U��>fI5�`:���f>�v�)�z��g��찮La2��6�U�)_�N��Uܔ㋕|�\���!�Ӎd.S�GxM2�����^���^c*{�l+�ў}���Po�ގ���Y�E�,ӭ�rc�nYw28�);y}x�Q�9�Lr��"��-����h֨3t�h#q�R�L �d�O�1���eG�ӌ�v�q�"�
u��<O���X����[����޼�$��ɇOy�����8iI���
�`?���֣:�O��G�� 	Yױջ,;����F�l�@�`� ,����C�c��ڂ.���N���1����<��\Sg2d�T׼xus��s�U�ϾQ\;_��g4���2�b��^R��8z�� �ac��.����, �-RV��NW�]�Ml�����3IqLz�&��
8)l�4�՛�H	7dj{���K6)������w)M��Y���P�GU�0��0ꊗJ�\�Շ,�
�ҽ��4�z�b-�0�Ea�=�u&���W�󒑸:�֑����!�E�����@G+��
:pR��"6*���0T��5�@�0�bA7DK�{e�X���EA��R��M�����'�EA	IZ4�PUU���S�O�/	Q���^�;�Z�|�Z��>8w΃y ����QY��Q��u_�Ή��$�wYu��Y33�ڣ��]/b��4�Ty���� b͆8��r�,�U`*V}�D5������t�E><J��B54gðK�q*���\���W��h�0X��)EWnp��G*�C���1MuD�A
�[�b��<|��;J1>����{�אb��R6>�2`f��_�}+R� �و��1j�}�Ѫ�|*1�`�r��N��P��:>U���N����N�v��cfhd���d���ى������w���+f�A ��Ӿ�+x&W�6kv�`�Խ.//X�tttDYe|���!�g�����p�t���[�BA�@�{�x]�>z�X�3�Z��'��A�bo��Yv��׋J��!�^����	�"�(f�@^��!�pm�8�P�p�P�;=�G�[�]:>�uh#����Q@��=H�B��9}T�4ꪵ[@���5ٸ͵�B4��t{y�o��e�q=c*�Ig����������Ў�H�E#��oH��5��3w����w��%Q�Hx���;Lf�1��� �T���f����������~��޽{O���B�Ы�9b��ꡪnM�{�����Ճy�\I��L�o�FUI1y/�ླྀ��A �x��)m0p0x��1D'j�������_�ϟ?���b�=![P~1��L�7�}�{��jJ�`��5$�KM1�����;����X�$Tp}}�^�x��A��y^G�&�D/�?��8�]a�� ��㡞K�0U(1�TY;'�"� Y�	�b0����]Y���m���)��Fja��^�O���g�����^�Q�� ���d3s �Ƹ��K?�����!�P�O�кDc*���^�)�Ǻ��Z��f+5���q�h�~�R4�2k�yc5 ��p8�5r��o��wx���Ƞ�b �2�Z=D��@F+9�X�!��wmmE<���G�R���[<�0����g���3k9`�c�|�y�|0�`z�z%�D�� ��IC� � BU����Γ�S��N�ѧͭ+�UGI*@L/��;V�z]�F�8Z��__?��@1)�Q��\��ͪ�g�EnE�8Q܁�zYgJ}��=(�7\��1IaJU�4�����G���f�.s���	.�C�%��EݻMl������0����j��
�=X�h77�{�����%6.�:x.@R̾FW�N�2a0ư�׿Q��)v4IޢVj�����ܸƧ��V��Z�V	+��깄��* G�:�-���٩m]��{��>M���l�T� �S�gܖ�	3�U&P!�Z�E� ���K�iv�i���<��k����R�޴���o*ס�{]������2��V@�1��T��:}>,.;:���q[,fW��k6�ny�:���p�#�!�_�S���J���֊�ߵm��yRӿn�uЗ�NV;\�m��i{����k�ƙ
�U�E�$�F���L8���S��d?Ɖ��}���I���O��Y���:?lRۨ��,1�!��&�kH�ZB���Y�`�7�۫W����%	�J�I�.X����¡�.��Wc	���N�����+��$<����I��P�PPy@C�67hqa�&�s�}�&C>C9;c���T�g���uGR�P��4�R�V�-��q�$���XMg�^	�mzbE��VY'g6	o1��u*rl]�N��̆���INT�i
�W��bkgqx���VJ`�2Z�oa�Q2��b0+�s�K�����R�۽�#����h{{�A�(�5�IAޓ�l	Яܰ�Z�`q�V�N���C��\�i��ت�pdx3�_��ts}��#z��	��ܠ�̼�P̓�bk{�~��?�?�`����]��f�����ڍ�A��\� $��+kkg�� ���4T��������;����)M��^=����$T��/�ҧO#)? ����.2 _Za������ɑx�&#!D�r�ҙꊶ"A��e�sŠ�@�
����y �@�g#�tzr��%��r��5�U�l����g�z�4�
� �A^���"rv���1����wp���� �Y�cO�?^j�2����p��!x���%��B��=�OCIf�i�RZ�ݱG&�}qvI�<g0���5����|�>|@s�t�2j�����zfP�l�Q���S�2�³է�%����ޙ�`��� ِ�}�|�w�F$E�'���֣%\�8p�2ȢHF7�óK���,� ����I��R�J�^��)��:V�_� J��=�O�0�l����`ei0�mJ|>���(���:p�X��@T�����S^[��䷙��L⹯�^��OT��b"tI��)j��пPx�|M�K�t�b�S~�9"Do��&��/����B�#wvؼT~�xLd��E��8�۽`.2O�Ҷu��u�U[||}p�8��m�+M�>'����Z��%���:P�)�,�R����GA,:��r�RwC��ɴ� (����Q��H �Z5��@�آP��wм��I�\�\b���W�_\������{%�{��+>�W�M�!B��`)Ư�YC�_AjF�yԻ��o褈e��}�>2vA�l��������ti1H#�HlC)f���ҘS�Y��.�o��k�hk��G�S��Su�J�[	d}���8���JpH�ɉR_��l�^$��,T"s^�M���\�M�[�;Ԃ3��3P�kkA1�z�����,�i��3�DS&bm
���ZR���Ja��x�hLMӵ+@����k�����}a�zWm��!au����(�T�CĬ�\5�o����}���E� PZ�Z�6[����UJQ�=Yh��iB�"���� `�(x
��|E(7bG�Xc���l����#d�*��UE78E��4�4�:1�3%%ؐ�	ؓ�v��4V����R�DA�P>5�G����dx��+�y�xʒ)�`�re̕d��(��ʺ�Q�D����eZZZ�'@5�xz��ɻ���6mm}a����#�T���U� x�$!)"�p`�
�X�\���Z�Tv�D��͵ZN�k���{�����"=|t����ݿOs�<�W�:��y�������_��w���-uܰ��N�Ί0<	f��לIn�Q�x*NN䃬jkk��יx�����ۼIc�,�\��YQ���ٹyڼ�R7����x}� ���X<Y�zG��[W^˳&
C��AM��.bԉk�bJ�y���J�&5� ���XJ����D����9�}�����H<Z�~� pO�L�#�c�4���	�B��=~jF��7����!�0�Z����,-,��<��e�0������0��:Q�ԭ�|�b�S��M���`$k�� ��k�%ʩx������c^������I�`o��i�^`��5�aT�hz6�vF#����¬�N޾u�n�ِ�@�����!�o�lB�"�UB㯐�6�3�0�`y޼��zi����Y�P�l��\��(R�� Zų"�)�K���#2dD�
c���T�"j��s`�o4}�s��*+ʴ��v�Q^�뇏L�Y_��Z?b,�Ē�W}BdfM���� $�gC�>���O���.�Ja��+R
�vctҩCq-���[��PgoS֋�c�3�QÂ13	G�*��$]N��0$�� \��[���<Y����d�|�t��p���
B\u�i݊����PP%a��NV�Z�jټ��*����sO,8�k�θ:�S��O7��,۬��U����0(�R:��z�+j��➫0�K� Y�Zw���+i�h��ʰ�[�$�����i���r~7o�ԦtX�|��{>�p��4i���`�C��k��QhBtpD�'>��`V�F: ��@JJ�)I�tg��:u��#	��`���w������Y�XK2�Әc�	�߾ %�N��޵k�w�k=)�*F�챾��X����t/kʹ��S�0,��� -˼R����BF�����W�2�֓Z͸��^�1t�6�p���w|�P��B��J
�{2�܀|?Vfu����K�bLɫ�(� (�����0@���ͻ*9S	�������Fk�=����봱�!,f(�~q~&
���x��z֓V�#y=clhYص(�M�B��L�1��1�yP�{$ ^����x� �� �P�Đ+��f��������r*�\;���9µ/��x�1ә�`₩�V����>�I*��=%�|*�U�	Ӊ�NFa-�P�`s�2���*SD��zMP�tR� ��XO�B�) ���6���]�FG(� �[��Z�ho_	�_՚; '�����W}3)�E��o���B����LYVZ����|yc�67��ɓ����}���I7nܐ�N�W�Y�W�Wdv���O��0�8:<+�xF� �M��
R��<f�r�wA{�҇"�XQ�����3)p,�3�����s~8��<<���97��':nq��d`|�A� X�f�uյ�Dе!�=m_��i�X��F����r0!C����	�<h�!g0?���O���/���6��S��揲�up x�r�y�_�s;��` ��D[/Z~@C?��?�Έ�7��V�fiuy�V&�<�7��=0���l��0xL�U�]?�:r Q爂�˫t/��;0���|�@KM�/۟ū7b0���L�ˋt���`_d�BeW�`l{z�8[�Y�K+t��=z��>ݺuC���p_B�GR<��|.���٠��Hv���!�U��l�D;\+3<��WE�},����V��svir�]�?|�u��m��W�?��������8�<�~�*��v���O��S��_v�����X�Ik�GQ�9�R��:c��	+J��+��8|,�w(��N��5]������眃�F:*>��(a�Q�LdmUY��f��y��R��*0�-@r��g��:{�\׳ڳ���ʣ?<<P�:�����v����J�`ls}�R7V�Ea	��Bӓʕ�>�:.m���|:;����r�kH Y������C�bHl9"J���k�H$t6c:�-�M��s��U��s}�܌�t���[(��M� ?"u����	+�u.�����B&CZdY��b^�cF킫x3��aŊ�-i�%�G,@��E��6EH�>~yÐ�τUj���@#f&r`ꗍ9_+oP�N�%���o'A�/ �}#�E��hT��
(���i���ן��E�-�3$�&�C
�6V�Պ�,������è,oIR�@���$1�S�z���ȐI����f)!��0W�ڴ��~�뎒���I�Q���z�����	�)rK@���'��[�����Z���V�Ч�V�$�}Y2�㇨$n��Hd���d6&�?kt��fYQ;�x����{WF� e�0 42�gH'�lj�K���q�0��KEf��n	�_8�d��V�k�u�cr Ԯb�w8�a�$Ӧ��� TxI�	 o��c~�ٳrp��������(kǪ�5�	����!�U�&�d�'�'� ����'d]e98^�dm�����k�,xvr!
4r�@'~zv!�A!�����G�,Z�Z�.���KC/��*�bg	�S��P ؗ5�"�<��w�.��/���P�#������1���9��O[���kz��Kz�a��PȘ���ãs��1}�ڥ_{O�Y �YR��AX߾yG?|�����x�P`� �Q��2���ݓ�����K�{�m��SaFm���:�c�}�a ��xp�E�ų���"-.-p�����le�!%@ ��y��x���<w7�ރ{t��m�Ɯ�+ɹ<��_vh���c��*�z_o`��6heq������]:�wZ�A�ph9J�!c�_P�
����	5����r��:?7ī%��ܒO��mq�Hu]�C��o�/`5!x�
�5��&c!�3�&� C�RBኁ�;_��ѥ�g�cõz)d��i�2���,�k���Ѓ��ie�S��X���MC���D�Y!+$���v[��[<&+n�9�Q+�>���-/Q�+Oi�� ��JBYҗ�]I����Vr�n�ZtSh��u���mM�q4�Q;1�&�ycJ���6�1ۀ(��#�W�����l�I5��s�rIo���`�RA�B�p�B#$H��r/iȯ'r/��ε�</�dd����񔜨Ƣ�Ҝ�:1�c���o�gko҃C�Et�)�����J�׊��S��1Z凬qrH�ʮ׺���W�s/Y##�f��Z�Δ[l`Ӓ�lC��J�uU51o��cYuUi`S���2��dr(������{�b�	n5��t�nʠ$��ֆ����+�y��
	�8I.M_�v�]䱸�]/��j�ʶ�t�������Em?sX���o���&�+F�,�.�q4�cP����%*�����,.c��n��m����L�)�2�bl�Q��e|�}%_"�>v�X]{��;��!��T ���V��.��&�������p��Fi?���)����i"_y��{���<G�d��c
�Z*d7AXC��5���~4^K��Z�H�����z�z��%Uܳ��nߦM�?P�?��dx���؂b EH([U|��h0�b�~7�yD��B��=ɽ ��,_seYko�P��d�Z���6:S�Y�D�"�D�B����3 bQ��,�Fb �=亀�\�jMFl�(�wߏJ��!|��ˠ�� ��}u��H \�b4��'�
I���4
��',�P<}�z�׼k�K:����
�K���>����A�u���֌zH��M���T�V&��~yG��s)xN��A�!DN��(&,/FñP|W�!]k��&ҐA�ʝ+
�b�2�,���1�Q��HH+�_��uemE�ó���g�x=(�$W�DG߂���/�˯?Kn���a.�b�IES��ޥ�_�����Yl L���	Ŗ�0��S��P/��7�k@��� �L @&r�旤�����Ȟ�5���h��cR�\0�s����j�/4~�(C���� kDc~�g� �{x�6�ޢ���&��7��M�/J��g����yF8ܓ������&����m��柳����s������%O��g^����ݻw����vC
�{!	YS�Cm5�t�x��r��S��F�o�^���2����P�o&�X]������ ���P�Ë��"l ��C=fv[���<J��(��9��3C�f(�Sa�k�D��t��f�:�}���L��u?Dv���Op}�L� ����'����w]���M�x-^{1�-׭JV_��uAoE�\F��̖gE �����"+�T��t���z�yL�_��
��古�_�-�Ϫ�;�F%�z�cwJ���r}��c`ˣ�,������>'f�2�㡅��[���x�<W�ۚQ�SM��r=K���d �|r�Z���U.P09VQ��3���R $�(��
B(�L�)��'^@Lc�f!1� k!-��P�A�\+JJh��|����19C`���-����N�b�'�3��-W�]�1�~W�ɬ�Y��+�ff�`R3ML9�1m0{��v+CZ�iZ�Qw�%�i�RQ*��l���ڕ��T�ƅ~Hc\���M�v��_z����8c�?ߧuKFa�s�$߮l�;x��Zt�oI6z�t�Zu���7��2�����}�+���Xx�-RL�N`LΔ:Y�Ca�)]����&!G
QmgI�j%��0)�'�S!ԣ��o�I������E+S���:�W}-\�CVaȀ��,7)$P��*���=5���H^|0�[9�l�x�͑q���N�0$�i��I�V�5՗0CX_'R�B<1 ���Os<���(���湨�C���[�E1��Aqqq&�S��o���X�D���{u��MڸuK h�%7����s�r��8�׎�@ѝ	ZWkF��P��G#��(�G����X@Tk,�Q���X���X�`S��J��75�@å���
@_h�t�}�"D*螖#VP��Z�2V���Me�5�c�so)�)o
����7�J��n$�Pjy]�
�,�?3��[�ſ?��!�p��g���6Ä˧hL�5yq�N^��Q3F��M�6�F��S��0���7�
���=~�>}Bw�n2���:�,�!�i�޾�@/_�L/���-����:V@ ��F����z��� �3��o�~���=��>����R(��{��>��ѓS��ՕV��4�6j-Ó�c^���kV��o�)$��]�`�.,.���"��<����hH�18V&D��łY���Դ��@kyu�A�����v�@#�4hz\��� B��k���=���c�{{�V�fy�����6}�ޢ�鈆լ��D��"æ&;gy�n�/�\=�wn��'O���ZY]U��kߓ�=��@7Yh|��۞N!�M[����JX��s��x��h��J����:�8����T�� X �"l�2�0ɒ��ȏD=K�@O4lZ��0:����ʦ)��g-BQ��h��)۠l�=5�G-��J޶ɝ6{*�K�!ev��B���t w��Ώ��ĮW^�Y��-�E���'�s4'��*V�u<r�vij��)�� �0�ۧ�dp��o{��s���3EI]�p͘i���W(�E�L0c\���;>�A���!�n�R��`��������Y�nh_z!�G=����tڔtք����z���v�W��r�MgB��a{�p���<Wmn�Fdh<��N���<
��C����Z��2Q�}�`����à��zu���rn���Dz@)�R0eOw��Z�q�	k�K6�>��`W�<�����V��D��]�Ok���>���l�g:��_6��^�I��eDz��㺰���۽�Q:�qᒇ���*D`����,&�틉����i�����	�Wy��k7m���k��]�����a6�5�_���De����N�b'�{���ӂ�'������sa�Io�{�6c���u W�-��% �s�J`�!z�0%5I*���A��Y�>�˴M$��ļ��5��Cn��UV���S�E3�;D��$��R���wK��^�g	���Q0Ƞ�\%J>0�Q��S+�[����gl���~��u��])N
�����#�$�w�i�.�Mȵ�w�.ݻwO�lct��"$�#����kE�+�B�P6�]��nN����ũ����x�dG��!�0 ��F�Ov� ܨ�p�(9i})d|�
��X�nz�r��fG���6 ;0ƴhD"�~��1�7�5�7dz]�B�hgE��KI�譬H��^�~�(� ꙝ��������Z\���E��ب�t*�4�=��[�)kn��N�s���(�ijE.[}��)�h!�d�w6��/��O�?��%�nǁ����w��痯��}x��œ�����Ȓ�� !���sɻ���@r�1Cqe�"@�Tk{�e�F�ޗ�:�Ik���V��~Q���(�wzzB��r'9DM���M%�%g^��Z]]��e��B������I����\g%`i~���<r�Ԙ���?'��=�����������ڸu��M�ok<�}�,ޭe~o0Sk��,|x�}n�H9�gXwY_��g�����t�mlޥ��5��UoM4�Dy􇤼fP�s��,�C�\Eυqf4O	A�����D���,	y���w�j&"� ��� ?{SY�/�D8��T��v.x͜�sa�'�`�������Zu:���ju�c��i�Q���r@Io/�#�LI�>?�����Ͽ~$������JgjG ��y��L�vM���#�R�}�dvү�TJm�z�:~��Y&W�\C,k7\�$w��*�Yy����w�/8v�����������xק��X!����h�-e���`]0������[�V�a8���h��Y�_�(�e$ZA�_��n�^��!����V�*��Ҳ�σE1�q�,T�����%՚ɓ�j��'OJ|Q�G�ݐ��9ޔ���V�=1�S�n�%m���&�]KLnz�g#���~�<J�9|�|L�b�C�P66QI1�g�Ww7��]�Ғ�����<���s[�n^<���Ụou��y�}�M\zc���EKO!I ��.�� "��*� ��{�Μ\�-dE'�=�B�Q����PܴmId�p����	��b�a�� T���1�]
�ot8^��å\�}U&��O������{rt��[�H���Bk+�_1��[ĳ]nb_�F��{�y�*7�~�%I�BY�Y�F�p�������z��?�kȜ��DQ��DŘ~/&/�*@���&(!P*�vV ��Z[]��>99��D�+ZBA��1�nnn��G�����ρ�yX�Al�\���ma}CQQ(���N���2���E����,_?1���7�C5��F-T�����Zkd)ZO�(Z������Nd!hnՄ�>��P�kZ��J@g�2A���^�0&`�X�jZ�I��^8�SW�����h$\����s�LUL���B�.���͜�G���V�oJ�W��֞xp��J 	JT"_�U�׶n�,�Q�L!%�j�>�����	!�s<�7��X=�?��;z��sZ__�~vv%����mVo���^���vw����rxNzF�����`�}���Jj�M���r{��|a`pe���djޓJ1�����q�W��Y]�!��7�h�b��3\blY8>9b�-�� DA���=�8c�����7�:��q�H�q�ӺKS����'�f`!����QWq"����8���C�jP���3��L�����eZYEX�'�7J���wf�Kj<?���3�h&j�Q��۷�����{��kfnqE \d�^�98�MWM����ole��-ꑳ/xdQ:��0� 2�GO���*��m�1�,P=�нS)rݫ�t��pB桹�X��>��O��)�5�eLz=3��S�S�s�����'x]���|�x����(&/]���~��<������;�\a�.�Σ�-y�����f6&�ś]��I�2QE�_���J�k��%}�u�N�uGg�w�\�����Ǥ��t
����H�:Sy��������q�RW�E�ϕ@�z�b|�{nKN�q��`��פ�mw<�k�NNza�{v��k���<���>���n�N�>�ZI;����j��<C�`�d��ڗ�Z�TDr�$Y ��pPNm�abz�[b�x�l(�'�E���+q{�`��Dcؕ�#���<_c8��E�#Viz`�"Mx��*<o^�#^��|�^p�.Ql��1�Q�ɖ�Ґ6P�v2�hb�,���C��c8�02`��Ҋy1�G��u�x<�b�����Z$���֠d!M,���6�YJ����i蟬��AZdD,
�J1:�
h�^E׀��|;�#���Ū��RP0���& "{�i1c��u�S�f5V`])��3O�:j�Ap�m���ݕ�\���N�~�C̆3��*��t3�x�B�yT�R���,
-#����b�-D� @�2�����������I�xr�ʇ'dvL}�t��r��t���j�rb�~_�ǘ�R*��ub�C�I�%o�e��b�����k��W�І��hĲ�,�v�UJ>e�(�A^P:����	IQ���]5 s�a�ZVS�Ղ�}����9���ק۬�F��4/���ʲ*�sttt(�
�"�J��@F��~�����gz��+�G�C�dC��(�!X�@UI�ub� ��W����G���3�����-b5�^��ANɗ��Bn�ۛ�B��ZN�a��z��p.�{�$
*C9�B��(���cZ�2-��A�2xia�Pś�묀�(�������>���<������ǐ���_0(d0���G��9<���1���HΚ���ZE�©�V�~a�H�noH�=���-�桸1r��#.^8=��R���,�n�y�ڶ @���V����7�}��X��s��Oh{���8���K���j�B��5����|�jp%<�i�U�n����RR+Hqn4��"֫�����&=r�=Z�����+�{������˟�& ���T)�͌k�M�9j8�4j��t|)��uF��ynjH��sP�g������@��D�Hi�v��y;�}��U�yk��k���<5߷9�+�5!�l���	��⼑�B��6����t��!}��E����rJ�߅�99�@f�\���9���������<yD�K+Va�Sȭz��myHsKs�{�r���@�&1%ss}XC���Dk��n2*�17#�0�!�Y�������Ȁe˖���,�hum���*�����	j<ѵ<5f�����7����N��o�v��Wyn_)�A_�r��h�޽}C����ayqpr��j�֖nJ�Q�੥��V�>d��d�}����M����1��3��pd�Nin~ 9}j�����b��|���H��z�ɤ��(1��f��{�����>_ 07Lo��`�R��$}&l���+/�MD����W4Q�6�nA!W��8�?��xd�
��o�6�f�g{��Rh+�=Qv��cJ�lU�3�Nٽ�,�on-���֠�~E�Cȃ��H��Iu�)YX�x��o-�>c��w%���`��Fߵ�W���\猺�R��!Z�zݚ��"_zٌ~��MTW�Q��D���l=sE��i�Nߘѷko�*��k�T�zX{�Q	�QO�4���*��Rv�ZcF����P�k1�Z�j����,�<\�7b�������
&J�S�������'���P,�	L�~�
���".�v��L��:�4lE7~IMN�R�ʰ����a$�A��&�cZ��FU�=�n,���",���cR��Qp�m��'o���翩�>�+O���S<ܥ�-E�Y=��:�oZ�y澚��z�QH�<��|�u摼	�B�<D0	|���3�>�
��t��U��C--�%�K4�aג���V�C�6��r\0v�e�x��!l�Vw����ϒ/#���Ж�Mc�B!�z�<�)�]�Y��0|E'���!k��!�zJ�вd@ ����p(fB|����nӚ#ۏ�*hcZ�B�G�atސ��⍺s玄by���~{��Xy��CΗ�=0޿�^�xA/���6n�����<�K���G������������	�8�q��q#q�Ԡ/
��bܺt����hJ4d$	�ތ� ��!d���������������?�;�����}�}[i��E����i�5�(*3�s?�Gp��^7�Q��<�ux �Ϟ=�y�B����iow_<$ �5�G�M����pC��KI6�3Q�5�P������VV���e���@H���ݗP�_}E���y�d����Hs�:ڕU��ޓ����@�������Uz��>��O����s�o�7<?k���'���_���W���k�.GS�@I�"i^��SDP4���De����f��SO�l�V�`6�p�{�ٯ�o8������e�7��'r � T~Rޯ|�E���L�e��yg�@�W�D}!G 3ߝ�;<�x����=:�;a٠�R;@����y^s������������?��@�̆+�|y� G�@�0���3h��E���=щճ���J\csa=㉢��?��QK��X�W�<��T@/<Y�7p4�c��'���16����UZ3PC2g�^��:���Wx�/�~�����/���W���{�a���a�~��޽+���\���=/do�l���ʹΞ���D�J?�a*��o<��59��ɣ�Ǳ'
z0��>?��G��Z�����o?�|��
T�Wϒ��� ���ſBi�����
­�n��.hC
�����C�]E>�7�Y���rt�7B�ú�+9{˿��aV�zt@�zV	₫V��]ӫ�1�L ��>%�ϗy�(��v_�g!~�H�C��yMW�ڽ~�h@1�4V1U<ه��?����\����	N�N���R8��z���B���Qxj����!���5���ޗP�P�v�D��/�F7���PY(xh��B8��P��+��J�K���Jqgϕ��4�1i���!Zbc,�U�	���n~�@���q�� �����ZSe�Z�w"������-Z7ȕ��3G�/IZ�&� �.%pJ���i��K�������/�BS�N��B~���[�YM����_�e�hG��[���x��yni
d��'���(�=p5�����Q {B�3U��˶-|r6'�Zx��b��7�uM�X8Ut�l�A:��-�dg���F��� յ�}��^h$"�b�e�l�(LbZ<(1h�_р�C��l`�-.�� %�q�#�er��	��*z������ \�T7��X��P�����e�J2�,$�R�`"����h�� ��B8  ���ڍ5� ��%{��x�@����18�π�ɓ'��K"�@P���6�z���������J)�Z=�I
Sk�3B��@�!��Hd����A�~M�h�4^�ۛ�������?�p�`,����ϴ��B�$��q]_ߐ���L9J4�H�x,������fk$��c�vKx����{��ٳg������ν����K_Ծz��~��:�?��Dܠ(�Q��y��aZ����)��6?��ylVto�P�h�EMw����w���{�<7�D
A�0`�iba�B=,[��`������6
< ���������~��w�'��З��+�~��'�������+������n��h95�G+�	�*�7�\��O�m�ڲ� �����6.���.��Kc��+Z~����K�Ԧ�O�����%��5����B$352~��}b�z���JK˷$��:hϟ<~��
��}�@����]NDO@H���5^��O����'t�ƪ�a�<o��i{�����9� m_�&k~�ԥ���dP�߱H���f֌ 0)-#�e�0�����a����p �����3��tqcͼ̩�Z�D��J�P?0��P�d8 ��]IU�Y&k��Т��{���y{��>}�������D��H���G�����k����>|�=aӃ ��l�΢J2<:A�4\Z=��GVN�ݺ�ѳFΨ8�~��]����e���߲!�\�NJy:V:�)ǌ�6��`�T�+�%K9��1�BT��4ÚWu��eDOzI=���Q�h����;׮���3~��4��������~�b
݋ʁKw���/���׫
��AW��ӡ��L<i�=3`j;�%Y�q=�л|�=��x!�W�F#�+�-j��n�H=�t��b� �AAVsX6exhT��/�b]ʆE��z7�t�q��78�<�wna�f�$�V, +mBmb�Ѷ�F�麳oR�VJ�P��n����� ��k��n�C[�<,�*c9S�n���䥶�ī�P)�~w��"h���!��������k��<��R\ �M	�aj�OwA���1%/A���֋�����NX���=|�HH��R�Ĥ�֑�4��$ ����i91��Qeq�/Ni��H��K.H����ΓGc�ߺ�uA� Tt	aiR q���`)�%��r��u�˘�v��E��3j���5˳¼MJ}5<��ʬ�r��|$����2�J��d:�^�P�3�
�ȇe��{dMY�A��*4���~xX2`�1X@��:+@=1�\^����>+Q�$���
��E�t�8Pam766Ty���� �@Y�HNSCY	�m�����S^n�·�VkU���
��4�7��<��H���;9>��Q������ksk�P%��@�g����я?��>}�@�g'��)�a_Bռ�<^�5�E9�C�� Zb�u��uOj(Cl�z*�\��u��޹Cw���o�Pzs}��Yn�0�!�O���zxQ�9+�������;tqy.
����i:�dR�ȏ��{����V���Gmq��ȭ��ۧ�<������3�� �Lc��A��,?0�H�G���^��[�Aͭ��YB� <�k��F�y~O%������{��$Qҕ1()G4/9yT��K���p������{���������]^Al3X+۬8���5�����7�D�9�0_Q$Z[��*0 ����9?��F�`@���cz���#�s4 |��!zW�'�+j�f��Y6��b��w�B5�4��2Mr;f�]r8\��[����^Al�����DXW�x?���0��K"z�wu��&��gi8��y:�_ļ����=�K�������3���xm.)��gg#��r�c�Ko�~��|�Y R�!�U}� M9�̈އ��m%�	�q Z������S	�D@��1�3�����|R�JP�{>�ܠ��O.�=�J ��*��NS��`՟�\��.s����/b�9�ߓ{A�ݿw��?{NO�<���6���#e�wq����d�b���R�i�-1�~�Qk7d�XKn��L(a�8zvR9Og+%�u7ڒ)׮���m����MQϻ$�]���,��l���{�!���/���܏���;KO���U!���q1X�D}�w
��Q�+|����l�}^<w0�_,��[��C�R�G�6q���u����ǡ���V�vR���N��5�w��q_>��e%e#ՙ�l�sos[�ؿ�o�>D�A�ɍfIi��{]��13l��Z��hG�a�1	�#�E���;j-,�� p Ė��hi���yq���꾴��Lj�T�q��6���[w$q
X��|h��P��X�h�K�7��H��^ڏmZ.T�M�Ap�K�J����@P���3e]�;�yU��u_R!���7���Ȋĵ��"u�:{�������%���N������[f��ŵ�%���$���u	wlӦs�U�\^�g�DZE�\������J,U�� �4��B<}��P���JƏT?�Ș�`	`k�2c�Q�B��M�'�1/�{�wQrÐ?㌟r��<^�%�Ρo�,:x���N@��M-f_��ܤqѨ�b��:~�3�gE�+��K(@z9���v10dN�7�<)�;ɱ�@5�Ǡ���X���S�07��eV���'�����9�1��L\@�Aۛ&�,!Lº7�B��Y���P��4�4���6�$b����FRK�ѐ8�����0xZ�:xt@ ��ht%����F(���g�� �W��_��7�嗟�m�rOI6�����MV�.���H
����
�v0�mn)$��yK�g��Ʃ�T�� ��e����=�����qSI�@ų6��~��W`k�<�T�|�y
زP��B��7��V�k�۫W�tI��7�"���8,�M��&�<�3n2Hø }mf:�=!�P����+"��
�t�a�*R_���� ����J�g���w����*�ٌ,D]������+�<(�����Z陔��-%��F]��A�&(����O������?<���o3��ϳˆ���~�����sgg��}�	������R�� ����H��@Pį��{�����c09��6iyi�����>Ӈ����H�2f��aN�����{�?��"��+t�A!��PVƼ�z֊�!sR�As)x�Ծ|9�������3��u��=>��d�k`v�A���n�ܦ]��5��n;(��l���j�6B>�����𸽗�ĳ�K�8ǚѺj� ���� ���~�Z�iȥ� 7-�}�Rz�Z��<:���yJ�a�K%"���<~�x�r�܀$�vb�f�=�Ԉ0 ˰���E?:<��#
�d���2 o����ѣ��
��\��b}hʅ.P��ə��Y1��mg�{υ)Պ�#�r�����[ �敵mqp�aV��*���BL��"��=f
�$���V���BD��t�\�3����R0׍B�RWꯛk�w����g�Oe��ۉ�O�b���}�S���H(�)����GLzZ�Qa�@�Z�}�Yߕ���қ�(1�f"����G<�˟�:�}(�1��d�ۭ�!�:?�#F�����J?�0�½�H4\�W2�t�I:�şN�]�X84�ٕ�$p`͝�T�IҌ5a��&�)��T  `�5m��m>�b�(���b4!Đ�V�F��'
��%�]Đ��`h(1�tWj�:���ܨ��b��O��y4	��.ZT����
��1v@- ʂ��]l��Ut���uW�JH둨�h�̃���;k�W�&���VꃁI�L:���P"�Ћe�W�Gٞ�mK��Xl�h +;Q�����R��6;��T�y�p�bI�j�_K��,\���s�hW`�x +Xج�Qs�y��F�Mdy�.@<L*ʚ��֗��R��ei�)��v(�[���Y\fe{%I�ky�&Z�X��e��v�9Rae�V$��S�� ��[UQ���&�^�7���r8���X�d1�F��\�^%�h�,CF�0\ ��J蘗YiX��F7�V$���dQh�Q�
(���BYxqZl]��$V+ˇ�@+5�>}��B{{{R�
�
jJHw�o@5yM��lo��q��-�9!���v�����[;���� |�aN��H���kW�_��=m0�}�_ʐ�,���P��<���{V�n��[� $k�<h��R)����iK����9i����AaF��f�@]IX٫��q:�����, �>mmӻ�� �aXS\a�	�	Jt1������ B��mEڍ{ë��@tU�%/
k��x��sW�u�@ �H��R�g����%0w���ھ�@Gh���/������Zz���a���6nm���{Q����{���y�4S��4�N�EQE(}-��������Z^]E�t��{��Nք<jl���ӓsǼ&�L˺X��x!GPvG�F1����7��	�B�Nk����77à����
�����_!��B�P�����������CV�?�����G4T����t�J��g�th��R���7b%�:�C(���z���熐� ��X�gy���h��b�G6�B��h5��g`A�X!����#���/������9�7#j�|+��s�K.��m}��@�h��-ޛR(��)Lkw~@�#/ [D���I^)1����@L�l&�W�'>�,���=�I�p㆗("��ٍz�p=�	³�~�E�	a��}}��x��#
�����`d_j�W2=g&��zB�6�꥙���]�����H+�甤���K�Y���v�Z�>���d!J��'��Z���F���1f�!902-#�G� ���=)�N<�z�㋢M����.��o.x?�_2�&���S���hu�{�@>��))~�k��?\!�3I�3�E��^C\r4R9��ʧ��- �@��C�P���!���JA����g哊B��\�Yp8�-U#E.U���|�jL�Pғ<n=������1��	J�
)� C�B�00�'x�L���ޤ9ɮ=�琇��wyeU��/0�I�&JZ�}��=k��3��n[�0y �J��&BY�*'�� ��Ĳ���ү͢a.�`�W��wi��m�u�䐍�v+YuY��^ʿߊ��XsH��N(�w���G�l>s��ro�5��C�­�<���)��6V�4��|K�i�Ew#J�"MkCj��QW�Uބ����<����İ���dAP�L�����_��p��?�wؓ8�2�^x]�Ȉw�A���&`�y�E�8�J�r�F<=�4��%vJ�n�����iO�ѠT��T��\�@[��R8���&�G�u�a_ydx��h�vS���)9��`~��,�	��(�Pk�I��k=݄B!]�Dy���C"|v~��
+%[��~!lY��Cj�pD���&c�sG�)X��-��Y�9TU׭���˖ ]DV����"^q� ������3�����D�ֳ���ua݇��|#���~��޽}+T�Z��/��2	zyak�1���ӧ-	�ڐ�m��Lg�3���/��B��{J"޵9/�g8 1Ȳ/AFYVHONϤ]?�������>}xOǬ��4+vP�^�zM��	mږܲ�w����,^V�gn�P!�
ߠ!G��Ѕ��V�oJ��B���v��~�s���GY��s�A,�^��eo���Å��8�E���aac���4�z�F"�jq��H��Y\��0;���+���QB�*K>mS�W,j�M��Q�`�H~�����	����d�$c����q��rE�� Ъ(��9��r�p�d �sxC��³�s\�j�W����//��u@��C	����x�� kB^�hiX���V�d=yH��<�ᬆ��R��O[_�����R@j6� 4����%���@���-���1X��� 7n,�8,�����2�� ����y�_��D��?�����%��/��� )w�	����ؽ�ޟs4�����<���s4�w��h��-���D)/ ��eO^c 4���S0PJ�sA/�7)�k���?'@O4��06P�x�{j���0V� m�A 3�; �e#�������#� �G�Z�6gr��Ѻ3��x�V�W����d6�Wtuq%��R�OX�ղ(�\�&�%�0U?�=E\�5j;�\�qcbR�]�v!�'OL�(��gu�,��t
�\�.޳3��N�=	)}>7}te��o@���ۮ�;���}z�iJ�l,���U����h�c�B�*� ;�Q�!��7�J����;XV���C�%].�u�B��	�Gՙ~�Rp��� "�������t��S׻��+�j�.f��3/��X�e��z%L�l�4��(X�J�ߙ�Ô�h�Ee*Ҡ�(购|3DMx'��+�$U������5��V@-Uٺ�J��*�����{����?a�{b�c� 0�_�3 c��0#��RKb+,fʹ2*G�kۿ�L
�~C�;������\�����d�g�w��!W����j��!US-Ti �&0X������j�C��sE���hs�p�o��NO\�_]��X�'v���D
y�P	��$L�
�P%p�y��ڕ���`p��z
�P9@N�,J@K=Y!�+��cN��o�}m�;�G�8�ly[��ࢿ6CM ]��
|�&�_rLE���d��D,�:v"TR�}�VԆ���J��
FSY�2%KZi�����ߏ�����`��>����`�	�~9�j���J �ｙ>��a�b��R�D��H}+�	�D�j�������/�� Z7*{�%�/Le}BI��� ���H�i�XC1��)�1:�}&+H�i������q(�g(iPvԲݣ��%��<>�-?���x���%9T��+�� 4y�C����P��h{�3���,^��`S�+�`��Ç�C���r;ЮF�o�bYu;<[3�����zà��˗�3?�D�lB��32� @�����A����g��xƞ�O��d[)���pr(�A�*�<uW>��v�7o�(%�Y��ê�!�E*�	��t�Թ�7,�o��d`
>B����YY[b�F���Ʒ�sLg'Jiک���C`�v�j�%(�ȓ{��}���I��,��I����b�!�r Ww�ޣ^����Ԑ` ?�0f�� �P������^9E_�6e*C� >�e���2X�7����U	�G����BY/E��xX�Q�Bx���=x��?}Dw�n20���C������:v�o�L,�l�!��ى0r��p%�3����kan���=�4޻����.-�H��`!��~�~{�����+��_�w�>1 ld������dwO�(S
�^fI�ݓ;K��X�B����\��r�2�s��z��恀���>��tqBtq~*��3ɟ��<h���u�K5��S���{��&V���`�P_���A�	������z�縞h����,��m02��Ix`$��ԺU�8H��~n �xܐ�5�0^�\�z���BV"�mbaϾ%_�\�q��{&���@\��SQr6��܄[�k�sEِ�B��4�33$���s�T ��@�� [ű�����{�˶�w*������cy���l�4M�b�{�����v�sʾ�(�]����������I�.!��5o�#S���KI����DpQ�A�mC�fe���,�*�Iţ���&4��5�՚������D�EV���9�%�U��6��n@mku̻.ʤ'�������� �j���3>��T��F�EV��S�aWR�����{����,h�QOu '�(�.&c$���3��,P�|P%�d�F�֨�[V��^Kj\�	�^`�%e�=yš�UJF9�r$A��^��R����#$���� �������GǓ(�/r���' �
f�hc�:�J���(����{������U>L��*y9Kp�k*�`�b�y��M54ή�Ԍi�:ZZ�����!�^�Cr�2��>��N�W��3ot+�,����b��2���r��������)��H@�LL¾I��ͭ@�C|ASW��-ĕ"%���G��irɊPZ>K���+u �ܺ�F�����FU��2�ɱ+{LSW�(V����K���`o��7Z��2(}}P�Q�����X)��p%�N�6� h��#�/���%�Bc�K+�дBzpN_X��������O��dmw"�9�Z��}5"�.��\��(/h��V���}��Q(�_�~%��
n�߷6�jS�� ���ʊ������ep ��?�
�����	��d���� ���JC���U�F���������������!��8<&�痴��/���P�y�l%ލ~oUa7%L�9.��S�K���a"�`�����>��'�11�FA)�����׿��)��<����v{"��o���TB�P�ރ��2�~N�����Ǌ�:��]��3B1d��˺�~��+�K����=z��)}��0�!�G�va	[a_A�B&����Ν39O���j@�$�����f�1��/�w��o1�>��K�	��PW�x���hc���Ɗx��A;VV���i��'��+�ȭ�y`s<�}J��;w����Ҝ��Ѹ�5��.�?
I��הU�*b���0<��\�}fp5'��E�x�Qdx��'���YG�5x��wtp�}�D����׿�L��~�]���s�7#^��4��*��Q	 ����{f0g���� ��|� ( �s�<?��m^�~5���H~�C49��R+����ھ����x=���/H�� Έ�j��JH�����B���0ɡ�,��o�ߤ�;�����
�{[r�"��&�ΦwȦ�H�~�0���ʊ��6�%t�!��c%�q�T�j�G�NT�p�*9�JZmf����o?�Uv�=����ua@5����T|������A��*�����5ݨ %��g�}O���֙r�C�3v��-�G��nX�i���\o�x�Ώ�=C��5�d�/��	�0���fZjF��*ӿ�74�s�_=�&瀷G�2�Z�:��+��S4hs�� ���+�������I�֘P[L�H�Ia�K�*�΋#����1��
 �������T,�.��#(�_�\r\����|�e��M-�C��"�0���
.{\3�hO����h�.
�N�A�^Fxhq�,�j�f�y=��@�%�������YG�l_pk[7B��B���#����|�̫5j?�� �tW��k��k#���b�_-��#4#GKs���x�<�M�FIh��.�cC*`��P�\�V�&�{�P���ZP�$���R1]T!$�
7ɏ��=U�"9Rq ʶ���PLd7�ήm
@i����*d�ؼ��V�� eoq��A�\*E��Dp����u�XIx����nkD�ٲpKߧ�vA�$`\i؝(������7At��X�lTzhaK�l_2D'�KIjX�����~5������T�v�~���( u�����>��Յ(0H0�Z]Yb�lV�,!*E�@(����9X�3=�� /"��	��M��@с5Y�=�dQt�W��q���u>e�[QF�+0�{���p-�/ݽ{�?z,�&(!W�#Q\?��������a�!��T�1ݫ����4L5��Y|_(<�f!o	}F�ٻ�����-V���Xh4҈ �(w�HK1c0��(��� �7P$�Ub|a��}Wi�d�d��x͟��cem~F�$Ǚa%y=)�9�sY<Vgc	Մ�fv(�5x�2�Ax rӾ��2��+�B	��N��C���\�B�)�����A�W�{g���>yB���H ��B_X���
�e �� ��=��FXj�j�*X$A�����#=��=�Gk���=����kyJ�ךZ���<x.A �E�KJ	���c~(���)�y�^���`~��1�����}���������G��[ⱉ�2ab��e��kx��
��Z�[�������^��Yx~���S�t�y����+a��h����<��M��^#5� ����O"��޻���=��g_䪟9 ����;�>nѯ������R�E������x�ʚ��Pp�0oxB&���^P*y!�V@~�A�LJW��2!�2-, /TA�dt��($.W��x��ĈY��`�`�a��c�X=,: �����Z��`��V6�^hd�{��}�T<�h�^pz��5FE��k:�ݐ��[�7���� O /.�/�	�5F�8�$�M��]/�,��4\%0�Z��`��d��g{�m�L��E�Ęs��SNX��A~FW���0y��l�(�nsJ?[~8��1�U�gYxwr�H��^7:�����Gko�^���IE��Q�rV�����u ���um�u j�mcnV.S�y$�w=k#��Nґ��>g��V�����sA�҈�@�q9T�ߣ���c�VK
���!{���哅Gc�(y*�pX��j"\�ȭ��>U���X<�V�фu�a�EYGmT�W2���N��j�����<;9��������'秴z�"1��|� �
�6��m-�> CH��i�6�f-ͱ��R�!\x�P'������}f҈�\��X�%�FcJ�OI���h�V��*�x[Q��D]"�6���8+��o��z�5�ԋ �����SI.������,�Xp���@���:�.�'�m3���.����*�����)L�,DE9����M�4K@��pm��j))]bI���I.�VY�za�٠��WZ𖬁���rm�N%T���`��	K�&�$�|����=p��A�T!���P`mM��7I�k�]�%	�Q�����@Q�G���J��N�H��̸!F��4D4b1u�ZMm-1�e�,-���F�"Ct[r����"�"U�ȉ�ʀ`m�*��(WR�����z��.%��L,� =�U˫�_�F�ذRQMY�a�n��!+3��g�������KZd�oia^ԑ_9�K�"d�Xk�)�ҹ٘�
m_j�)U?�m@+�1���WRP�D9�uED�Mm{��Gm��[�ö�dq�t]�]�듷��c�V�`�����
o}�P8(ħ�Gbe�2����a�E�Idu�P�Z<�jZ�H�G�]Vp���?2`;�SV��<;e���EN+�����xb����믿��ÇBV��I��pN�
����;ZP~@�,�����3r� ���=xpO�
bc��<?�ڥ�<���k���;V��<X�9���:�S�p[��9����Jp�W&�Z�ƼBa�<"�!��;<���χt~2�Rث�@?9�C����2����;7"��;��	 f�H�'v���2�����-K`./��A\@��y��N���E���aHK�7��Jk|F��Xf%��%�����`����2*q�:�}u&
R뛄���//�38����@O�������((��e�|f�������Kݘ]�����S���G���~��/�	Aʙm�)C�(��1i�l�y���c��/F��������O��۱B��"�	�"�=y?��Ч�����������3�M���[! 6b���
��3�Z��W��F۞�n'=�^���C�#7�/���,]�c�:
��jg%����k�|�C�O���6����=�;�S�r�@��~qq�^��'c2?#�X<jʴ�cd��+	��ܼ�iq���KTueaO�_�s:���;8���g�ߘ�i
#�y�<�����l&����gR�Rz����S�7�wLO���1��tV����X�Ы&�) /�_�PZɋQ�ߏ[?�=�W�n ,)�
I������B9�!�*�d.�E��dYԍPTj�L:H����B�>��a�~���M?�3�xJ@��e�fA��G�y_�~�o)9��48]��z�0
$�@�'My�`}�/x2;ک�t�y#�U�ͬS�H��ٮ�%1�5��$=ud R��LOml=��*zʁ���)�gzq�?�"Q�d#���&���9�&7�C�DYo[�h�ԇ���1���VCcԂ%�%qSa,�:��/���:���
W���u��!���X9�sq��0��;�%�n�T���A�h:o�+n��d]5`5�J��ˋ�X���I��Z<_"G,q�/���!�^��Ѵ��E����+���.��k �ݩ�Qt�:�j1�l�u�7b%�@��]E�x+��0�קv|a D�VY���riԢe�}%M���,V�T���-?ʀDaM���`aȪ�I#gt���@V��0:�	O�$򢥡P�����>tb�m��d��4�bsF.?�*���I[����.6��z���A�̨�J��U��f�Z�RRfe�U����I�Y�A�g���$K1% ����.�����́4�T���V~7Zܩ��|�DQ���J{�罨���dI�u��3 Xk�9T�Q�>K�`�B�QI>�D
nj�Pf3H���� �!�WRc���a���q�T�����W3�������u奘ˊM�Lp0njAZSDn�P�hx���@�ݛ7�%dzwgG�?�!d@GqmL����6ա��
��ayk��SB��/���/��[��Z�7����ݼ�.r
�P3 ���>J���H�Dڏܷ�9G�*�L9���5��c���>|�'�ak�����"Y�o�xOj�!/9i(����7�;<1(����+�66�2ȁ���\�� ����(�xSr�T�hhU�ʱ�aB���:���S  ��IDAT̉�><>��_v�4k`d��js��P>xL�"�q�M$G����i�u_"���������bZ��gE9RBY9�j�P���r&#�X�����ES 2�oo}��Ľ�s5~6f�pK�9 ~c�O�@��9�q�G�Ϸ�W��B����	�-z�����!�O���ؒ���~ۤ�r*�ڴ{����x́IyA 7�+C!��W���6�7o��/�?io�9r��"��Luu�o�����I����x�n���u��<�x��@J���K[-U&�# |8>�?�N�����Z;wp��������~\Z��Y�3�aYý͸6M�K�YJ�:U�^�{�O��?߇���K�>�Fz����>������ 
@��� ��)�"E��3:t�G�fOBO<���d��鶗˽�k�\m��u# ��S��~�,�%�N���������*k���[��7��ҟ߇���ɢ�*W�9d�C��H��ȫ_�_kmڎ�ݳ�~�R��)��h6T�u6)Ps�iȋ$d�@w�@�r_ r��d��$79B���3������6�a6g��_�QCa3%�� !n��!p"�q̵�JO�ڣ;n���!�q^X��_<3��cd]<"����j{��y$�/������(�3ƋgX,|P�s�W����GÁ�)�8�:�Ѿ(lh�h�C�46�֍��2﵆[*�R�鸉�o�%�XD�0��Y8H�E���j����Y�!M��
��;QZ�~�����v,d8���D'F����Rh�Xs�E����?]4u�v�oYL�˞@..E�����A�cDx��K�k��f�����y��#��G�S+�,��Л�5�f z���������MD�ax�^���_�|�$wEA�ׅa� `�7SB�1!(2Ȳ����t,;M�R��(��o�kq`&�G-���l�"Fx5%��	���`D�<k�!��Q���X}�!G�X���{5A�W�)�j�W�T�Eo��8�-K�m6���fAeM�4������}X&��B���7~J�ؘ�ƁtU�}�����M�4��W�g�ʵ��p!  ��* ���B��)=�����<7��E����d5��n8RAV ���p������$���:�����'��Z/ɳ����>6��@�D�$����
�1x��l1�f�Ɦ6_R'a5Su�5W�̵tΜd�p�}cS���fundN �}���fE��>߉qĩ�y�t)�:�%e�7�ނ�Hk*�wsxX�/�ʅ�g�4nd�|�2�ӽx ��H�8�&I��Sl����ԁ͏`q�d2�� )�h�� ��������q��Gm,������%�pNKb�nH���a�E#X�����0�U�#��f�̴X��9����l�N���J�b�l<J��E�������;G����D$B>1h�*A����9���An����$Փ��QN��1���L��;Ⱥ���-��}ׁҍD����]}~���{�{f�"�؝Υ��i����i��}�u�7�Q]�?�C�?J��$���j����pv"�9}�w�l�_		�Ή������_>�_��B��ؐ���ԁ K[��%Aѻy����w&�)�\��^�3X'��w�}�ipMz�}��cY@������C�˃��a��g �SM��H�F��`�g�Ʋ�{�ݾ���W���??t��#����?�[�)>�S�e\�L�Y"<\���ï�j}�w���E��x-0��ƈ%�~�ѥ��,̜B:Q�7��tZ4���'�Y�!�,��z����a������]���Y���=mo�hs����j��\� ��� �i�u��~����ׯ��펮��r��QIɬڠ�HV����y6B�l���'6[�M��d�۟Yޅ͚ı9W�#^ &�O��ϰ�B-h,�D���w��o�Z�b�0�N	�]�C��W|/�����W��S��[i1�O+�L�^��ɘ��J��3�T��T'����#��Ԕ��X�7V.����L���p���T	�ſ��
j�ɽ	H��A�`aji�����Þ<N;NF��D��a$�ﲂ�}�o.�qfv�ñ���z?��/���fZ�.<�1t�+`ⴘ����T�??p4�=�.����x��w�~�$Ju��B�F��\�Kt��L��F?��FGv��(^�XM��ه�kUKך����~�&-������=��~�W�*v�L�/�Ҿ+�CW�@�/�-Dd�s�\+�pj�՞����vY�1n���wxQ�X J�ӳ�٘�ٌhX�Xj�h.�x�f���U$݅���F��M��޴�����S"�|�Xr�ݫ�Zl>�}ZPȦ��M��/(�
�� ZF.��~����`ƟV�T��c S������X�<���c�j�F�ؖ�T�E�z�}]2��>�5ፊ�@q8�� v@Aafe�B|�=��b�p�M�ZDk����Q)*��unI��Aܱ��'f�c�0w������D�W���`i��jS��ҍ���Z]ܩa�
��������(�����[4����ɕ�r�ԟ�k�WB�`m�`.U�#�l��-�aQѹTZ��Q�b�
�ES/&�8� o��:5\��?��0q�/����:r��E�
�h������?>B���!����h���oZɌ�I�e ��gC�C�W��0��8hq��!;	���e=�,fB�Z&���Ͽ��s�A�F(HLB)�:o4�5B3xc�~k��j�/6��be�b�����-1[������ sǇ1I�q10t�(�F[g�@y�� ׶Ѽ�����R�6I��(���P��@�n8��2�?��Hm����g"��v�y/�5���9��鉃��b �����s�K�_����h��e�P?I�������[YR#Vt�ǯ��:�痝b�KϷ�4M�������`Q�� �˥��;�p�׌DF��m?G0/���r��e�Ao�C��{������^Rr\q��Ԕ`J2^f�ʌƎ�z������i��37���~G��=�������g��׿w��W�GY>�"D	d{��������B׻�~yw��у ^H��������ϞӜ�|�"��3;u�n��w��92k�n��8�"VXK�� ���紶�l���Ѷ8i����D��|>v���.wؙ�v��5j�����b������+!���%��tIs��h�ns�ן���,�e�:���,#�S�3��
t�69\�	�|�?f�%| Am����q���
h<8��b�`h7��W�(`5�O�9ŀ�ܦZ��r�,���;�|��-�l�>*��J�\K���e(�l+a��R0G3ta��S�d6�Mj%��f�5��i�'��Sƣ��K��_�u�����>��^�ĵ$����<b�[�P��i���t(+2�
'�T�\�BF����!@�5K5�GC�g�õ	��I���׃��a#���^���кy���9�_���rz�k��ه�����pE�},w��h{d�$�^3�9Ӯ��=�2���KZ�W�hij�(JzH.j�Ա���zE��#��M7"ľt����.|?����E��[T�Bg�۷R*J5�m��`v�S/~U�mp!Mn��v�(�C�g�����2��i���BL�%�7���h܇g�J:L�t`qV�`kV�� ���h��b-AX�14Xr��J#Z[JxWdY�4�� `�ջ[b3#�^Dn��QmS^��G�_�x��⩃��^�R�bϘ�/fM��FyL����rN����]���QxlP(���\屮���n �Ƚ�y�UYrt��$I����0���",Ni��I����}7����]�Ԩf�ũC[6^�ĩ9ӹ��Zl�m8���f�r沓��ٚ	+�'i�`m�lM�p��5�s�5�����k�uX	Izc�lAn�P]��lk��$��Jgn�~��P�9��^ ��%���t��KѺ��|�(��pf�UW<,�����Z�N�L��;�R�E�M�<ZƆ��R.���̕D2%���h��?�O�����z	�@��в�������{��	R�G�b�F#Gy��D啂f���3Zj�*��^��"�d햲,�w�5�oU�B���s��2��̑�B�R�d^tN`�D��1��/��IH[n��Wdq�!�1m���T$r��N��A�߾�g7����{qH0Q̾���^ +Y̪{<M�?j�M�<�%�L�Gqx�zd �����Hth����jc4�[1,ذg�;�X�y�[(n*�`���;}fq���Ϭʾ�>JB��s8��h�X��<&ֿ4h
�}k��OR�z>���( �jx-�V�����8s�$�V�sa���T�����mצ�;8����k��O��?ӟ�����-3��Chf0���~���&:��>S���Ӟ������it����{ӟ�H�o6���+i��鹷)�������Dl�M�kI3d�.��|"Mc��
H70��Yud�s��͍�$r#Gy�3�������J}������Ͽ�����?Gq|LS�����i��|�Z���>�L��ng�^��ׯ�����;�{&�8K��I�U����<%e�H�0�9�(�޴��d%v���P��0���f2����l� ��j��@�f��9 ��Ek��_��F��Lq�P(�_ �8Orz&8��ui~�D�^/ca�t�mR��"��q�+����QʺjI�����>-�*���Iv��oώ�D�S���6J?�^4�˾ی�y#����h$��kh��>��$�/�j���Q��� !��Kۈ��.g�p\[QL�jWu��٣�!�2��\����$\P�b+���99"�=I8��s�y�P����٣ָ�y�ǳ����nН��>���p������Khq&��	+w-�W"�+"�5'��Hz�����#!r��Q#�e5{"�i����.?���OR��������p���i��B$"�Y�k2x�6�7�9E$K�e�ۣ)Si�j����n��౲�ɣX���L]H�b/a������N�#�q H�Hn��s��H�� ��=�@�K@e�C9wp!ilO�i��)�����J15��`r��hhIjp��z&��,m.�O�fP�4��,��7&3�0�X�](p:$�A��dGEcuX���B7�z�����������������j��*���7z�=�{a�tP��Z��
�H�9uP �>LM�����MQp���d��R�r�{e��f�I���'U����S7D�U���@�� 
�k5�d�����Vj����Ϥ���
�{U��ښW��1�"7œ���G2���P�\�)�#�N�2 :YT�A�px�Hif�7�93
���WС��;�O������k��R�l�� ��=�歹�G����j�Ǡ����Xg��U� ����59r�ԯ;��Ԁ�ApJiU��N�A���|,W���d,E}�P��Rܨ�D*h1:'�{#@����qv���tv�#���nS�HWUֹ���IKI�T��f�Rŀ��i�@��Y�l?	��6B�>g>���8G��D���]w�H����O��G�
�T4N�UgA�(;oΗ&�OH�6�y��3�t6eq�.���(2�Z�7 "���h�~m���Q@ܤ�N�R�u>[4?׫�[���ΧA���4c�_B�"}�9�&�7x_smS�t���$�Uk(H�,�nN4)ʬxl�X:O'e/e�K�����@�����~������~���Ы77⼙�6!_F�a?�?�s��G�� 돿���?ɹ~��?���}�#�cx?m�o�N 4��Z��2k�-�K5JL�5��[z��{��/��/~9E�/?�W�'9�~�w�����F����~�H��/��plt��,6��rK�� {v�tJ��[mH��Vk���޼y��o�Ї����$-:�Is��L��l3��/ dY��Dg�>8��;���ȧ�����l��o\���J��H���0VcPf%5��$��:C�7^�+�FS1.�*O%㥗}(��"Yޗ�%|	�Zb����MY��<=Z��8�->v3��[+a��q�
'�}۾��H�0I3��������R{Euq�@��Jq&fՍ�'0b��]�"��
x�"E��l���B����nb�I����E� Ā D��1�=TM����fP�{����/Z0y��y�
�t�3{u�����R��7�pwGGk�'1a�:K��x(��=����������j>�Ë=w��k@,���,5�u�H
�� �5�� d��r����/7�4�9�>�n��d�bk��,mR��H�μt��O3���
:��Ѧ� �a��9�3+�Z�Rf���-�nx������M0 ި`�"Q�-d�~x��Pý�u0��@ S��)fٓ���d!���b
#��c*���󨛋Ә��E��ż�&���N0�R+�tq$Xҁ��Ʀ��P��Р��������F��Ʌ f��\����BANzD�8F�� [�3�jQ�:j$K��ɟR3�#����wb_6ݰ2��,F� �͛[!���w{=Юw��F�Z��k���l�����K49�J��zI%jVܯE�*hD�ܘ��j��c	�Z�ee�![�𶺠o��DI���ãʎ���!��6��!"ZcA�x`��g�Z38=�^ӭ �Kx��F����=\��}����"WL�����D��r;��-��b)A��5��ا>ߓ5��Z�4�V��=�>P�8S�V�,��jT%�7]$j�^i7H-�ϓ�Ċ:���:�~p?�dq�O?̃��}ux�2pq�.�g���@��x[��}�,em�u-�z���$/_,bXl]i]g��{@��ϟ���G��9ʺ�te��ȋ	�������˹�ck#��$����r�m|<R�w�T�&��BU�UЋ�rNATGZ�y��<�U���O�>jt4� %/%H��A륙�X���쪓�]w�@R)��5��H��4RVd���R/�=�w"��)���[z��D��m�j;p��>���p�rmӯ��mW��?��?���i:.�k��k����O��%�i^/�+��e���܊��SLPss�)�L� Y9��y���E�Un�o;��N;���h� �kp}��<H�λ�A��8-�K�_�l�e��./��k���f�dvM&,b3i�c5�ʨW\J<�����p.n,�����&��[�5��k�_3Y?��F�P3�h��dz���)��i����+]o�~��A�Gf�M��"/P�$�e�L�\���nYA���?2d{���3����3v����_�.�邰����78^�
�J�lS��<67���B����#=�4-��3���'��fmXk�p0����J1��rʻ2<i�:Y�	<�n�"$�>2��6YH�m
i�J$^�QH �@؞�sWbG��6�A�]�����P�U��)s�W=��x�t&��Ȼ>C)[���/�20<�j�L�fL�.iq'�1��3Dv>�"��4G�5=J��� "=��'U�H�)5"@���ym5�Q�O��3�*��E�XT0���/p�����*���" �ٸ��p������pQ�Y9���D�#��$��B{@r j���b #��62?	[��`lN�h/Jà�FÀTAU���J)n�CQo;��[�7���s��0����M��s���H��#N�H0��yD�`�Ԋ�|�k+b�P�Ԑ�ؓd^��ޛa[4R7V���d��쀪D��T�ԋD��ջ0��JG��bg��U��I�����k���ry%ulL|fB�&��k��� ��=)kb(8t-9Af�� �����4=���nyf`�+�d+�(���{���.�)3�H��2�5�c�;_T�{�twG�t�+��' ��֓V��ƞ�职����=32�g�D�s��K�M3^ԁ��y�	E#��Ob�_��j4��ҵ<K�*`	5�x��l���&e9���:��I#�7�q$�.I�z=�6t�EJ>@h.O�A�T)�rP�6�-*�~�^#fD.����ߋ�ІF��P��T��j�.7ZGp�y�6N�9u9*u�耋da��;@u_$���S`��P3D5P-�Utv�#�4r<�b�Uu��9>]�1�N��� �jd���u;�ѻJ�r��PN�Q}�Q9�$B��j�K�7Z暻��[ڎ$�r��d�`���JP"@�,)��Q���?|O��o�F��AS���6c6ع���ͩ))��NR��RS�&Z�Ek�X�����)k�~d<>��������������Ҩ��w�������iډ�Fō:��gà�$N�42)��=&���i��9�h��f�Ҟp�N���4%Yp����{���i�ѶŖ��r6<ۖ�3̖�@X���(9t�v\��ٚ���t�(�]ƸЎ�f�ȋ{����+���������s��-�,�ګ��~�5��ZO�ث�L{�8�;U;�V�J�Ɵ}|{տ��#����Q��@�b�7�Q�ƅ\�C˹�� �	�'�e���F�OA���By�o�^N�C,�Y䛈΋v�,�X
L�j K<g��$1#��*�h4���I*�Vu�p�E���ffZYn��78�w��I	��q�T�y2ᥑ6�J��,�
5 ��
���C m��եM6W�K����"�iιQ��ʗ��f"�Zʳ�HV�6V,��H�J��Z#.�q�z���ᴲ��M �`(����2�ūx��(�� �9��mY�X�fT��m��I�,V���l)w�F� K#M8.��"_7BC�qa`��:x3X�`Ăv\@�f�j�`0)ч�_���I\�1i^�F��p���W�9�+�Â��g��w����+��*Y0ގ���!�yb�В�k:���i
� A��lt1������sc���r�U��3���r��*\�O�A�?�_�|(�	���L4��&�I��.��SN�>�ȯ5	L�՚_&�٭(pm����+s�n ����ѵ�F�U�{ehp���=��?�i�2� K=���2����-=�pZ��{�AOӵT���D¦9� ��Hu"��K�Nѻά]G�f&��4��Q��ƴ����KBb��t�N�k�T��	�4�<)�{�����H���ِ�}�g!��?:>��̉�C3�Tv�<�S&��My��_�j!��T�Ct]����@dMf�>N�f)��'u��b�Ҭ�],�y�0�����)�j'j����2~�6I�0l�p6��T"�p�U����Q �D��� ����S��R_�3P�D3G�d�Г0�im���J�BAFƬ����X����me��z��wh}�]Vw�}�6�{��7>M���3"I[�쒋��st鷿�-��O�~���#�߲��l�*{��֢�ɬ�6��F���I-���ZC�i�l+}��I�7�e���;�����W��O�J���t`��#�B�a=�xl�ʖ�ҫ	Iپ��XS9�h�2ʤ)5j�YI}�1�����!�'�N�F�)Fb�,l�d�&��ζ~��#&:������grV�RE6�؋E�r��#a�d�ǆL�Oj�l�Ȳ��}�9f_�n)�8���`p[+��tP�{X}#^�f���f{,����H*�{�9����5�u�G�i�vB�\.Cp��#S�G��,�}J��d�<^�W�s���Fu��F+�lS�;@r6+eĎRoS���D���D�D���Y�=��N��g��JF���"
�1�'OG�2�M(�B+�HX�=�O���N��u6��� �d!;�g�2�)bF}�s<�t����D륤+����nV��([�EU�
3�̈�h�V6��ї�,�6/ܴm�%��*�Xn�f�xj jK�䝯y$�$-�<zs�"�i�:����Ss�3R���f����}����.Wf��e K"VÆ�r��q`1�r�eQ	Mo��8������H/��M���0Y~�p�ų%=j֜�	 K<���g{��u�XA��jQ�3E?"�T�2fC�(�F3��H�ٌ��m����^bh\v;�-lB�@�E��^X+TN�@�f���ԏ0��9�wc��'�W��#�dt,Nb�wC�[�RH.b��p媠�Z�P ��T3���k��`��8��y4@1b?cA��&c�~�� rK%�{�� �2]0�Y"�3�d=�h� �@ `"8�,������Q�,�һ�� �^�5��E�'�!6)Ϭ�e�ً���d�{��0��
p��j���-,@�3�~�B��aIg�@�6�O��Ig����1�k�8 �ؐ:�<� $Bđs2� �Mk���u�5"=��5;$�\)N�$Fh}!5\b�������S�ST��Պ�Fn��.�@�"z"�����1��Z��sP��X����OY�TgJn�^�����i���lp���$:tk�}h�����1�
.������nNRw�La��xGu��c��6h<[]�<�4�>��2i��(���������ՙIm �]i��ka��¼XrJ����tu{c��B����R�-1�fc�$r*v�R#�����l�>~������&��3Q3�>���a�-!���]W��k���8S�B4�`������gЯk��}���t�
C���iy����ߐdL� ���0[�f�-^�2H��ʹ��@ӓ�?����k���#1R���j��x)'pȀ���{";�ln
���}f��,}帖l��~/.i���L�����\������|,��jp%@�^5�+�`��9����g��������B�~A�?>"�w��#�xw%pb��:캬͐��{ڴ~�Ej8.������1��u6!Q��w�W2�#K��V��f��ӣ��� _�,�ZxX�ޗ���1�64e�b�Z6��2iL��׉D�q�u52I9�^��עobr���.��Y�ॷCO�"���lرTcSrg6�'S0��ۈ" };
%[=)���	H�a��lYx�����3ij&ϝ����>l@�Q!M#1c�<��)*��f:������g�Z�۫ \�W�Ak�O�\}��髯
Y���&��F����j��e�+/(�*�K��,4�k��y9�t�i�x�`����E%���ה3�@�/��W��e���4�1[��c�S?�G�4BaS�G3�������=�D��hF��z'�X�D1̩���f���t�TE�T����-�O��*����^�Q6NK�V[D�̶��D݈`C���?�Զ����ٻ�[Nfl��*{F'u�ؼ��
5[��7��f�u�bc~����WCY���{�5C��% � K2�y��6��l���΀iW�.���+f��hf��H�O+���S"?R$\b��&�������ٞu�juʑ����	)�� �`D:N����PCY.IK��;ZPrOБ�m�f���F��2�fn�G՚Q̈� 2��!��R��Q�� -C4N�#U�$�ȠP�+j��p��B��q�ܒn�<w[
됬�("
:d����9�|����?7�d���C�3���>7S��YJ�|��;���p֕��"��,���>ǚ��L_b�A�pa$���S���֨R]��Z�ό����*p��׉Yt��]H�@8ⷫ�4�g5����˟.P�������׏^��[����n��R�}���)ά�6r��D��|�}ݝ������ N�����=�2���A!����s�������>G�t��ʞ�z�q#���������'9gYS�{��^1�F�eo_��v4L��m��n����n�����e	}-�m�i=q����HvW�F�����n�js+{�#���{���g�������5q��R��ƽ�s���א��0|e�*��2�S`�d[�����d��s~L8���p�k�����QkUf�_ (K�8��a˧�P[O@cp^�߰������L�;( +!���'v�ۑ¹e�ε�@�5���q�ؽ�6)"���OC���l*���P0w�jJBܪa�0��sVK�.G�� 발&��Z�⎸��@��Yd?N��avU��L�}�&����5�:�q�G��f<�<�aa�/U��E�@3�vH�0<[2�9yF�<~d�6&g�,x�?���a,�i�~�?�d�N4$E�ض�Ľ;K����h�k�z5�axM�V���45H�K($�bQ��/��C���@Ϥ�K/�	�W���E��W%�+����3R��X�W���� cPfl�x����(<��蹿yme�0!36�ʢ䩄aiFX��.�$����%��D�Jx� p�Ir�(�Z�)���H,R�Eb�����z���9�l�����)��%�>C�x9o:�5s�[� �v^�!HB���w�=�%lS��R��zp.��b��-Gij���Z �g��tGOg�2�qc�����r��w�����K�r S`z��_L.�ΌM�:�S���Y$(/~x����"�XyP�n������>&;�.��
�sA@a.C� ��E�Fe�O�W�c�.��~�w�~޲q��|^|�p�Xg�e_k��$�t�l>#�tz0A����������(�x0��dcN��(��g�����bbk�[~�n�{/��x���j-KQ�$�9M�B����/W��������Jk>���3������z�s��Ŝ��V��zY	J4�0j���r5�/m��\W���"+7�����1<�C���,�������΁&�����;Lf'���ST��.����.���i�y_E�@!�4���������E����֚*Mu��!�U�^i�����o��;�t��\�����n�9J'9�G�-��Y7܏������k
+�r0P���^zLt6[��F"���{*��܋�m�אR�C��j�mSB>ۛY޺�=��l]3	��K�#U�Y�NU�#��_��D/0spY�����^t�%�䕧��Op���H�s-����i�*K�xn��j����0�+�4Q�=G*8"��:��W��^h��`[Q�!F��RS҄��N_q��ǝ�ǲE8Z���2a���Xĕ������HX�b��ٌc�)�b��6e�����O�5I��V.+i}�F�b��8��@�_�_���	E��`���jot��j˥��������ym.���\F�\�/1�νXZЀ�[�l�n4g���^��D�=K��7p�i9"��S<�Q�bf��b|�FKT����N�=��Ȍ-�tt2�_e~R�/^rI��������9d�ژr=���̾���j�JBek�����zl,�F^�.ml�S�}�p�	 %y>d�䖖FdLY�ʎ'鰳�aJLE�P�&���ԧ�g)����q��F� ޵�]Y����G�D�l��ɒ��}�ȣX�
5Kj��>8i�%��\ �gOaӾD��~��	Ʌ�[n<~Q�����}6��#�Y�[f�N��֔�;M?�k	�i���y�_Y���m�ձ���}KO��Z}�ϟ4��`��[qG�̔0h%��#Ҝ�/��\��4��}�Q��~�9�{�2�}O��qkdqy�k?X�q�uq�����4��SJ�#	']xB��i:8V��Gs�`�'�	��^��|��R}��׌}a���ƫ��W?M���)E��E?����c/ғ�HM�E�O;	K G ��@۫�v[�m�g���`��?����ʺ��dZ��JM���rwG~��~������]�y�S�O�=����,̤Zfa0D� G?�>��I��؁Չj9e�)��}\�Ax�E�}�����~�������[�����G�gg�|B&���.�9���,3{�웦v��1�}���v��,�}ΔZ���a+�L	�r��µ�R]��LSote�C��RD&���u����3��o�/����p���mip� �麒7�}C���R�c|Iqԣ-]V�s�M�#�M�B/��L��`�6��o�8n)c4p���x�y?%�������5gcK�G7�d�X|2� ����V�I&��-&d�TQ꼙�i������pV���܅�
0֊N	9���v8�·\��~KE"1;�Ӹ��OV��i~��/g1b��l���M��Aɡ��d�⳦��x�� ��A	����\��"�I�z�T��mo�e��H;��JO�T�YD�TI��ڛ~?�Ft�G�D&��V��!��`n���I�d!*3�F�1ҵ��+K$�_gw{#�J��C�r������E���E>p�_��.88"���P���D���*--�un
]I�pi~"���J�+׌�������3lL&�LR�B������|��|��oi�Լ) Y6��J�}K���2^�.T@�^�t�ev=���`\17q��/�Y�}��.8���Չ����1y�)�Yh[4yV��Dt/ʨ(u���W(fpjZO��q큥D���D򇅯��]*ך�'\�O<[�����H�_&)L�TeR�HK��G���4�.���-�[D0��I����R[����*�b_��g���s6��,�vh�k�0o����6ʓT��#ti�����fD�,�dl��i�4��! �5y3Q��|-�?�-xώj����,�V��b5pN���j���*�AŖ��lu��0<~�a7V��5}��~�||e�o��<p5��u[���+Z�C�|W}&��9b��="Z���͖5Q4sF"_��١{�6	�P����g$?���6dmh18�HY��#��>d"��`N\�p8�݇_�������u��A"�ls07�z)�����%,���b�$���EK5��b6���R�z3R��h��m�o$���G_�'穃A6y^������3[�ՠ��Z�u�����r�%5\9u�k׸���R�	ӖN͈Z���ľ�E��%J�j���j�@�꿼X��5l+r9�B3�e��-���� О�@���W7H� �%;){�Rʵ�i�_��g�웬�s�R?f}5�m�C�>�����
ף��5"p��<�Z�P)�+]��,�`�V,�u�)�-�JmB/�R�:��Sj2/֔w�HV)���晥*[-����R�YTl��@K��p�	?K��DiVxu�
��Q�u$"e�v`j^*R�qs{K�߼�%�f�m��) Y�l�g{W��6]�p�L�]`q/���\i^&��dF��Mj�ظ ��L�q���Ak�T-��*_c;Ҷ��7J����4��_ǣ�0���9��j����o��Q�e�"c�Hg���g������qcR."e�.\�R}3���iZױ9�2���� 	i;$%��H�WG�� Nx' |YH	=/��C�o#O6��n'Y�D�x�ڬt�)��.�c�֒aޘ�
xYyͳ��7p,%Ad��(���$@�s����� �4~����Y./?Vu!	���� ����l�����|�gL�j�TI�[�9G�"H�~&�g���:�'f'�-���.��� ����w��[��W�ܒ� �c��b���(;(0�P0�~[K�����3�K�Y�'p=�PZ�_l�O���=5r�2�T�EW�F�\�hF ��{G"5�˹�Z@'��@v݈,�C��� C�̇|�����Ն�/ Y8��v1 kyޗ��i�U��8�r/ޛ�KIp��o�`�Ͻ�o@�;�(���B�!�]�˹Y�Y̪���<X3X���+�Ϥ�z�nv��:>^��� ���C�g���F�R�bĎn����qs% �)ݙ���������{���>9]8u[�ö��yRL�KݬQ{N��cc��J�������p<��R��A��7;���O�{����>~����7u@نm�}�?��ǩ}�@��Q�R�~c�S<���Ie{��jE������ck��[\E_m4鷲iZl���ģ��N�2�y���n��lW�%��K�z=qO}��t�K���_�{�X��~���u���!����9~,2�}I��	'�G�Ӹ�=#d�Zk^h��W#PMzAj��b	!V)��b��RgCE��0p*�mέP�<��]�qc�y�T%UG PHA��;�3���������w��/=gEq|��7���v"x���N��"}�8ב�c^�^�u?�b#��,����ة�,N��T�"� h�q��N�p��+bVV'3���_I�ُ�-������]�F��
������'���"BdO�f��mh~�T?j&��U��4�ݨW^ݬɥ�h���kƁ@M�o�LR~MKB���l�Qɷ_m��ePc5b�Sr�������o]Հ����^�d�-�����u"43��9�c�� >�euN_�n���Vg 43�
%6��K����s�́����Kz�w�O�x[V �#�������3�f�hQ,*�,��~[?�����0~f�*iHqMPW��]�cPf渱�>��20$ XYY�k�۲z�E3�k ��\��$&z��0�Xq�E: &�`�Т��T�u�gJKe�~[�z���S/1�(R\ᜐ�# �9]���UO� y�7�_Ȣ�I`��@1y�e @��D��:�b߈��Ȕ��"�|5���Q�C��E_�~<�g_
�J� ���X͌���&�28�f/�p�Kk��Z����ۢ3��뫼̮NN��>y%��F?�웑�m-�ϩ�U�.%ֳ�.	+�U���ݾz%��fk|���Y������5��R�$l��q���y6��p���8e��������Ý��d��ӑ�rqKvƾ�7�[�O�H
�Q�W�=SN��,5f��ݽ��\��� �gϬ����L���;j�5=�f���~���=}�l�͵~��DSy���3G���u����]&�M�m��>��/�t������������>7;���0��֩�j�D��7�!Mu�p�@�������[�b5y�`ľY��[�/��ao��V/D-���lz��2�x�Cǯ��}d�������M\B��k@��w�	����vYLq��WG+�[b.K���p�%���0���nB�Q�7M/TlYld�:���3պ�	l�M[�h�"�`���RT%*�ӼDgs ����p%_�~�`"6�A�e����4�RA�h��t0g�C�~���Q\i�(��ז��J�}9{(j)pQ:hUL�J�����?������7��4��w�EX95��bv��}rcW����r⽲��`+�E1�E��lk��u�y3�~�A/BX�mQV�d�p�����v'�O/{%o��t=�1* �0f�33|�GX3#?��p+����� �ആQ��<P���NѪ	@���r��Z���4A���D��>e�oa��t�z�U��3?sS��ML�V�s��=h�m����{�I�y��!��grD�X��z���'��xj��0n��Ϸ@��3�t�PH+�ԣ��k�`�a ˭K�:�G�P(@3���5]<��"��x=c�_��9Ӝb��>��TrƄRn��+��̴<o�7�8"�!���h��a�8�K]�=�Z!ڊv�!ӞeM󿗢5�.�6V=�?���;GB X�o�,��랆�ќT��l�c.��~m/,"�Ͽ����BJ��~�k_Q/��놑�p��6�fo���ߔ�di�P��h�)l��k��Zh�Y�v��oz��][�rΎ]�=ą��ʀ��*f=��%N2a�4�A>3Ď���'�_�뿄����_�Ç=}��ȹ�K��h�Ӆ�w���+���M���<qSa�v{`2 a2�H�a~q&�A���hC뷊�>�޼����4�?���v��wwCu��v��~�t#�,f����.ۍE�L��w�hہk���x�h�o#��y���͖+�ֱ���T4�C̰��F4A���N����A���{�%�}n�'�υ���~���9fm�@w'���6�|���;틗r�M 7g�	���2�r{½U�V�߭�o�k��*\[�֊ke[V
����.�� �Vq�*��30*�ƺ�_�zi�e�Fk�(y�~��&!B�!ۏc[y�%'Y�F7�*�a[?n�������� =��1���x�6	Ո5�ZQ#ɱ��9��p����4����W�]��.�b�D�6���C��W����׊q�L��#��$s����=4���B�1�Y��k��g��q�?�_��.��5Ee����\S&5b֟K,"Ͼlcx���5}"}�����e��Ә�@�믠!-�A]���kzO>��X��Rq�7^Ki�2,꼗�(F��ϗ�3��m��!����R��ĺ��i�����@�O:.�nT̀)*��r$q�$ a�7�7�>i�� x��2~�{2LKw���A�?�֤�{8d���GjE�T������?>��16�(\�b5�PI�^/��F0͘O���^��hq.�z�d�����������t%��۝��9���;�i
��f��ǎ���3��6S!R�́Uc�#��
[�Ѭ��{�II�4tUq=��c_�!:������C%��T��龮c!,�"	Z}yx�֗C��Z=q�1�=�"����Ʉ��Ky��Io=����O�/m��Ǌ��0*��ތ���9L�%���J�F�ƪQuflL���\�
��0n��;:s�vQ]�8�t8�����#`�y�N��f��rՁȅ~��gz�+��t����^M�;:7�L�ǠuNu�6�L#��{�s�=4ay�(�T�ڼ��d���۸� l�����<צ��������ˉ{���Վ����U���n�]�T���"��\G�j�yg�.#�b�L��E�.�mƠ)iJ/5[Z�U/�Mԃ�C�I	A(CԨA^�˺���P�2ÖY����u�Q���ٷNa�Q5�,C"�8V���F�����`��~}|�f�`}��.�R>�C-��Gz#2|п3r3L  W�^��<�C"7Էi��)Odx-縤(VF-@���o�yi��ت��	�+��b^����n��J�8E6"Y�m1�
�u�Oּs������SI4$�S����/�|������r�y8bé~')����" ��j1�`�8�(��'i�)�wq��T�B��c�%����sށ�fT�W5"�(Q�N}<'���Y�5g�>���2dʠ�t8ҥj���i!D腣��Yo��&��M4�J4kF.[[�oL���KEIC]YM�i�Ya�6?��;,�LZ��F��ی~xu ����#Y�[�Hx�+��C���YVܾ0β|�;_�ׅ1+�!Ƹ��� C]P\�u��y]{s#�g�����o%L�H���.���K�V#��oZ̑�����L����=�-Q�%�Q/��If���j��C�k����ЬY(�@��\S�SI����1%��Φ7�j���RIs�s��!��W��W��iYCZ�-@��⓶��m1z���6���A�os����4��$��gfK;k�6g�h"�p@���FX:?9
����.פ�a��,��=��gq�4�b�ɢ�A�K���K`�׊�����eV4���DgjQ��+�Xy�|BN^D��_�4׸Ƕ��8�e�����s�~�\�1���|��/&C3]�	0�~���&s�ʈ%�n�Y�������n�k5�'S�a�/�`Y_�tw�@�����z�A��~G%��:p���{�����2��)w‘�<�jKĮ_s�2���H���q�/{���FG�_�7I�)f���ҹ_���0�E#X�F�X9S�<��@��;&+G�ͩ��-������5W4��4p�j6,�7�R`��s���[�Bp�Y>��=!�x��k���"0`UC�%y���A4�/+��N�4���y���w(�~_3�� YvD��Ul�;J����}��^m8�w��+=w���?!��#Yf�/��������$�4T�|�b�ػ���0�w��`�|�Nq����'�$�� t�D��2v[OC[��l�Yɏ@��<���|�>�J���1j��X��Mn�ť"�xC\���m�����E�� ����O���?�g�%#�����Q�<��oN�8� p�Z�79�@��>Cd�TMkl¬7��� �Z�l�'3N5ϹM3�Zd�?��;s��dr�QG�[e*S9�d����v��q4�CJ��|�ד��^�,M������A��+��C�������aa��z��Z)z(,ms?����'68��kk-�[������K�N�uSY�������q.=^��-���)�<׃-���!y��i"����3�������|f�����aY}��vȥ��ڕ�����j���$�yB�]S�渺@��5�"9C����Z-��$� 3�|��[(���N���7׶iJ���»���_&�f��<�F�Y���� D=J�Z]����P�8]5�Q�tl��NvM5�[S�=��3��� e����`�䵼02J���ri�Q,�稷M�k�=��ј�Z�uʨ}� ���W�l�X\=�Ș�${��\��笯��fY~u�2zՓBL���3kV���d~�K�KF��u�;?
���Rt`q��(��e��C��w�'[G�,�#4��#��ǚ5��e�e���wN�c�.31֣��던��x<	9���$���~߯� mT�=s�Ij���^���L�>0�OU��v��{�ƿ<���@��Z�]����X����I��s��uWG�$T�B�1rM�e�A���N�}֯9��z��Hֹ���[���H�9l qW�bByv"�&v�$�zj�t葴�IU�d���󓟭^z����E���~�]����}�Ԭ����������N����P�;!���P�6+����C�]��S���;(�읭dC��#R	���C*� ,�p���V�m0|F�Y�&V`V^��t9M%�����&4�r�5HR4y�A\��¤$���L�ߵ�T��_i��,|������*1�����
5f�aA�-fku��?���B�z���6IZ�ty�s9��c�5Wωe'5c���{_��2�f��w���#�� D�LA X��W�G7��-
��[�����h�b�!�A�;���-n��4�@��ECdPO񅻧������<�V��~^����*�i�a�\OV��=`�<���H���Ʀ�XD����㴖v�1-�Zl���G!��`������Abѿ�j�����xH�bl��Da���d�5W�P�޳�����s^(<0������焒�!0cRy^5���X ��J����i���"�[�6'��h	²r�A�����e1\,�]�?AG�(��VN=���%��raKB������������aV�)C�7x
���} �-�·��k�Ҿ�Ɖ�b����j��,�4���q~I���MB��x�1��pK��᦮��F�Eܫ��bOD�1E8��x�� �Y���	7��Bf N��Ʈ��gc̆:�MYi�n�����XB��:�ůz����QU�"}�GrJa��0Vw��,�v�$Q$�̄>��f�,���:a��cL�50���f�ۆ,bC~e}M-����������QS�4�� ���L{��s1�v���%������J� ��ܴ���]��?�G��\=����27g��09�+:�Tw̚���p���U���- �8��`2'1@���M*cL/k�RԐB����1p2c	�}d�4���z�8�����]�v�0���e���ϱg�x<0�n?	�����6l#:��>��,��_��\Ӊ6ӡ/W����Xg�������u��;γT���]�үה���y^�5���
�>ڋP��х.N�k�� �T	2�a������z$}#�֐G�ڼ��dl�dz�@��W���'���j'Ք����Mqc�[��۟�gg8��[T<��~>�N_Ƶ���5R�P8f��^��j��u�7o-�,� �oBo�mm�L����yK�d~x��^�H���]>�����w�2��D̥ޫj��oM��d��d�p�����бԦ_㲡�-�ڌ�N#"h
m��Ƶ�,1�Y�qCPښ�O*�m�P���	�w6����h���z��,�o��lƢz�����v�ܼ�V�\Jϋ'}o2�*��3��Rh!Ȱ![�i��<Z���)��R�V�5[A5�h]jd�!�k֯KR!X������E�PmS�?��� D�(l|/�/�t�7�1�o.P�N��,z�h�)]��g"h����o�F$]ϸ�\�����=�|gAQ�EV��V����N�����w��kϏ_�!�1l(�ed�$E��s�Ꚓ�L7f����X��ă�ZknԚx5Cҡv���� FI��>���x�\�,p�{6z�^�a�<g؍�((����v�B�qv�E�T(��Oc[�ƪ2J�\�\aد�Ӱ�� _��W^Kc@d*�q$���-IS����xB�*��� l��gN�"�Β�G�X�PÚ \اgg���k�M�s�\�� �z��z��������r���-�ULCv�4�R�����(�X&H��1�@]̦�qۏI���6��������z!c�G[܀��^��Kո�l֋��daDn���LFB�T��Wa��k9���K��q��x��M���-��0��h�,���-}���������o���r8I+��z^�CA�)�b��ii�Q"[J�e����&���n1+3�����X��	&���Z����G�v'�^�_�i{u���}H:�%&��Zw�'�S��6c�7Gט���n�uka<�:��<�C����뿷�3����ҪՌ����0�)x�Z{�&#T�$������\;T���)6��ߒ�!d��"E�@�3��\�o]PFa�s��'_v�d�BaAI{49�	�A�%͋���
���/?:_Kc\��&E��ĲF���&'X������Wn�e���C��ӈ��c��X��
�4���ζ����}����0V;�qC�V�1U�S��]�R�x�F��"��(N���{6FnJg��D1PW��F��Q*��*Z�7h4#|��L�� V�7jS�K:&8DiJ��	gD��r�H�Zy����.l� �T��U6���t������)��Zq�偦��&4�V�#��$4�CI������6q��Hd �%���hk�C�6X�ޫ*)u�-��[ $��yld,���xd֥�j�0_{�t�ǧK�����`��K�mXx��(>y�s#�H���j?�#���x���Lq��`�ưKK_���R������Z��m�H��J���s���� \n\��1��A<`��,�z[��k3}g}[k/Z���X�H������h�(�1����w(Z�{���y�\���u��!�n�A��n�<�?Ͻ�?)ת�6VL���ϳ��͐σ����2yo.8����%MI ���K���'���ޝZ����9�:"?fV�f�)�dj,��)43��}d�v��w���Rf��qpTP�@�ht��\�J�T���u0F@�1O,g��=���q���o��{s���w0���������^�̭RfI��=��(��+@��^�&c�v1]���gw
��T��;�R��,?��qh{5v�s%}>��O���޾}E���o�����y�r
wv�"#��-=?o��Cu�?����V�p�$���̋�iW�������+�����W�27�>}�H>|�O�?�;O�v�J뛭�m�<r$�J@ڍ�%^o�d���Ӈ����=Ng�$2AӮ3`�[�G���8����_�}~���(��Ͷ�o~��޼~EW����p�R������J0غ�����J���َ���o%l�G{�@Λ!ޒd��zj.?�ڭO��f6�I"�]���6�寕�jv�pL�m�/���f��n0${l�Z�7����o���?�Y2�2xl����RA�H����wV������I���?IƵ�7�sFy��%���h�������Y��j�q-�n
�:�� �Z�H�z�ʵ4�a�)b^���Ƶ������h\l��4����"Ki�菋/��4t����n2
�>苡��'T�_ϓ%�Ǣ�P�"�J����<��Zg���8.��{Mn�;J��lB�&m6��hih�<.����}�(��j֍'}��A���G	gW�^�"k �B���l��	T¥ M���\jja����
���!�o�w'Z���+j	��T��I��z�M��r<!���X�`e<�>M�Ԙ#��d+��8<U�`�l]<s���y,-�S��Sp����������������k��k%�)��f������@[D0�܃e�V��񅘂���h��x��;�m����O����`w�g�u���ʓ�����|g����t���S h+���q?<�k�Ӛ~�k&O� `m�	��y�ߕΧY���FE"�T�K�GM{�P&u�P�ڦ*?#��6�<�cieQ_
8�RQ#ܞM]�g�b�,-���V����]�n�5�8�������O�0���@za[\w�׺Ο��#��D�v��Gľ�-;'����sk���O����s:�0'�o\^�^�S����4k*����:Qp� �%
��<ď7��HyY�l�,dn���P6ү��L��{{M���Ex�{�}M'��?��xq �߹� ���c>�Nt����"�Ɯ�T��r�)P�:@z���� ��τ2���@�cH���+}� K�_�LKF�W*����,��I�`��Ӆ>��u��c� �pI��k�)f�^B���NR�����':�+����w���~���������؛+�oU�k�T�K�3�9UR	��z��ƣu
C�f����
�C�ւ�b�����{�A*�M�nF�)9F:l��p~,X���I-խ�n}��R2.EM2�VN���^�yHuoy�%l�b�br�䒋��<-K|X�~_G�>���$�"�W��p~ζ��*���،�]�;��R]��4D��*	N�b\Xm6��'�h�|�j��Y*��zS@�s8|(��<ۊ�tӌ��/��\�D�
Ryd��l(Q�-���`�R
�J�cy��+/�L��0#B���b�*w�H��҆��4�e>��pe�� ���ll!�h0
9�E�~���9���5�:�@��f-���bt�>�&�H�(�Ř7�@�Xɉ���������A���e�i~��o}o�>��'4�X�/��r��#>Լ��I*�,!|��igN󗎦��)�!�ʜ�^�b>?�Q����ɥ\B]��8����|��O�eGj��#�9Ra�ŅqNN}iOXj��R`T�Gc �QYX��0L^�|�ρ,�C�>�_��߆�獽/��H��TX��>F��'򄞑��zdSn:KW�v���g�?#e�������U��f��3�Xcj���=H�
,�ʬg�����X� ���,^���%�i(t�I�٦P&5��P4-:�G�2�+�`֠g��Fc�ϐVZ�����OiQ��ҡ��qU�7i�%�X�7j�#cc�
eߙ"��i�~��e.�ҿ�5�e�Jq�F-�3�����YZZ��=��U��6ը�$ �-R����Y#��h���.&�&k���oZ��mP�����U���=��o~�W7o�O�W������w�@V��W�JnũH3�6�U�Y"P�`X�`K�3Ri����ۛ�fJw�x�10�h���`F���\lc�z���������H��}W�Il���+p4l���r'�Z�x��6W2���^�p���$y}��۫��H�fv�J?��3���`��>!��VߢQL��B?H)�7_����N��ng�ba.�p��[ġ����u�����~a 5�eD���J�/�B�e��'i��D �t�B/�{.��j�����k����e�ws����¶�ѡg_�=���������?�s' �3P���y�SM�'G���jӧ��j4�S�V#*F���yl>�id��=�Ց�����2�5`��JOnJ���+Đ-�y��<�)��D.�����(@x���2ΔGd}�2�	���6�y�X"��iwX%RLHŃ�(��?Ki(��,Bz��k��� +�23�����2�-����#Z����r������X��ٵ�X�P���2��h.�4��y�����7A:[�oF:��|�ۑ_��BnT%����W6�<s����~Ԕ����a C�w\��a��#� 1F`p矀!.h��Ye���`ͽtp�b���Jv�q�����ҽ�J�Y*T���n��5�?�\P�Ӝ�ԁ��5��>	" �ҁ��PM�T|�)���9�װ�l?�.��xS�{��j�� 1"��}_�(08��J�B�������S˚��i��d8UP԰�2�N����'��f��뎺����ٵ�3�����㴩}Y�9�P4�'d64\#��vk?dVZ^�s�o��� ?ovҵ�\��8@�_7-���ϦYS�K���9���(�$K�cÖ=[�u�C�&ǵ�?"5Jj
RTa1�hQT��HfT�	�T�CM�@3�Z�N�|d#�vV'1�ޱ�v���$��:ZOL-�W*�ɜ������L_���Hono��̔��S�q��۷�;����Á�؛��I��N��,=��r^)�g��H�`ե�<�\�Ա��Z�3p�����72^iD�S�cC��g���Q+�z_��a߯s�:/�-�����LDF��^�pu%-j��t�@k����1 =�JCev*l%L�dc"d�FnJ|����Qkc�M��2$=�ka�&��E�,�/JС��}�"R��՞.��k3����Wg�y���s$���n�YQ�~,�#�g��C4XA^��Ung�������������g�=	G�l��r��$�
է��#�3q�����p��~T0�Fjf#����XEc�ثD�j��~�U��"�}��� X���L����T�C��G�E��SPAm��'�j��S3�e��D[����f6#L��lv��`��ɍ�Ȇ��&�t�8<j�>��(�� �.�
��h�͞� W0cK�C)����dC�$�J�ڤʅ�����{x8�f�N��2Bާ�+"$3,�#�](R�
R^^#t:���1+'�r�� ��"@XY��Q�JT���#AV5T�=�j��bn�� �#�:���a��ۂ֮�(�D��j[�d�Hn�Ry�2+MB��_J�+&���PI&?d�u.�41i�K������eD�|MQ��GV�7*�;,��1a<�Q�Q$�o0ِkj ��lMy>`�&��� �O�w�W���c�b����]�o����[�_(�&� N���z�y�C���r~�˷�<�k#��Ð^F$����@����W�o���s��L�$N))��ܯc����UQ)��uF"�Ym%�9X ����؞��X��G�s`��N�;�¶j��j�[��/��<�0�t]�b�:�0E���D���3��I�.�p����P��h��!�s@����b$&�%�چH�R�f�?�X�1;ǳI�"��ȋױlyYI�dxQ��I��%?��V��̨&p��j��xι�q����"���oh�9>}�pO?��+}������l:��w�u�����'��e/�� �����:���,��}:��R/&��R�)P��k0����s�5-R"T`�u�)�y�8R��Z�Lv����,i}�����v�f+��#[�M�2&�،[���ͱ�BNm���Pa�/\&����]~鿛ջq�a�7̤_�w>�}����:к�mJ	IZ�O갯
��d���^�ER���K@#�>Fōcb.��x՚���>pc�
��`�V�^ނ�R�r}c�KY7�Y�vFY��hԀ��8��j32��>M�e���c�*�0{!w�^:��B&���|>������bn&�~���[�w�AEpH똕��:�c�d5`(%ճ���lAB�L"�_Y\�P������?�8Q�\>G�f��s�`��WY�Na5� Q�*���`���EP�I#r���oB�
kv�(y�͍eP����z�0<ܠ�\��B!����Q�bq<s5����I��'��E���s��T�n���]@�pԄ�����d����Ϸ��r|�7E�����L3|�-�V� �KX.���F-�oŽ���Fs2l\a.u<B��$3��~oV��cܳ����Ec_\�W[Z���l�-��֔�+�F@��O��CUdkx�aa
���S���ӡYE�Σ=XC�z�1�󃺌<v�.$�njY
��ZF9v�p�y���>���
�N�4�a�k��:�eEU���yq�/����S䛮Yt�l}dY(H8��ga��[6��������|�}Y*���0�"�s��_�
�Jڝ-��P��vnp��.qv�)M4��������k��^`%�S��v|nѧ=PB�y��gJ��%֣�jzcK���*�s��Tmz�?�>���˲�,��a�{���ب�^�\W�\�-1�����J�(�k(�0Jt�f?&�C�]�(ͲF�ߓi�B�9�ˤ̶\� �M��%y����6��)I��H
�EOh�Gb/d4z������{7��ñ��M��:��8����=}�xG,����ݻw��ի��/Vw���,){�
���ς#^�$�ok�X���Y�	OV�6;���}��wd�0aE�sf��/g%������d���YA_5�u#����k�Kt$W��� 3����7�Y, `���V��+h�MwU%����<�Y��>�`�q����{��}��~�xw���}�,z0lD���^�8X�g߳��6�������d����9&?>wo�3��֐DG�Fw��V�dXT�E�=xP�a��=�x�!F�=������<�`"��_���!]���./�o�Mو����|;�wf�'�5{f򴐕�le&�������3��{ �4�]��?�z�S<�d��g7(�1�٘ధ��3�N2b$`���f��L8�l��+*ٔyD��������zH ?��>��<�A���ES��X���{&}3���8�V] [�.�u�q2�ł2�� `�Af:}� ������`�9��7�?9M�1�p$�2r�a�CL1��F��X�J-*��\R�b��=�g�e���c����ClI��T��8�QEھs�>Y�^�_Id����D-8� ��dX>Ԕw���\>p�����q�M�"�g `"k#��6@f�
F��X�������:�~q����4�_����e�Ѯ쾮������	L���}���n����J��k���K6��TdL���a��l�`��s���ϰ�z�=E�ԧ�L��!����I�5h�ڞ>���)�)g��CN��nL��`]�a4�@0[ӵ�y��>}�cK�����u���E���u�����1�H�e^�o4+�g��O�I���� �(��\�t�/g��e���^DL��C{�d�Sj1GxV�#Ac�7�)) �_\�_�jd���cn������;�9�r�m��6���A׎y-�H�g{��A��ǴT)-<h>��E p�y�/+����a����� 8>�$�Y6���,Jc0��=����^��$�X�O�IS�c�`�g��#X�1�q�	;�Y@�g���
G��6e�N�lGK��1�e�2 S�������|~�L���8����-���Oo����&�������������J� �3���.�����cG��}�>AG��,���o�߆L�g�����`L��)o��Ck���^�3H�(��C�=C��}&�Ȉ�L2��T�5����{����>,��,#vgh�A������qXVlYr������>�����ڻ�3֕ɪl>��K/0;	���Wͤ�3�(���>�������xN{I��X�c�ſa  �%�����]�0,g��U����k��-�Ev�ٵN` �%v��L
6'����({�6�6�/L� �v�7�4�����x�$��/��t���f���Q��2> Hd�q�w;��@� �� X���B%k;=K%y>V�5Ʊ�vQ�{$33�Q�}� �h�9��r|�ϴ��W	b43m�L��/��~g-D��m�̀�0�,n`�u ��́�R�)�f�
wQ&(��0*9��53X%�hZ�W)���2��Q�q
������e'�ߖՍ�RĲ�i��\攲�4r�d�P��2��dhص�P��˃�em)�Ң��I\h�X;��f��-�ӫjڰ��h(.ݤ:}�:�8�9qN��?����k���s.\���282���{@5��ε���p�>��`;0�,͆7��ÓJ���<D��;���2�i6�K��o����� �)]��^ T�F�~d�,6}����:��ڗNIǥ)���Y`��v�L#�����Ĵ�������&��#��6�PDڄN�&�6lY����C��`���%딞�x����'���9�]��S�*����y
�'����Hd�p�!�mBh��� ��X��t�F=��ؿ��ٺjd�]�C-Β�U�~I���:;�G�����l
�|Oc����r"e�xYK�~1`�g�4���"���8�X���&����� 'p�*�udv�V���d\[��,�j��y�'���1���X�>?x�#x�ΚVެV�Y�����>S�pÐ���n>gk�-���p���L~��#�K�3�ʒ��$���X��?ҏ?����M�$A��k^ӟ�����;��I4�p��u�GR�=|.�Ѳ����r9�s{Gs��Y�f���~ֲYv����5��0~fc�T�v���/���:���_��<-[�6;�]�ΆZ>X�ˁ-���7�o?��X�����D~X���d��U�p'	�y��=��YX�#��_�T̸�O�B�3�LO	l)������+���ffv�Z&�i(�
�����Ĺq�tHp'�X�Y��v�~�6�.k�MĚE������G�@~w�=����	,0&mH����ZGX\�O��}F�>|���J��O�n�-������d��;��w����%�7�i��3P���zD��;��kُ*��t����-������齾��i�Ǐ��ֵ���Y�jJ�a>���@AO3Y 
{�xA[}���v~��P禯m���Ȋ6{E��TwD�2�eG��!$��1�008u=�9(pg�V�V��/��=4������#����������4E���IfʲX�Q����	��6
��cH3t:�;�
������-�Á��^�l��L�s���j������v��sgϟ���0Fk�tV�1js����6%ƶT9�$�:�E��׮��ߟ�-2�}�<n�2�?3�<s�F�� g��H�� h��a5H���ٝ2�㈧B�q�m�ߝ��w��n��֬�������4m�q@�6�K����� ̑��.�q�ı:XP�͍I�:�:��U�V���* ������^��ӽ���S=Y}�9�V�B�!���3{8�yi-DpF��9K��L�d'!��8?� c��@&�����sH���S�_(�ߧ��{ ���X'�Ԯ������v���VOa?�{E�۸^�F$_�V́�@˝򦎌�:�y R��*:�f��(�C��=� `�pk]3@
n'����V)lm��2�#P���s>���$��|{![`Ү����4�z �ή��u@s�&R ��9{�0ԑ��b���Y�A���uK�tZ��8\@2�����Z�<�t�\?���k�'UX���3�V�9���qb)��<�J�_�[�/�R��eeatm��K���hI>ꐭm��C��7��I �.��B�̓��v!l�܁a��h�j���lHaϝ+��3����8���RC�[�2����9��y��&���wg���`���ͤ�l��O^�.�(��g�r�B���~�q^ε�U���y^{��5/{��z� I�N�g��G>q����g��w� ��D����g�~�y9���Hp�^�g�;�<�Xw>�>32�Vwۚ����Z�_���V�2��0��h��`M��vaC���v�dR&�3�@x��a�'I��9M����^nA2sŉ�a�w���~>Tb�2��;.3�(��~M?c��p�\��+<��Le���ۼ�1�g�7��ƥF������=a�c���QB|>��#$dP��T���v�8|f������|5��d��Pܝ�{<�j$���|���_�/��ג�˹�����=�1�iy=���iH����������g��s����:(���Nx�Ͷ5�춦I��CNbl²##��,F@�f�/w������T��ڙ'�2m�hM�ƗQ,�?�d�m[��%�?27Άt������Zpѱ����X��Yw�F����.;9�JRF�\�@$>c����1u����E�Ƣ�S��bl�1o����k�ͤ����ۦ4ɀ1j?.��BL��{2 �8��fW��Ej��?���ϛ7���=���������d �ۆ<�ւX���p���1��h���2���#�u�%���|��K&���أH�,�<�_$1�����Q�=s��q��6j;�k]��/Q�>�_k�[%�#f���!�X�`A�O�aY�S'���M�H_��i8����ݰJ򗧬*����>�ufG��`�`��4
��Y�ܐS��QfeЀW),�h�8P\RH��5�����Ĕ��7�Z'����%1��Q	��Ϊ�{��e8�Y�Vp��,��Ӻ�t[�� "��c0�(Orp@������
턚�}̀F�~C$eO��Q{�8P�3������k�qNVݳ�8�6��ـ/�D5-�%�o�qsRГc��)Hn�/�����������I���� �r�WbP�� �� �
�W��$2lCM��[5�Ώ}|Ě���p"o���g$�כ�M�Ο7�j�� hג�͛5< MCF�^ k��FӺ?�6�?/�����������:A�р����B���mD���V/s�z2����jX�	WW�=K]��VM�Ŗ�X�
<������e6 �x�������z��@��B��B�а�O<H�|��č�	L��[� �vO�Z��G���}���Ϣ�U
��d]��Z���JFa�ڹ�E����z=],3󞶷��d��<[ق�)�%��ygR��~h{Rv��֪'��W�g�?4b}1��bӄ�}$"�B�	;��c��A���,��� чn������W�ִ�q%���m�y��8�~6�m�M'Q�S
Y�t��/��G����6��h�S\��3#lB�J˨�̬���q�岔P t6���<����VGM��y����-��_�H��^N�Z�!������׿%c#����_?̨����MCg��;X|y0}ѹ�{D�ݏjGpQ'�ߦ��e1�R96�l &4`����C��Y�	��,�l���e.a��!d���#X��Qa�6�/�2u��3[w�=}l��gK|1�y^2x�J�R&`���Ґ�\ٚ�Z6v��r~5���������A��v:��A��!~����i`O��>�L/�i#�l:|3�kt��d�gP7�N��}���r�]fv̍mt'�2>�F1U�U9���s\�7V��U��M��')�� �	Rt+�Z���هwu������*Xtm0��Y��5���@�,�$��|�R� 6�Qȸ�POP"�?�Ǟ��ٛ?[�g�^G����7��=,;$,^H��֎}�ݧ bޯq�Tɩ�k�C�9�v�9x��L=3�d#e�|?��X�)Y���s�p0������Ҝޗ��/�,�=���c�a��LdK��Y&7�R��)�';k�a`��7>Ypo�>�ŵ렰�
\v�v����e�� ���V&o�kw��?>�.��x{����/{ۚ�eo�7rҐk�@1��<pd�(��l�@x0�y̹H���l~��w �gd�q���ޒ"c&��L��,f��^_O�\��	o�z�g�����q�md���#�pʠ���~%�Um�%| �q��{pmA�u��9�0�������A�	� �h@��S��Y}�ͩ�������,��֩����-���$�AP�q���(E2)�e��_���}�WqϴV�Q= ������}3�Ӽ�N�$�D���S@Oӥ �������-��{jY]�u6n{L2�Y�{�g�e���������0�t�mf{�}�΃f;-�2�&�ڷ����1�l�yX��ϑ�D� ����͂x� EAV��ߟp�E�\�6�z1"�쏭ӝуd�2'7�Yf�uY����ڼ>,:@ڮgdIAa�r���m_\�.�}����l��*۾�<�D���3�`S��_��Q 7��bd�>��['fml�=�~V�e޵=�P����h��1�sP�E���E�q��Fw\����!�,����`�~?ptS7|����[������o�ŏi�v��oo>I��G����H?�O������pc*�ʉ��V��d�I�n��<���j�R�L�
��L�Bg冰���jf�vv�I���T8 4-q�8 0�3'=��� J;ke*$�9��֦E8uK�H�{�������	Tn_�-USð�A�D���7����<`��dz;/fP ʳJQ�ղ�����d�ߋh_����|4�2s� "Z�d0]fSG�X�7;�p&M�� �s�{s�1o��f0�9�BF�~_&�p
�̖����c� ���<��qNb!�(Q�?�k� K(�s���_F7(J=��k�9_����^�Y�A��>�������d؝Q��j}����p �{s�g�)�{��N���`�F�2�h6ޫ����Rݘk[��Y���[+��� P���T� S5���ܧ�9�1^��
f 8��Al��x�����S�`�)�Y[��f��k��$+in�����:�Q���L1�^ #	Щ��/!
�{�,���od)xUW�-���� �DKZ�\��m�:�1V�E�h�l�σA��_�5-�1G
��0�Z����]w^�z]�t���xm�@|8@�����~;�uv��}��v�J g����2a~���l��t��ㅀ���Xw܅�x�?Ab�̌I]�!�ln�c�.
tV�ӧ�G� �I���a_��n؜x����������1n/�a@2���m�?�;����3(ѣgDV�&ɖ��u���Ԝ!p����~�Y���9^������4��2ɂ�j�Q/~�6l���Aֹf�Z�Eֈ�Rg��։v>h�3�,��@���Y�|�؍��_����ž�#��d�H3�ȸm_���Lo(Z�帐k,(�(ݱL���胀 �[��V/�hDf&�QH�>��+���=�����;,Ve��J�qш ���9�����ϢM5�����1J ���/�geA=���/����q��H��oه���{�����W��n������m��5n����(�7�0"��fa2g���&��rd�J�%��i
�
�Cm3!#%���7��!<��� ������q�,�Ro��Ih��ӌ?�'GPw�B㐅�M!��v#�3eF,s C����A:�[F#���A�r���t/ˉ1VS���X����	��^����\&����Ӱ����j��:ۡ�����ցn5v�83)hY��c%���#9�ZL4nF9j{�as��o���7�`T�B�Bc��@���X ���:?��>.�>$#�)g�)N�hb�^,�{�XoWI�(�c߫fFp2���E|[� Y��l��8B�a ���>�:7HP����دX|\`��Ӽ�̙���Rϒn)+�hUD��<E��˸�`/:]�ra2���z �ؠ��"3b�)�|<��: �N��Ui�	c�3��Sf�F�b����]5n��#�F�� �-[;淉ђ3`���Ƴ�v�	��2�����I�O�g�Y�n{`C����d�2}�!�||^�iئ���z���0���X����Or]�w��t/�;`�"p�,���e7$EP��j�s��-��?�CH:��쳣f��� �}���<�6�r�D��Sm�ϙ��ImO!��� ��3��5%��K��5>��M�wI��-�_2�Oҙl������Tw��8 �d��3�\�,)jҨ��3��M��[i;�ǤϞ�8?_?��]:��$��Ɛ��F�i���ll�56�*dzE\����[e'bEsc]�t��,ɝ�7U,����9�`at�[�8@������e-�B+�I�"
b
%Q�۰��*o�ߐ��^�@@��׍ �g���/�M�|� �3�?׹H���/��X���ﲃ̵�Sd-%�\=Z���=2 ���#g��׌�{9��W�����P~���j��Q�k{�!9upU5�\�?�:��9�n� �,n;O�wX�����ؒF=��(��|�A��p�/�Pn�,�p=y�@�bJOR� [�iJ����g���y��J���MA��g�1v�T����H_31a��P2$��5���:�MJe���ʦu��ݳN��T@iY^��w�:H����?f��5P��fi���D���.��1 ��s-�|��氈�&���X~���l����b�&�+8���q�.A��t�8˟�B0W��陟I)ݖ��8�q.�2`�]��b"KF� ����I�W���&�~!#)�h��\��vF^�YV�ۭ"�8c�#��c�%�fA��{��ype�	����dޭ��{�ĩĢ����zN-p�D�1�b����cM�bOς�$�n�ϒ����}j������d�t́����)�~����9�D�%5Ӥ+�4����=�y��n`u8a傰,������!Δ�Fv�Á�݄�A��+��܍�rM�ϱ�w�{_��t��������X��xV��a��5�7;s��]k�2KR�%��TOsv��1R�f��(�/L���\+�tC*��Z�׶�X���x+wJ`���_��gn�1���5�h�����Ɠ�JA�`1�2{���e��������<���|>{'��y}�4l�@&A�5`�&ʹ���o��1�+k[�3?N��p�vr��=�ޣ���Y4��<��y�͇�b̩�����r���߇������d9�8��V2�C͍�!m�oE:��E�5��+��i�7���c�33���a�e�)�|{!�N`ڍ��|�Ϛ&���k�G�ˬSΚO4ZX��C���#ö>���
E`�'I��}�f`�1V�Y�9�S��E�A�QF�-�B��]dݳ�y'&M�f{w������)���$!u�NmHa9! �t6\�=��ᫍ����.#��p���<���H��ߪ?OU���o���c��1z�#[h��پ�fK��l �,������+��G��g0��-���\l��dǻW���b�D��_ $���Q]�,(yy�#DV'L{���q_�$06�˓����A� ��u�Z�wϽn[�0��R��]��>H���?0{����	����v!�0 P�ޯ������^%	csO�P)��
j�
�}�B4fZ���>?�.����"�?���v;��`i�P/fx�|��l�Ҽ>�1�b8��=�4���L5oPa�8��{ty�<�������5����S �4-�=6��u���Թ8��P�+�h-Km��6o����ȳ� ���2���#hM�[67�u����{�ӡ�j,䗕as�sڼdG2"�#Ic�A��桏�����P.@��@��CAe_�a�Z�Ns��]��f~�]D��\+�rGS��|��`��N%��c�9N!��$�m��ps4�h$�V���>ajp��J>Nd%�s�dv-����2� ��S'�{	r�2����O;�wJ��l�٣����&i4|ks2��k�Q���|�=��e��:��/@P��k|�U.y��)	����Wx/����T
��n�&n�P�L�+���s���Y�.�Ȥ��6hX���[f� ���'�"���̊��.3��- C��̌��lHQ���y
vNz���+�5�7m��O+c�?�0<��H�_�x[Z[Ԉ(���Ե0�X���}*�A�� d�.DǓ��t��:�.�dTcC�<:4A��d!huOR�t�ۂ�m�I����s<N���3��H.����;�ct L[:F95d3FVA�?4�mԵ}I���L]`���e_�:i�����)e����,��O�)�˙YI1��]�P9.��ͬ��������j��MX&fʳ��y&�I�Z����N$����Ug�t~���7�� �� �h2T�oG7�Yz���a�,������؍z���رo�@������$�`�^rY�YZ�O�q�N������2]^���c��C�|3e$qzxZb�fP%K�@�$N�}�#ٹ\���fޫ��f�l )�P��o�ĉ#��\z��@Į�{I4� |Jd��u��}{?¡�%��f��v%�l���7��i#�w�� �5P(0��>�:�f"�Y2������1�sP� �`�]�H&U�g��؃ �}�i�H��۞8m�����|sҋ�%�1��e;�u���"�^$��}q�Z�>�;Oy�R'��l�C��8�hCҕ� 3�l�`��ݤ�݁�u��jo`�Uq�� �����yl��<����ŐAI�� �T��q*� �[��k��; �Bѻ���C�q���j�efM��*�*�$ںm�O?2�H� �`��T(5�z?l7����r�q�uW<A��;�9�$��D�(+h���� �wq��U�~܃��
�fɠ;�C��:�f+�?�����k�q�u�����KV#��fsn��݂�-�_�*gC��ף+LL�u�/���;�C6���0r�6�@8R=��k��<�hsV�b�݊���RfZ��A����i��=+����T��@7�s9e㷴����T�K���{M ֆ:����54h�`EVN˰�%'�r\�}Ee�gH��J?s�P%�o��ߩ�4" �c�X	{�d������_+�3�k7w�^�5���m�j�QeTv�5Dۯ�9�돡}�Yu]�F#�v"��5�`���_eQb���;�/���k���@�5�FV��ư_NH0�|lh������a�;�*�����'9~'�b�
���L��A	��E(��iĀ ����ut��D�@�oZ�g�Y�tߧ��	��b<q��a�Х����&��X��(����v.{�{'�S�Q��<�㡝]G�Gz]{X;�r�7g���F��<�����l��}填��[��E�L��H���~�(7"O��g��o��˵�_�fNC���oC��Y��<>�������	`�z�jI:����z�w;�"���=Q�%Fĺ8Bg���Z<>��A��tJ�b<|ܿ���V�T���!9S+��LR���N�1���ҩ���X=j)�M��E�ް�<��
w$m!p�}��2eH�����4Of�j�٭P�S��Y�\��/$Z����0�<���fV�wӄ��_��]�o��$ݜf���9Z�ɉ08����G��-y�ݘ�cH+l��Q0��(|�÷��1��=��������-��u[�2��qtx+j�2bP�JL�\�RcѠO�����fy�h3����ʂ\���o??���%������k'j�,Y�)�� p�N)2'��|��
Ճ�%�f[`lY��n�53�F^_��O���:�(�������Y��V<cP'۠��g4��M'��r�mc.��2���0����SAV�K���w?Qo�Z�Q���-�-#�(WDP_dAU��!��,${���o�٫�3����/7�8 x�
����gMx��KTvd�s��| 6[��&�m�2aFlZ�È��FDyC���l��%56�#�P�
6�t6"9I� Z<L� R���ϴ�����,Ka�@���p����p���/�Œ��آ�]�����u�si4y0�h����3�[w?�σk����v����ȍh3n������75P��;� 2�	l�Z�sj�7f�l�X�ۺ��C��M�c�V*ز"��`��@��e��s��7���Pn��� �H���j51d1��$w�������] Qpݬ����,��֊̢Y`�aǗؙh%�(����je�t��e�FP���&cN����J��A��V6���n�%�z'��J0��,b�ʵ#�_���m��l;�� ��QC���"�m�ڂ��}���o�>�U+�g�z[���fj�4�|���Gcɐ᧐9�IHL�d�����!�L��v��#A$_ٳg�gx8�D�Ğ�ւ�~:��,���H i+��X���{vxXc�W�2�M�T�jX����^�U]#�t6���cC��~�{W�~��`��H[�kq[hG�Z��82�0�&	"R�������S|^q����8qX2�b�&AvHF���}%tGB#<u!�vu�m2�YF6�]HIG<���E��/�v�cR��U��ԟJʁm.O:�������;���Oip��c��p�(P����CA��<0�{���e�XoĚ%�/l+_�J�S˵2���H㤭F��F$SF)�nN���Y�#'�����R����f��z��A�s�lHmX[a�³?��i*���
�� ��@�hJ�Sؗ`��d���W�-���*��L�Bd�w1�9�,�kР�[����.E���C�V���Ԃ[��m6����dg�����%ż婭7Z8�?�c�Q��}�5~[F���,ey��Νs��~{M�%}~,鱭I���fq�fK�������A ż��c	Ш�%r8n�لCu����`��y/[=���EY�Uu>��rIjn��-y��P.����A�k��g��K��{ٷ=֝��s�:/"f��mԌ�i��w8�l�i'۝pQ�77O���` ։���y�)��,` �Yu�/�wR����$\��7w��b.��vW���)+���@�����^_٨b���#{t�'�pm((s�ǘ��|~b���ܢɊ~n�y�m?𲫓�u�L.7ּ�.�j���F�2$���-I^�w�n��N� �s�l�fl�GÁ�%,����Õ1v�����ϫ���ϻ_�l��o�8��#-�׆���ٌuYY���+Y�$�/&` ���^i���Z6a=Q��~ν�UBpF�ۋ)w��9
[�7d�17�q�_�"@ݭ:�dÚ��ԃ�vy�R"��u��'��!�Й`��؀H�!�*���ױ{S���$���]Y�ȩ�4�	��f����O��F�@�3-{�hתg����vb���^�S��I%�G-��ܯYc�\���I�//�p\7�͵ZA�s���Q��b�NID��5��y���YX��Ȧ�V&�	)rʨW�yde�=I�����-H�����\�w��3����,��l�n�����{���M1�l맆�lh-p�|n�䥉�R�8j��g2���u�^�����H���1<���k�}`��Z/�_{A��d�u\`����d�˙��6�����Ć��FS,���-���̔Xg6B'�c-pAp1g��'t��3��I��'c�P �44�2����uT
�?	���25�����E�R�N��,��h(ceْ[c��,�N�����m��u|�� M�J����h�����M`c<�������x=�����}o�
�b���QF��:��h
 F�i�����#+`�9ǹ��W�/ms��(���8n�(���nF��2[��r��X���zs��c��E]	uߺW]cy`2>z	��3O-t���$����E��
f�~nI�b�ͺ�����	��&���B��`	i����-xH�!�T�S@��SmQ�Q2��_j��٤`�z�`#��pS������At ����@�w��j1l�,j�����c��FM�k������>���j�2�)�Q�-"d�>����@��1dvfk���$aYu��R�긌1;t��&�t�y��!9�W���/@F�5��()��?7����S4ZZj�q��{!�R���*ӳ������O�A,@M� k� �h�=�M���tU��FG��7��ݱ�&���Z�@|�5��O����e���,l��Mk�b �,a�H��� ������o9�T#V8lNk<d�GMm�
�%����@��:��l��t��������l�,
"�`{+S]��#�k&�gu�侲���_q�ѡ�KTy���_�����xp�]3��Qy���5Z��@�$43B�I�,��� �.�i&�� �$�� ���T�A�ƾf	����l.LZZ��m�ӹ�i�ed|m�X�,�%u�h�l�w6���s���,�e��t�'a���|�+��Uh�O��	�'�PO���z��> ���՜��X���p�K�L��ΥK�,��7H������_(��+���0u$�Ϙ�?�:�Raoa	�Ov���j�2�Q~1�٭X���]�ި�|���v}S�"�o����W6�S��M��$�6Cu�<�K�ȏ������=�IY�J5UAL��0����"��zg���~���r�    IEND�B`�PK   �n�Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   �n�Xj	hY� {� /   images/a580090c-3dfd-4391-b47e-11bb84c3f632.png\|\�W�~�UڪмVq (D�����L��" Ђ2�2Dd��W���!2d��ȪJ���"��d�a�B��'$������7��s����>��w�Wc�M?����m�?�k��m(���[��"���?��������'�;2���=O�����_��[S�r�>��{������7���#.  @������9OGo��1�8�n���/��F:B
v��q=�J��O.m�1>vմ&kז��s{�5<M����?	�եy_kj�r�A`зUM���R~~{�/ϻ��ｧ_�����,Ͽ���U��e�X^�P4!�jWb�bN�T��x��j�eǬ���oq�!�����N��Pa���4�FͰ�*V��҅˅��S�[�Z�ԓ���>k^�dL���C�S���u�)a�\�{g���G1���J:�ލ�H5-��9�K��v��ELk�����~�<,fD�ݧ��ֱ�6��[.�b_I�y�3�:@E��.�?������͜�q���j��c�A�_ϔ_�OT���_�S#��!�ry�W��'ݦ&�:4}'����\���{+��4S�N���$��І�>��5��R�ю�̚�Uv �XdXd�;W-+�#�]���}oC@*:��>$�DW�]044���U�.h�GX��^1v����ސcvt���M�\=螯a�Z��4�K'���G��)��ø	9"��(�g"D���tX�j�:티7�/�����E�{�7�д�뽨�:�9V�����P�\�����5П�u��qj�_c'Kh�Q��y�a_��{�6J��1t�xgۆ��y�/������cM�V�Mp��O��6NQ����jiȜ��v�o��k�_4��K�r���O���C}��l��MȖZ����ا)/�gn�^5x�rL_8�T��
y�uW��<����פּҚ.�8p@l��
��ۋ5X�����5#Xv�9��3�h�Q�>���Qz�����4!��ݩ�c�����u���1B�9E����{��_2Xt7v���yz���02�s)aN'�q��s�����OԜ�Fخ���W@��ʎΰ�_>��b���3��宒 �|V�)�s�޶%Qf�}��HS���I��.��F%;/C:t��j�R
<���Dr�x`c�b���]��=�"��:7F8}�l�o|�2o��<�{B?����0G�Sc��[�g!�Y�Ú4���k����+�����^��A���T�0�?�5C����ƙ.�����4������
ύ/����i������ݻ{4��Tc�1<�8%j��7��I��6�v�QMg��}�b��h4qu�O�6��������x�CN+[�0��=�Yv�zִ�mG�r���o�G��(������y������զ�G�-敱-H�.M�[u��W�CY��D��\�"7�5��[}�p����K �tf�Lu'/�.{�F�Pyne�677��w�p�)g�����f1����R?^����ƚξ����nV����=׸��D��ܠ̋���]%��ޓ5��ν#aa��I�n���X9n��f���2����T����R��Hk&7m�Z�Ew��J��5m�#�h#�)�;d�ax{IV�{#�:��}�9�ŝ������Xqn���_z���7�Y�^�t�<���ۆ�c݁C�� >���	�����9'Db��OV$"zҨ��_==�b�]�m�ӑ���y�Y�T��a��G�ku�ۙ�q)+D=�!������]E��#}��ѷ�fj?RK����g1�/Z�lv�Čz;������qM�Vu� ��̋t�Ř/^��|���\���_nD�E�Բ�S���2�&H��%L��/؄�{��]�˧���f�*�G�O�i��8<r��'���6����jV� Yv��'��ڸ~��Z�
y�L�;�9==�\�9֒�t�����3i+5Y�{����5�G�8r��|�3'�u|�(Ed���������-O����q�������X�����l ��q�Ȉ[o����O}1Id=�A�e��GeW�lkj����d�NY��hx;-j�5fci��E裻`����}��Lp�(|Zܡ<&�~H���k���}��V߿�jLo��OL�py^;1Ɩ�-�Zd�A𬄐��,5��0�l$���5����������c�����g@l%������4�g�2m���Q��(��Sv��]��� ��%U�o��(fI#��2�sD������4�W�IUo�\vK\�c��6/���������wT�!�Izz�Y���U	9�&�^}
8\J������Ӛ1B�bѧG���Qf�t��[^�e.� Ԟ �j�$pۀWjq�\�w�tY13XOv�`vqy�[�<��|�w�f�]N�V�Ј�&��>���\�6�5~^L����R�s����.�y��'��xgxx��P���a߲̅?��>l��L�}mJ����^L͓����X��L&nJLI){�7F�إ�m89��,>gl����Y��vh�_^�ё�$� ���3��T�΄�ۄF�w.�p�4�N1��F���Ba���XgH	�X�x�7?�ONI	7�uԣ�r.�D�X�c\����{`�ޜ50�ۆ":cѝZ1u˧�`�ς$��*�E�J<_, T۷Zl];Kss=���0~݅U.i��$�(JY��_��{�`lԝ�0�)"��t�5D�f������5�����	�듆�%fQ�C"ٞj%Z�~?�âx&n�	N4�M� ���y�-"�e��W5(����X���*ͯ_�����Q�w��oB�E����~�G���~��-�E��5k�~��u���ٗ�Q�e`����>f��Aa63؍GhkG�=I�HvȚa����u�[m�/�Z�����d���Y3�Q�h\��'�b:�\;;�}ݓ��{�cEf�a4���O���7ɴ�6���>.ji���,^�`����&��aA�|��"�|�+�>�?
�iU�T��i��ʡS���Y�K����#��y���ƙ�2IV�	���nZӐT�OY
OnfG\�1}�gy]E�������c�M����Z~�w"..��+\��2�!�
�4���_�4g�̍iu�p��N����Ne ۺ����Q�|�^�p������0��<,��X#z�=�!]e���Gt��V5 ��5����$o"pQ0=�K�E�-7�v=�bo Rm�b����qx��b�ռ��x���k��3i��w�i��S�\=�ke��N#D�u-������9	$�x_Y��-����kg۰���k�t��g�h�bCY	����[�/��4$:3P-.�-*��ӝv9s%Vl���=���L��ɒº�Ul [|����@R6b !��^_ꭲc��s��ZPg�ߠP]�׎w��g�!�ڝ/�
,�����ߟ�����L��	�ĖF��`B��Qme���2��:^����}õoFFF���Q�쫮�x�]G���/�F�]�6�c�3��g_}�w��j�y6�t��
z����#�J��\SE�8��in�vHLأq�	k��aE
8d\TiOp �&\J�8z���+B1HJT�R�j>��y�P�=�(G+�O���s+z~�� ���1m1T`�`����cÞ�Z�i�''�����p����]8R�Ȕ����j��c7@�waF1+o��1��e� e�7فX0@���F����/�2��[�H��6cdT�儾��k)������� V�1&����(�Yh���X�g�իWC���rQ<3r�s���l"8��St�,����H�XY1/6���̱�8;]��)͢��w�eoŠ���4��8m�6P�m�K��C,���`Q��2����߿?�,��/����,1�5]�Ɋ�B2�p�s�bVL��>��d�FeǄQna���3���c&�5����h7��o�HH���gk`b;�5�h�Υ����}Ց�Y�T��5��G���ᘏ��M�sEﰬ�{�)͘�F�'u�
���B�$Yc��í���#c�Baǔ���G@��u���8A��]O����3�)?(kh����?;cJ䫏c�<�+MI�z��P O��W�C�x��O��a����[��`���z���1"�wʇy%$#c��˻#~��!g���f]A�~���5��t�Ҷ�hB�T(�����~��Ϛ��)Ѭ>�%��q���Pv @�ʫl��5 '��n2B?��e���c���~
���+������PU��2��
��%!>��!���e�~H�dz�"���ȏ��x3m�*���s�glbll��~)���%S�1�j,��}�Ҳ �>s/�ϔ��e����sԔ/-?'�`!&URl�0���


��X:�%c�L:��� �䜓�ǀ�.&a��	=]���1����>FĜ����G���c�8Z���@�b���(�����Ϯ��X�e��.}v����wy�"��Ž0g��A���a0X��9𦓳s��x��h�?���1�R��5�����M�	���@I�n���욕�3��ҕ+��I���\՘�A�����|�q�Weee�a_u�>S��펈�R������
��A�pr��Ih+	��1��@VU:(�rK1#�W��㚥
�ZvU������݌��̬U,���
�2�XHC����������q��q�2���G4*���L���r�E�����؜"/dOILHH��ԁ���'�[}��(��-�b��J��65#�,��涍��^�.{�����e�쌱a!v���k�iMNtU_@#VFQ�=0 e��h�	
U�Z�z�%@���y�d��Օ�˻����@���o��~���yN`�N�惭A���@+��QGk؂����QV��1�[!';�Lɮy��lJ�����w�Bбt�TD.#��			����j��LWŹ7�'ˬ�FSSS'W��s��~���w7�N�*����b�G���Ì���dS
�5����n?Ћ��)}U�˩z��<0��+QQ��n�e[Ft��u����59�T�2N�r�n?�F�߸�<��)V���)��3�0Fw�)�����3jShR���9 �R^.0'�n�T����XSlZV��`.�n޼�\�&[�B��w��#O+���{�6EE1�@�ǜ��!�� (�]X��N"'��� �խ2��1sqџ�t�&΀�v'R֚HS睜��	����dn0Q�@�0��	&�k{�0��P��18%)�HoF�1�ܯo��v���J폾�U���aH1ê�2c��w o`�g�ΝChsϥ�҅A�*�z{{�_�F�a�p��>�>�����	���a�D	������b<�'�:��q]�FUm@��jI����a�e��=L���Z���oU�y@op�8���%�� ҍ�7�t�4j���,�Y�������� Ȗ�s� ��I[�)֗�T��v�)c�#�+�LL���Lk��Y�ő�gnE�Xuk92��VHx�U¸&���P�r�Y����1����{)��d�~�������?�hk�	�L�L����j�Uz8��@}B�Y�1w��ȥ�tF��3X�x�^���_�b�)�.%�Q�=(���@+Pٶ1\��)֢^���Z^]]�&�Nh�,�
É�)#����30 ���<�=�%�Ş)��.�vE�2�A-q���v=��F��_�X��O 8Hhc�	�h۹rA(��%�K>`���B�"n��V�R���uo��$��r��.��	l+�[�ӈ���](��Y334j�{'�ѷcU�����9t'�g��)+O%����C���n�iM1iS�»"1�k�@/W[^�\�9�#K\�[�j	��*O�P{J{�1y@\�.���iW�6'&p���&)��Q�a\pF�����p?�B��	1*���MT�LÃX�㭮�����'��m'x�����r��L����|��x��`�r<�ff�j�|�e��~��]TYhQ�ueD	�]Z+2gO�\����f_!�a�.�/=�X�=�D��ZH-pl���1����!����]������3��:��o�''�- �F;y�S��B'��w��P����i�(�T�ǉ�A\����hC�!���Zs�õ����6
3h��h�w��6��q�)�b���eݍ�SJ�N.�x��k�n����{Rtv�;�%��Fݞ�aDrn�*O��)�@,I���^֌��֭KOy�/��_��r�bQɖǒ$g�w>�f�$.!�Zm�C�Z�cם��<>jV�5����B0��s� f|��V�ml���n�)��b�����c��RB�b�g�b؍�%��u�?�d2'���|)��#;n�ø/a��&�V?���p� V�b�Z=�e�<v	GF4a�ޫԀةd��o<�'�a��>�	�/����4 U��b�i�!ȉ�X�yQ)s�~ph(�P�)��7(�St��.���~�rr�x��1��E���6W�1n�����W^��X��������wz2��t&��:��7`V�3)�:?|��ow���@��@�a�_��%&�2�s��sZ�P�v"�=��O	�1��=1b$m���f�R��-�]�������#Y�����?�U�1��e}Έ�**Z|Bh�ĳ�!�%De����OO���`�����m�����҅�<�G^�S'oG)}z�S���6&.����qY�"��F�h��V�0]C#
"�!l��}��Vk4�Bv�O��R�1��"t��ޔ������ލ���Kk�tK�.Q�csL��`�P�mb��/��5`�!a���_���H~�Ә8����BA瀎��S�6��a�I^�,��y�7P��=q�iJ:5���_t�P�IK&ݽs��,L��s���h3�p��hRL�>(�"ǧ|���󱕙�}��2���Xůc&d&m���6�;�x�?�8�Y*�K��ANk�vu"����p��-bóf� ��Xb��Z�~?�Fr�E"e�
P�X�� ��s�@oŐ��	䜽�k�+��m,%�Aap<�JhhU.�L�]?��g����= R��867��)ڝ��uւ�Yݔ��+'������+`�'��4�2~ɒ�r^��Ӽ�h�Gp�Q�Vȓ&�"߱g�M&����y��L����T@�<�l+�lz�5�֘������;�
�DUA���}�+W�J�L�gaOqj��{����.o��)�����z1%��6`�DOMr B��_-0w[�G`��,�B�$(�u~��UH���ڊ�_6cK��cKm������H$[=�r��7�]��K0[ �1;�ы#��N ���¶%E�\�P�)��G�0j�S��4��'7���a�T5�@	�	b{�ut��s��4C;�L;�aZ3�7ȏ�ΣIܙ̴<����������vcU�L���޻w�������UPOGau��t�lE��"��X�~��s7}	:~4����l^��1�t�¹��|Z%�H�e�32���RY�^$̲��<l{!��e1s&�R�ﴓW"��a%���W�/���о�c+CԁL��fyz;b�2��S�&�T����u�&�Emg�M�SZ�����M6�g��+�wAhmQ��]�*y@�����^���w�''&��Q�*����[`dk4���/�^��8���`uqq�X���0����	�Uh�)�A��V鄋<�ƙ�+�QS��>x�i�C;�E�v�B�	�| մ��`��?��Y,ӡ�BL�=�(��Y�N�f�ُ��,����Ӂ��^V��\ysa�`�Y�Re�>z~}�܃�<����י�|���?�O�xr6�o���\�=��p����+w����'^�fL��U�R3`}h��+ &�[�'X��7EVHa5T��RGt����(�,��67��'(�X�m/��B�_�ڇ�7��y���T����搷�u�G�d��f'$,�Ǚ��*m[tA��ӄ��qPEK�{��}.�R��%^E�Ur��"����XG".��ػ���y�ѥ�rD:F�sa�o������H�ǧV!��������\���w[I�e���~��qʌ���.���x���¥�[�qq���nu��j��@N�O7�M�\�&���/F��8#�,�>=�������V��l5���������y�P��7���-9ڢ)eh�����8��V���N��l�_��J��S8�[��@f4��z��-�Jy��%���s����G��SӤ�?[ٝw��c4�VH���{�ښ;n����!�����D��ziM�� �~���)4T��.���:�Q���Q9?0���4��3m���W�(��C�jI>i�O������y�7�b��Ng�Fw7�g�P���5u)K�� ȋo������0�D\��á�Lqv���on�	p��iM��okю�9�_{�Z���1�ihF�}W��!����ip��������:!�6�րE�5���l�r��<��k�<��������G���S��W/�M\r�m�}|N���e<|��?Ϙ�����~�Ӗ-[�N5$(�|V#�s�6#��}B�O�Gw�]�+N���6��!�t���,-n���a��۞�^�Qv<��I�n'���@�����~�R�
���`�`���k댋k)�����.��\����b{C���̀b��ldN�h�S��O��^X_EV;���J�K?K.����t,D�BB���g���;�v��\ =J-ٗY�C"�ԧ_w e)c�gQ�Ʃ�"n���yT�sz�DwS��Fo�x��:�a�f��ݬ�EK��� ]MM�f겴R��P'���l�v�B]0�.ln0\�W�����I��- ��{���T#@Ġ�?R!ݹ1�e�a�j1�L�5���ˠg.VlRU)D���O)g��p}=�&9����γn���o@;"�+dd_�]<��)�F��a��wGǁg(d��0�>�lT��.E��ڊ�ӇV*��a�S�Z9������l�@`l���N����m��y=�����X��Y`��H	��.NNNβ����^V��Y?YZD~II��0�Pk�˸Z�m��>*'u�y�GĤ�cÎ����uh��zl_e1a��(���d����aaܽ�"K,��ܳ�`1m�텳Iy�r�`�����s�"�7z�w�����yŻ&�;��~a�@�o�ϭ����ӖEWD��0�Ia!n�����L�.��=��e1��6�.A�c�s�)=ߺ��N��d�8���-����s��֨܉��!o�58F��+p�Y�L������6t:}���¢��Lo���gv�5�v`v���6��e?/$��Q��ŝ��R4��܎�H��aF��^�q��8�f��"껩��X�D���H��f75�1[{�7�a>�qOꚨ�rƻJ9:�Æ�ER��6��>c�*�ҍSD�ӛ��p��Q߉��4��k��Y �r}*)#cl^�x�����:r��>���t�5B@���rڼe�To�d��^��)ʑ�Z[[k1 �>��+���:V��ˣ�����mo=Q�?a��Q'�@Mtw���Q��g�[P}4�TSS�9ܳ���D�E���lhX�JU]^U�J�2�=��(f7ЅC��sy{��^;�]��m8g��ȇ	�85-� f�e|gt��M�x�ʎ�/��Y�u��2D�7Iƶ��r�R�C\���a��2������:�=��*�� ��^8F��6������n���z�È���#���a%̒�����]�%i�������Sja0Tj�As����!����H|$_+��9�����mj agm��cE��aT�/���_�rL�`T����x��b����S�2�u�g��Mf�f���|��ho�+Z�ٕ�A]�E�[*����Y��}��ĝ��� [�6��8[����}�z��'Ɂ�+P��;4n��|���]k0���=w����|�o��|S��=z�>�,���X��NnF���'�jYɆ����9\���5N��/ُʡ�[m;pU����٩�rcY� ��ψ�N�c����1�E}Y��� L�V7�8�����z����<�BR�#�(;�z���Jz�ꏩe?��ZY)�4W��1{{{ǒ5ʤ%�I�T4.��
r`xN+[���O�e��(5.ϸ�W^���xCV�Z�V\3�J�do:���A�a�߲���]���gQ�������#S��6~����'.�X���/{����{�&�-?L�f[�,4gP��kGa��{���O�e��D2zO������VG3�
!�0o	Ы���}ȧ�x�qKkkNB�`�^/
�4hy6V�De޹a^��E}Փ�#+�0����Q6wf��h�xG�T�cj�^I:�!�i�ٗn!�V�.3 �]7��������n�?p��π����ɵ����%ѣ#k' `���{�m��Z)�A�F�ssn B�'�(�k(T`�ne�":k�W�D����Ь��������6Y��������8�|s��v��f�^r��n�X�����|#L�O\���nk��֔����{LU�N^�ߙx�f;^'��1d�a��PC�M����ϩ�V����k�����B|���G��o�v����(]~tXR��,����Y�����X�K�F�sYZ���;+�G����D���)D��0�L*h6�)-�d�Nג,���a���7�`�5����'��@"�ގ�txUMy��0���Վ`@�m���YT�7�o��ׅ�!�b�(��2(�U�Jے���"T%�����@�HNށ�.}��X7Q�;��8���K�\r�Q���?�6��m6B4������Ғ��ߌ����8z�r�pdt#��p?��3 4%�(�W����V,ڌE/�me��2ȫ�gYdq@V6;Z�,YM�'D��{�u'�d|�s����wl�G���N�U}�g�,Y�0��aa�v�m�3���n%�C��Z�?�&�5*��։�:�
[���n\E9�Q�ު��9u�������U�C�0#j�S�߀�>g0����O|�#����R�H�"e�p�u��^�.��v�Ȣ�?�2����y._���F~�[�A|"rAd5?��A[p��=��f~
������
,> C�T�t�ɸ;p q�³|V�;\���Ӣ����v�z	D*�(���Mr`��p���i�cyyyC��C��2�Q7����O\#Z� �vuj���H�*��,BW]��mk�r�5/޺S1� �A;�� sS0B���̚k��|�B.P*�=�ʿ�Ǣ�Ns���*�1��ۭ��.���!�N-65���ٛ�Ź�/]��bcR��_��7��:�d2��2>��Bpad�y�0nVҩv[�,o~�v���|�[�v������NT&iӯ��� ��Ɂ������VFC��5ۈ����A@���g��LՐ�}�oÌ�]��?�w����h���,�s;�{���M�t7��4D,�[�7�w�ӡmD������+�$�76.�.�s��� �V5� ��((�����!>Z�MO�|��)G�h�P+Y�-�M݋��7+I{�\
`|	},���$��ݚ�A,z�U~p=�ċrs=���F�C(��fi[sst���M绕M�2�L���YZw�Z�������>kn.r�<�[��'{��i:X���w�1��VFF����b~g���������r��"�[ J����-�/�*�\i8��"v���	4�)���}���cj׏�r1��h6V�Li���?X������QV~N�(��`(�u��G�b�J��w�a�S�Mt1o�Mq$�6��nU�h�[d�8p�G��m���
Uԝ��SHF��:�j������+��$"�<BB��o@�x/>`p֙n���ӟe�+���?�����}�ƍG���Y��D64?�PG0W�p����4�~B?A��0ɂ�E�:9i�B�Z6;��>"�[�����`�F�^��������0�ӟ��0�)���X)�����I�IE����j���%�$���d��:����`��q��'��(^�Z��C�MF�\��n{����Q���s�x ը�w����W�K2�d���S���[�`�n��ޡ�u���U���9�ڰ��G��`��p4%%����3�%$�ks_��L)��W��aC���`����M�J�h�b����m�Fw1�g7v�!���W��n���/�VR_�Z'L��X�6b �,��S�-~"S��5q�d
�=cڬ"Q�{m��yK���n�+�8^f�љ�9���k�v}���cL�9��LzsP�n�*{Gdir SE˳g�"Ha�)?1=;�N�ڎ/��)RctU�Lvf�M*���'TW�-l[u�M�
@���m����k� �KB��?�Ȱ��b��y�qG��g|"0���A�|���ٌ������exAz���Wܙs�DZ���jvv��Ґ��l�b�(r:���L}����J��к�2�Q����@�:9R���%Q���9ziMB�瓠�X>F9pV��/בK�wx��²����"�I()X�j<�B;5�����3�AX�Z�ؔx �
A��R�N	X"�l+()�_Xtg?�dK��n�HVI���<�Li��g%U��B]"����oG2�Hd�Z!ᑓ��F�F�ğcI�V-p�f �q0]��Phk�+���1衫y���'�J��R�K��Е�z���%5�17�lYMfu�>��=��� '����#z:����>joo�|R7� Z�4j��L�������ې9	�"ͫl�(~��ב���xW:��="7�v���� zG0w��f�s�n��i׳���+軞��~t�XD���677�A�&�� n�w�]�U�րlm�-J�H�2A�H�v
Ķ�ӆS����-k\�_���h**��A�X�;��8�v	�DN��	f�ѻ���9h귾�����DeLA:���?������UĻ$gd(� ��������`2���J�����HHX��]�`W��#���K&Z�j|P�wF���8���g;^e)�j�򳅓�
��I,t1��!f�mYIR\�*�&?�9��jB[;�c\F1=\璞L��f����k��Ү�CFSe�U��It��k�[,�hr����Ͷ��&�vve�P��L?c/4�-TRP.���ei��]��PV���M�-#�G�7����|7��]�A�� ���+%��Q3���D�^���^U\�Ē�M[g��'R�j{�9�|״(N�C�s�K������d�����h<ɉC�i�]��)8���
����wc=mDC�)E����{���Y_6��ɰ��j^�t�	�@Tߞ�W�X�6"�4�V���N��t�!_�A���P��x�L�6��P�oَ(Zd�G���(:R��jw�x��IO_�h���;0݊4|���r`����b-�b���$�/ͿC%��F�B�4]�T�b�`�{k29=��Sg׭��+��-�l��ߐ��~\1��m��{>G5����
��k��6�\�{+�o�:YS��O�1�$%{W4L-�^#:m�OP���ߩ��vE��0�����P�N��은.��E��T,U���qx��.���r�Lp)�lSDj>������M�8�a)3z��h�_Aal�W=N��m.�C�+�T���3�G�@ؑ���������S=T�c��Lp�J}]2F� lD�$W���$��9���=�����V..aئ�<��؈?��^�Zs��C�$��;�6��Oh��R���_e���Z����!�NAall����ps��'�V�j�Y�]ژ���[��y�~C��-�sv���� ݹ��DC׍<��tv գ$�p���d/�6�4>���:��Zy"zʩ
�=(,q�5�q+;,��~#z�q8�t��ܼ|'ޤqu����͠��W�vt�z�&c"�w�~
2*�M�^�NT�O�k�Y&���W���	�H�Tl�H��{���}�5�wǞ���Tө�X좥���� Ț��<��u�	XYsԉŢ�9��� "TB��
���"�ce��)�)���l��+)	1��64��n�+��6_<D����C����`�8���Κ��CmeUGr"t�W���sc�d�G�!��d�&��<:ULg�PZ�g�ѦȖ�qg�k����S��d�h����uh�t�I}^�X���惂U�>i�<\+�(�_ĸ'�ὖ`��BN���B@���Tp�K���[27��&Þ��owG�X�ۗKJnhX�F�q���K�<�������an�pɱ��No�s�#"�U�Q��B%�;dv����T�M����w���B�#Q��G��%���eSV�47q��\TYH��3t���9ǹ�K�k3�VV ����Qs(�������4���ϝ���������O\�0�}1BsV��/J�#�������Z�������PJ���[n���G���J�4��lBwGu�22�K*�pU魛���!��m���l�'�G��cfmeeU�pU���8on��/q�lv0}e.�}t���}D��ϟ/%�[`.Ȅ̍q�ȁ&��ԗ��ￋE��r� *uϐ���������7��z�sg�5��`�F�q҆��9'uG��H{���T���1J@m�=�˺���t�����N��=s�Jdk����W�.�A?ŉ�O!���hFx)�7 l�Y��\%{��p�f����u�81xmF��K�EM�mphE4�ai��1e>��V+��D��GK>>�H(�����������w0��������4?��X��^y�S��]�ͼz�j�^�,�U��ψgN��)�|�uG��|�� H��ɐ�N��n6��d�� x���"���`���o�@W��]t�	)�wG�<͋�~���e�f�V`�Y
T)�%�M��E2b5�飛�w�OG"0�A��>h�Z���M]�6�r�v����������/����h���yuE-tAo��<�Ȉ<^Y%�/F��.=J(T��<I{�����SN.��W�G�׻Rz]?	7~��G��$S�ȣ}�bx�U�<�$4�2�B�^��]h����z�v��f^�Ӎ�_̺��~Ќ N��p�����pM����͹���Vc��/e�VJ���-KBa�B�X �g��Ѝ5w\wU�(�/-~jJ�.�LAv�0�x���k���X-� �|�'�^�����jQ�ƢG�V�
��pf�5�����",�����JO��t<�)���h�)�rr]�y3�!22>����S��Z��]kp1
�:3�����켗�;�"��Q|5�GF�&4 Q:�D�ݕKy�� 0�R��j�[��8t�8�B*0W��[�m[\E�L���ftUx:�4D)z> �^���5֚yp�RJ@�8������`�^��>��r��-�*K��P(�<ǳ�o�p��ゾ�]]ұ`�����5���m<����F���c`��`{����&��V�z��ѳ �.�����+� Ԛ��� *��ߎ�Ks[�+ո�\3�����ni�;��2�4��򈴾�i;��5���>(/�����Aꆧg�ğ2��m�y���5I���5�M�n�ki+��wc������[���~�X�OYI���<l|2Xk8}\o�^D��c.�t�D�|v��b +2>�I��ي{{�9�&���#|t�}$S����� �H��߃��lZS� �Z�Y��t��|�I�<$� ��\��}�Y��k��}7�3�^3���YhRnۃ��.j[�˕��V������a�~(�y��gl�G����WZ�S��q��;��uEO�Ǘ�X�;�:8Oc �!n*;�����	Z���pMq�op�f� s��ߓ�����}���>�n�n&	N̢�X>���>�D%��Rq
a��][�r�~	�~���c ����7��^�J�q����9���W)R�,)'�r����0Lɸ������1�#�'.eϘ���=})K�ȶ��I�Ր�P��;n�0��+����ﶵ9"������b��MN��+�g�[�﹕S�����J=�j�	6R8;:����z��U<�3�UC+�Ԓ52밨���*>~2���d����/���b���y0��[�i�G�}��ܖ��^�����n[E;�Ļ�Xu)ˣQ��I�򼼼�ﭏ⶞T��+�\�,#����M�88�P�����pJz�d��!��5ZVJ��^�)U�nX���E�#��׉�u۽~���G�D|B�^�"K��<~O"~�6��Z�e�Zb�ew�l��f�(��s��s�[��]Bs*C��6Ћ����hTJ+{����:���<��9�8����I��uf4jdw�T}D�]���#��r�Y:��N�0��-����=t�t$n�1C�Y:b��Z����,��.�Ԍ!6�V٩���&�D��:���~��-:�B��������K֌�j%��jH���Ы:�(,W���߬�j��NY��j�=���[��(N�z �&(�xA!(e�����T�;�^�^�v��H�W���:��o��9���c1N
W����q���/?򹃨ʭ~uE(��._b��J2Ap����,�8�|+^o5c[�.:;;���D��y�.%Ú���F=8�?y�6|���h��T�j�,����k��:���=�z�Ʃ��	�����L޶q��m1js{�ѭl��iN�O������ktQ?��'���� ;<�� ���=������' ���H�,'C,#�!���9�.F~1�G��t �����E��d$���n����>�����C�1ϱ�� �� !�٥��?A���n -��ݖ�!�Tp1֬Y%�L����nII�1_un�����ߒ�@��y(m%���v ���7N���;�	ƻah� �צּ��u\fNND�Kj�T5Uv����T��s��7�qdǭ�}�kI���\���ѫ�U˙�]h�7��>G�qkr��Լ�t�H��]�j�5a�����T��R�?��ҒϴJM���.�9����!�4(PF�N�H��ye�W}�@75�#c��εA��d��+R��C�������G|����ww}�@o�����u;Ww3�|�t����[\mJw��+���CJ;�����8�
ԑ��/C��r�4�h�>��N.�<{�Ū�.��1�%ح�<R��⯊ˡNF��E�C�>���W���E�0ܜ�Q���{�g)omm]��%����h�+�|��֝
N�����<{�d�k"�ؠ�hϢs_@-mEm��b4����Ze����n����2rASԇ�N�����'X )p!�/�X���	�R�Lf�AI��U/� ����C(t�H�����D��p�-�T��BP�L^ 8�#�#���^��(�9-Sߊ/�z28�<sطk~�z�\^��Z�r���@��\�Ĵ�R'w~(������"˦�$��`�A{U�����B;W��U��lI�
9d�*f�s�	�z�^���rxka0JC��X}��z7�RV�j�#:��1k�+p�h�V�ȴ6$AO.V��Y����|#��80�������3��^�0z�N�����W�n�,�U����>q�I�0K���R*�Wu��˻#t5��;��Y�]ΜsLu4��xȹ�/�H9�މUlԕA2�}U����E9Hj���[���4H���d�N�I�D��8�Q��SiT�>�R�%�h�%�ĺ��p�dת�d,>��ut؃m�:��?��Z�CF>j�����v�uh�[�}n�p��ۿ�jY_��*�+��@�TC����Y��F����eiL��X�8X�CĖ�"���c8�͎h��J )���z6@5ݰbǭ��k��І�
�ښ6g���#ZMw�U��08�z�3�s��6�]� ��v������0F��{�\U�V����������"�l�J�0���r0�i�4Ws��ܠmd��#Vw����᣺�#+Tu+�����7�g��qu�B�۝9�Ë�u�ޮ�Z6�x%*CE��A����&��M�N.B������՛"+d�LSRWM��q���इ��42��F��?��ž��{<"Í�L���2�=�~"v�Hb���'����.�2Y��M�`.⽔}�D��1؞��y�g��\PO.�T.H�Ѭ6���! w����PʉJ�Պ�ya�5����q"k�� �t+��v[O�iw��>:r�Nպ �^e1a�-x�U�N*�b7��^��Ի-�=33�DC2xu�T�*��E�x�E�<e���6"y�� ��!3װ����c`��s=¹(c�<�Ū_��Oc##%�5�!�A	>�NB�\m<8�}�fMe�w�3��-V�))�Z��I���8b����n�J5�p
��%(�^f� �|@l!_�t����*6l�mx��ʊ�4�hqPe�bx4G��|+��<���C)c	�8�w��B\�*VS_p�tA����|����ӛ%�"ˡa��iZc-y~�@�,�f\`��B�Z@Z�Y�L޹*����"���~k�8��vx��Z�&=7��@���T-��%u�����J��[���}��g�AJ7�W^�,Ԙ�1'�o%����=�N�f��'P����D[rl��p!4�� �M�@��?4�y��%��J>���n���f�}�lf���,����Ȅ�~~3�R�F�g˕W=�G���k0����J�����&E��8/ �a �Dg����K���[��:ъzr�Ǝ5�6�*�'*�V��Xc��R�a��%��R�Hӟ���$ ����� P��
�����wpҐ�Y��GX����>�!b���
B����=�\,�b_�Wrׇ����,@�P�����}y8���A�nE�M��
!�"2T�B�J9�n$d(�����"T�24��\�i�*�4B�����κ�������yz����{�5|�Z����<Á�"��7� :p�*j���A�_1w�Yŷ�~��6Q^�,�@l,FgJ��{�1�mXp��k�����p�e<Z5 �Y�[����-����Uc�GCx�D�4 u�ސ���<9���.yu��ꑒ�H��z�{����w�h;���I�W�_Y��efp�U����N�A���{{=v���٣2�'oˑ�v��%B>�漀�/	��,�	]��H8eY���w��m۷x�����?yM���s@��a`&7h-_�|��F�6��欨���k�ˤX�ҙ;
���Є��������K�G�T��)ҝ�2e�f���E~	E^��*.R�H���8��6w!n���.��U~�M��-� ʃA-�T�5,�FէQP@�P�`�{�\w�{���i��1�腆���_�VM0m��Im�r3�oyyz~ラU��*��������A+5�K��P���������K4���6{t��P�(�U�w��{�����h�T�X�h=������(B@P��x����B�=�o��E`��mq=	�@�Բ��0��":���h�`X�)Jo�B2#��$��{@�$H1�Yy%*R?�(�6��XNӵa� �u���˗�TVW ��X|��˄D�5��^�%���X Q�= mm�U��Y������f��_Q�'(�?�݋˦'Xw
�Q�e��B��(�7��O6�H�T3�����B�@NnG���/.t��8G�|�����Ҍ4�2ʼDk�"�]�%vr�C�oșM=8��zy�g(N������^�����A�e+X���0��s��ʬSs�\\k���� `$gE��qKF��� Y^;�4�y��k��W:�ϱ��V�f�:-m8.�n6-<�h��H�(�.Ri��U=}k�.�1�l`�/d�H�+YH?Qh��}:x,:
I��=�E��Ӂ�e�S\���6p�`�޽��䏘����s1Pi��H�T��H�����p�v��	���c��H�e��0Z��=W�
RoO�����xF #�@�q�Y�W�X��������Gms��^��NЍ�e��O��5|i�G���uv�:�X���`�sFo-D+��C+">)h�pϧdV9V�7���چ��>�20�YX�[����T��6[$��i��aFo����ƛ�s-}���RM~;����)N�����a�״�Z\ć�/��z��M��kE����z6zr��;~�]���!
8�|��������g	�fWykQ�__��6���F�{S���:W}֩�J��fй�^uVBh��*~�u��,��En[�WWo�Go��'���	)܆�ū��_LD��񄾣FB�u08���9G��"G�=g�k�}{�v�G��5Mj|{��:+� 0�e���v�H�#��+B'\+��o���B������F���-5HZ#����tà+��>����霡|�y��I����)	�m��c��MY��2��M���֬' �i�}T)[Q�z�_`�p�r�o�
�d��%��6��h��S�����k�Ͳt4�NX U�@#��>����`u�ge�c�A�	ɒ{PQ8&9���>�9M�|ʝ�4�PnI�e�Ky���r7V��],-r�N�tg3��<	�rp�f�M���To�0C�9i�G�7��M�{t�9n�B�X�O,v��G�K��5)�����[_DM˨mdVNFM���	'��Ϟ<y"�֎1w��eS��r��&n6��w*y�p�ae��`;��$������l��c
� �.ִ6ƾ��.�j� �P+n3��$Mz���:��i�m��>�P��1���( �A.��o�3����!}/4~Ch���ݽ�9��Lk�4�ۉ���GT+V�0�j�g�h��X�b zy�:�o_c���6(����9+��O1cD���5q,�G��J��[m��Ҽ�s��pGG�������MS���'�^�f��lV9,+�عs�Ἲ���r��z�D�\5��t���k3�3��h��l�^E0��W��ԍ<�ɫC�%u���7D�y�]ζ')���6������j�'�� ��S�M,���bm[+�~G��5!��;���2�^en��F�㋽��C�pj�Ĵ<m'OOO���������������K4@j����5����J��1kz�x�'(4]�4!e����f�W��i���J$�����G�����!M]=��߂�}п6�H��V!�f��L���YdC����܇t�I�~T��{2h�M��V�{��¼4U��gE~�s������9����}�V��
���u�^��!�Oj<��|Ƥ|鷧�V�(�3E�П�a�lcW�c)<�l���N��,����B�&d	��\�X3,�8��9�4|����f
̟�H]��MD����3�x�.W|�bQ!�
���s��( 6���,��:����w i�`����h��:��w����O���>g�@e]�d���x��|r�#,�9���ـ%��(��8y
~�L&h$��;��]�?�O`{)� @�3��4��<��ƍj��]3�Aɿk��yid����D�-��,�R���Cy������t��9/鷏i��RӺR��O2\���]��Q�����\���A�AEE��S�6��yڟ��%A�����M��\����C�+h�K���i�������/�[@w%no}�&Lތͫk�e��N3;9��T�*?���7�� r̸�`g�]q�ǚ��AT��:�wff�N�}LH�0�4'�OcxK�6V 0��6��G��ճ��spt���GD�?��8v6E�7�WS��ˬU��ה_�<�V��۷�)�v�j~VyO�c�ɶ���|�خ,�.���7���k�Y��v��Or%�7\�k���9��ɋ���I�M���I���W<��[��6}򆝽m|bbb�\>��c�p�K���6N���k�f}9	����2|�G�U�;�Pf�w6���9ԏ�_������r��*�w��&���X��x|�s�e����{a�����	7����D�K��U����S,���D�9��Zѱ{��Q�+(J$�ǯl��s9-�� �[~S���i��Ȥ&G��3�+����F&SH2�����ɛ�x�U�o.e�ت�������][xHSY:�.�j����$NI�OH�1��,���MΫ�#aâĔl���4��T�vb"8L���%��`�������<�B�s�H2u���,�e���a�jEEE�|�i�}_�^%�m[�AY�R��`*�~����,lf���\jU������~�pֶ#0�X)���6�o�
l�Ý�*8�}p,���ƣu��|��qw�=/�d��m����&����G��8��(�sƮ�X&E޺��!8��QW�M�A��)�5��
*��ѲC�CQ1#1&��*Al�-��>�����u�/?vO�������$	"A �f4e+0��E+hx(bEhOh��T�+?���e��r�@�K	�����ڟi�/X�9�u|��౏�tO������෧�@� ������t=ȿ�ŻH�bY��Cx�D1W�� �������Yw�{�h��!Z(P3�P���������_��)�\�IW�	����=��\�Bg�H���E���"�����SÆM�ƚ��B�C�He8�~���U�0��s���N:�Z�P����a�򴹕�>TZ	?�Z��|@N�P�b���1��M IW��t�a���=^��j��+?~<���e�;Y啠W<d@����n\�V����@�i3*�F^0ܼ��";�����I�U^�����6d�r���9���~wFk:�H'�EM�s���g�<��7�X�̗��d�J�!R\�n�t�a���n�u�ÿ�͟�˷j�OjO�+8i���x�M��f��:A���P m���~��?��
gf�\�K��8��2�<�<W'�����:����~��B�kS7X�t]�N2���ŨE> |�- �H�0.l��i��EFY,�ʊo�T�i���8�b���?}��Y��a��)��:#W#�ۘ� :,l�)l���T�y�?/����Oi��e~^CLe"=�60��?8<��<���j�K|�o����1���f�v>iP�r�-[��Ռ��9c1(�����Т�!�|�y0���`uCg�v6-e�ȅ�X�U�Y��+���0�+B¯�uy��=�% G���|:L���vo͟*C�����R[܅��mj����י�_�u����>�i3�2�����yg����g��@���i����,&&v�����|-�O���7PH/v�̗��*[A;����j�,(��`����jjj� �[�Hj҅�嶣���gD�s���d��R����������\S�8�������O��<�>�E$�A�d�w�JR��p�����ZFC�H> 'ܗb��Xn=�~h��8Y&�����b��<!��t��s~A��n�E�+�s�rY>v$Z��o�h�Ι����@�cα�g@b}����+?��GA^2z��ٓ�tvt�
� 2���<Z�7���ٯ���x�,�L�� ?�pW6�0�$WA��.���'��1R�Bs3Sӹȥ3�D���H���g�Z3��=S�o�ㆇz�y�� �+e�Pf��ΣR��nƲ��#����G9�
�p��o��@���Z�E�C+�	]6YB
R�$KɄ�Y6߃)$��t�VX�h���S�R���t�a"ݫ�!�DpX��[�����L�%6RO�	m �������;qGGGa�X��`��4o��eS\�ȇ�i��.��UI�K]g�;]X�2ǟ��v$��Ejպ�
!��Bձ/�=�P�K4��޹Գ�r�#��=j�`v��?��`З�@W�����̬e�"�7�қ�j�2�#Z��}�wQ�� e髆Ic�@������/I^����1���������6]j��ݹ�ݺ���=h/�˃Q�u�gL����+�.�biۺ�-  l�nzS���C�
y�0����
�?q�"g�s�mk1��]��ZE���!KH��޵�:Co�5%��''��
m7�FJL'���u�-#4nڔ����W��YȘ'�@�A�ԱW�N��0o{�v5q��x	Sj~�W��k�W����2;Z�%��m��u�q�2��*�r�;���L��)-���R��iQ����!�A�������>���"Nڎ��n�:���!���2ڗ�[�ܠ���z����k��W�K��v��'��=>�7gj��0,���vj�mU�
E�Mzk��b���
�U;��]42����pR���0���ɯ3 ������_��)���@B��gFik���`ц��r?%�U��>X0K��Et��*}���cir����T��=���bt_"��`���k�չ2U�X��n�U��b�J�m�dh!,�D@91g��	�[N����J��e��������Ҽv����,��+W�5g�� �yu��t��I�N�i�c!�1��T
��G&>ŜX��D��T�%S��W���6H����i�+�k}h�4zf���?E�t�W�$J]OA��י�aΣ���v���`��?<����eq{�ƞf�&o�����b<����HO�{Ru&��.g��(-�.^�25�5E�ґ���=s��4���'�c ��:���&f3u�\������R�3P�\:'P�UD}��C�c���⨧����G���>S=:ŀP���fͮf�*��ehFݫ,/��0%d꒝4�iN-W;*�M]2���*AeM�t��5 ���bfp��Z:�lQ�m��2%��`6Agw%W!��?g��mxrU�����S���ﭷ�ĘG��fwFo"�C�)�8�}}8̸����������eoO�d���R�~�F��=�?��9͑emĐ�H2ϡۄ~��3���0jE�	h����F-p�5�(���D�@�(ԒD�W��j@�����c0uX8]��k�^�3��'n4	�����Aׄ]�a4�+ ҧA���d�.����Fk�Lؘ,B��sm3�N�����p�O��Y �$��v�S�U���E���dӆ�x
z�ô)y?�����VlD[7�$X�u�Y�F'C-uYTa��Bh(�� I�Md&��Z�sC��������l}�r[��*��YWM�B��&C�2}=�HM
�%Q��/����1`�$�p�x�H&&f�O˂H㸧�.h�[�N�.?{�Q�0�n坿^n��J��ī��)��BH*�ð��=k4�~v��0 �g�2
��� y�:Z�~г��1tr/m����ڲ�ߩhÈPҦ`F�IJ��$�a�nUF�=��cZ�}�PW�!��`��#��w4��;�o�IFrh&E������3^e�<�����K�G�p_L�&�Y��,����I��Ϝ3������)�J��x0�J�k?XFBcF�q�9�

ȌD�i/��P�_��,��=(�4��$��n�����\SHT���Ü;'R�a���4��"��zud*�����H2d�q�U �`z�^Q�@@��6�l%�8!ܦ#�54�{1�����E�v 8�8X�t!�s���w%���NE�Ǝ>bqnc�r�-�I�Ou����{���^���ՅR�y�=�a��s�f�p����Pܲ��r��tmTF�b�nOˋ���I��g�i��m������񝯦��X��q%!�������O)�.g�5ly,�������2In6��G��浱������6:� �)���ϒn��P�L\-WzR��2�:���q�P�� �3����NR�2��1	k;R��࣯搰�3��r]�	���>��g��u�#?�6�=�^O=�Ӣ+��xgE��2F	r���J��MF�y�w�J�G�N�BΡ?ƿTa�@�4��-33�.[�u+�h�Xd;C�'���Ƹ͓ʦ����Ԃth�n`D��������h��Cz��-w�}O��I�,�յ�ٌ�\�Ο2y��p�8�%�� �g02x�*���ɴ��`�"��sE��Z��Z��xX�t�ԁ#��`�Za�ja&Aii5�@��1n�����c�C(�)	�/\p�����Х���"��3u�!>l���,s������ѫ~�ɯog3��bU�'�*~�t�}��|�)1�A��4�2�s:��
��`�˟�ŏ+R �d�"s1N��a�0�Y�XS��)����<���.�L\��n�	z��<p��K�Ǹ1�=X{(�_S^��ݼxl�X��T!�eF�Hʳ� '��j���a6Y�ы?�\겞^}xd�|�)��b��[g
�yA����tj��'������IW���9�'��,��v�n��|5����_���T��N�������_���Bq?�Qı���9�7��ޟХFgT�9��B���4�%�i
*�_����*]��zsl7y�q�8�9���]�Ջk����׌=�i�$:�8~��_��s�D�|�(�=D�K��Ɍ
�yXϼ.pC)��v������1�"�A%�0\V�꿊�qW��4{ܧ������?Ĉ����?�}�d���.(��/�
2�4k7�R�?�e=���T���(_aY`7��~��N�/����z�0#�&�����V�̣Ӹ��~�3 ��дwM(˶�LӋy��H"���i�����<Q���?�R�M���B]���1�ni���.����%�(8�v��%c3�:�(z8����ĠAjغgW��B�h�؞�S7-M��d-$C�%��BS��	]��)��pl-vkkA��1�j�[�$YL&ꢹ��"����< ��ԫ��yu���"N�Hҽ�������ƃ38kg���I�2�m�nF�&rD�4�g���	],:�
S1�o��_�V����l�X�'9�mp�m�Mx�mZ���%Ff>��s���\Di��Yk��t�,�R����	�Π�>ұbY���X�x�q�=����\X5Cv�S�K��`-\J'I��gA��ItЅ����9�ޣ~�=�}0���<�eF�I��X�h�9��&[��U�
/)��D�e6M�q�}\ޏ_N�0�~Q&޲��|,�x��T�c�n�%�f��ɵ�g�G���0LCW0�CCu���x�.�Qv�0��,�Ĩ�!m����1>"4��_����l�cG/�sPd����[F'ʡc0�
47���y����d!zk��	�Z��F���{�8���oT�g�ۉ`i�i�|F�K%r��z�P����b_d��{ۄ-1�B�BQ�2[�.��XvΑ쩒3j�k�A-�ɚ�k�֔��w���w��9:�~%��
2��?��q���76���f+0�#7�|E��
k`"d�Ut>����`=Τ��zL�`�����<I�մA��<����e
���� ��Ⱥ�Kb�kX��w<��k�K�%�T�g�s[�o�=]�3����d{���R���Ċ WIV�O�	m@������Ցb7���R_w��P9�aT1* z�1�1u�h��ׁ]����� 9��.�S�.�M�/	�N`�Ӆ���S�q��V,�9fL��u��V�w6��ְ~�%s]���x����P<��:0c�&wS�����|D�ٔ�J2�7
y�,Z�9��w�6��uX�����DC>�V�ň1���tj	���+@�u�egh�	݇(��5~�^$[�y}��\q?*�|\59i>S� ��5+�4Kf�(��o{�N�F<>�G��qU�ת|�Q��1Hn��ې�������`��<~:�5V�� �p����94�OC&�O:6�0���4y�Tϊl��Xs�	�CX���j~�`�<�g$uwdu������t�ԛ�#Xb��<���O	c�+O��G;<����  ����e��2}���8#㊦I�-f ?Ӿ���,fB�)wK��VI}����ֲ�%��D�3�}�Es,@��e��~1Fd�so#��)�➏";�ύ~͆ky�I�C�!gv�(���v��(G�l�lz��t'i�Ab7��B�~�% �)&�� `�h�P*�q�DQ���1*�	�6��Z���54T� �]F�і2���N?v��o��R��ݦ�\��{s?ʹ�p�1����L0�����;��pm=��9��>2�=�tE�vl��T_/�����02 $��bE:X2�o���ج�^8�F��4�g`�C�� �<�ݮE;CqBG�7�`I������&�C"c�� ��MR^�F�ƾ�J���leŌ��3��4@�ǶȺl�.#Rߨ2�@�K2ذ�MN�w�UX-\�!�;N'!�i�t{=�44�8l��N����8���x��
t��f�O������d$a֘��&����n�2c��#�,2J��_����u���2~�<0��|�%v��%���H�	�r`B�������o⒁>��F�,mF��� ��o]/�*J:���(2�\^�yz'eC�����0��0]F�6jSN0C"J��T}F5
wm�y�L���1��Y��8�⑑���J	^���b�vn���tܑ���Y�QM�iz�y�����[���%����r�5�I�y�����kd��@�sCH�R8`*L�Tn���R�d,6 Y��Ѳ�����sF�9���'��p�
��QFG�s����,��]�9
9ʧ0؃*��� $�ֱ?�pR�E'3�6�ڇn���}4�<3̺$!��Tv�2��B�k��[��sR�͋fPo�8.{ ̽p�q���y�Kx?j�������e���!"�eø��Z��
�2W�B�%����/�Q�T~�s@�p����#��Ԯ,�Kf��s���s��-c��41��#IvB���ehwP��!%����N89�OV����P�v@{��O��n&�ȍM����Y�ɐ��N�%�k�ǚ��:��VCR�.��~��汎ӛ'\��73a-^)ZPP@����Xz� (K�Y@-(F���{���1sb�c|,di:(}���a��M`-!):;�]�t�"�s���Z���Mx�F��z�׭��A���t��(B���닦���ۯ�Q�.+����5���c���QD�M��͔a�Ԯ�>z}����� X�eT���c��9f�w�Y�i�''��wM����^�`<7�	΁�M~xn�?�z
��rT�q�#`ƍ��SOf�bN�wX%(=�1�O���.E0�i����{���?L�ɓ���E+-����(j7����x���i�����|�#눉P�I	_Q..�a~$_�+�c�Z���:�S�-�>�)�t�uy����k�M*8�ä�R�Y��MD�X����s?0r���0����a�1{�M�C�pm j��6-�:
���@�JNc�,%ch�g�6
q�C���B��*�@�k޽bɮ,%���4ߡ�Œ<��y ������A1X6F��+�"��`|��� ��R{2�o/��|;��(:ɗ5�3I��l���,˦�3��(�����/�*�<�$��C�$ɤ��gM�eΝ��:Mc�ER壔*O杯m��9(B>2ҩd-B�����(0�L��ܟ�a8�Q����4�:ЀI�{"��֎E��{�zV|ƦE�2��'ѵ��r,tR>2�m��4�c��[�)E�|�I�����za޵�~�.���&!tI��œa&�{3����G��Ү�!iZ^>�`����K}�^M�?x�(M�Hn��6�/fU`']|(���3Jt�9e $8�6~��
*�*+�yx�T���ih����@�<���;jڏ�t��֛50�1��N#V�gx�;�Sʮ���y�u��,�A\�B���հ�	QuV��ڝ>},	i��B�G�_��E�/�����$��huG���3> �0�e}d��ܷA��~ּ�|"�e��ݩ"ő�;���5:�+K��8�nQ@�]d��W�QwC^��̗��@9�Ck�g��`���2�N'����(,���3��P�e�k2����ܨ�\���k'��+��ۅ����h�����(���$�}�cc��?B�f9w��C?G�2R�'��X�6��6��O�?������O�?������O�?������O�?������O�?����9j��]��wN���\�	|��g�|��)�EV���L��ȟ��)�׸^�}`�?K{�c|����8�;<�ϱ�^I���,+�/yC��R͊���T��5Ͻ=� �og���wX��'1{t��+�,��2�7�X��1��e����0��1V���m7�W/�{�ߋ�^����������n�.�E�G�YЬ��߻Ã⿔��L�z/��N��&/�4�B�y#��fqqqUrϢRRSk�{�ZBۇ���(��Z����Vmq�{�nk~�[H�����Ej|/�5��4���,V�9�I'����sDb��_'3c��0�+�8W{p���r'�4�nVwuy������qq�8��o݊_e�5�+��ѣ�.��-ء��1��Zf�{����y���͊ϟ�����S	;yE9��J`mwسG�iy�~.�`� ݭ�66�QF`��'O�f͙JHp��`��vbJJ�e��.��z[��.ꑫk�:/��Ĕ�${�<�DHG�/++K3O�s�}(R���ߐ��/B���f555U3�u;�	��'c⋻�������۫��Mu�~]���}��'����2vt�9C|��E�S�ᩭ��-�Z���ji`b��#�x�"�}ʔ�ӛ��:p��X`�Lb�<� �g������S���:u*9--P��#`o�V5��F�[�r��AWH�8���8yx(kh<����~����U�-�3�O�����ʻ�g#&چZ�/{�U���)x/%x�M�M8��VF�X5���$���A�[�1i	�$ܵ��r�[EOmV�2lJ��Nk�/N�}�v�$ٌ��Z�St����T1�������~)R§ha�u)�oԓѕW��\obB�R��=k�aǎy�'O�w�m�A��X�[�r��9X?�(�����!׬�ٓ-cd���^�[����!�:4�?k֬���j���W!t	�p�T�:�v��O'(Xs���V��L�I`%+���<x�0�X�/r���}�����ʓ��W��^K}���T`'1Å�H�G�޾�kd<(5B������着���^�K�O@�cv���G�[&=��򺨦�܄P�)C�,�;�^���F�S��^����>~�T���Z�q��6Y�x�%���_��ӧ����O���j޿�'�D,`7�����3�P �P`���@�S�� ��{}	ݦƢ����n�̈�.Y��>i6� ��%���0Mߋ���MVj�M�6pk��$���G���.����!�x�͛7�}����[���V�H ԃD���t@���=-U�&��KU�ѹ```pYE�$�"����9��N���5V�7�������N1e�Ci�����OмOV;�ƍ�ܚD����$�,,�
�[&��X����Z��	��&���eə�3y��%^?^�hii	�_^����6Q�Ԝ+��R�iZ���v§�$hT�%-{}�"]�����$j��ː���_���$$[��u[����)�bw�v		�*8�y���~N�" ~�����6�bMW�L�ʿ,{Y�w��}�)���C;�?�嵺⧺�e��8k�e���D�oD�;�p�a�e��S��!q�zn�����D-?"��5)6DL)嬌��cn
�B)CɄ-�畔�Mx�/mve{���#W���G]QAA�1׫�:����[kRk�����j��j$�W�
o�2ۓGf��]��+�E�k{�����RI�(��b��@����x��\��ș[Iؽ�m6gř\���,_-$�='��<�j����B���-��࿴x�G[�Lיs����T��:�8��5k�f*F}߀իkZ�Pw\]]��ൄ����m0;cz³�9�5�*u$p�[�# k���UQ㒫a؜u;w��o��̑y�f��V��e�aª��Ԙ�$����
���R0�X��������U��$ڹ�5����W����e�p�r�)�2!4����'�Y��Hм�������Y�K捅�=+�@�e�N�nS!�6�R{p���1�o����.*�{{{���}�P�:����-)�E]}}��+��r�q���i���s z	���T�Hǅ%L�ˁ�����]w�q������0q"�x���\�׷�Gͅ�i �C��� �_x\�d������A�r5���ge��$N:ܛ!��B�V.%�T/�M( D�U�JEE������v�{෸�h+��[_\߉W��r�R��_ ���ոq㪡�z��_���^5A1��ʰ�y�&rr����K�WyT�����[H������h������{dr]w�Z��Б��v�CtO�{��FR�A����,����m�$E'���[�� lߑ��5��+��G��Ѫ1ah���T�Z编���˗W�|���f'H0���]9� y�**g�;���-a�_���������n߆g�kwI|׵e�&&�h|o^�{������:+�d۟���F"�)�,�5����������a���2^�I)�Q2t�u Su4kj�?~���R�
��Ɛ�v�Ty��L�w38z��uhg$	��W.Y�*�D�z��5�m�����RE%��W���yy�v�V�={6�Dc�3�M���OTp"͍6m���\��<�`2L��2
�E�V� ȁ�MKR�L�4Gww�}1[���Sx�8L��0L�PX]mA�3���2��]�R�w<0����h�M5VZ�A�𞔼+g&a(��Ok:�)�g��/7�<�����[&ݴF�zw�9��uJ�C��9�,=Րm*P�th��K�`T��:��l����;!���hEV�L�|�+`l�z�45//�$I����;Sm�ފ�i�6/rڻw�Ƒ��ߞ���s/�Ix�����O��z����Rww����(T�Olʥd�Hk���.\'
6�����	�b,--�A@U�lx��h�%��8�Q�:C�Z_I299ɁL�p� �hv��e�'�j��qD8�8�@g�W�6߬SxE����mA	����:y����	��P#~��	b��x�����LHlhH�l�m�t��mƠ1n�e�#�)���x<=��4pn~>8��������f}9Y�;�j�N�f��f�i�ƖWV��5"������긦o���O�.�������2�:��ᐉb��lJ5�L�8B���5�6�1�_+4��T�i�t,b�D�E}�poO�{�&`v��M�(��wB����Қ���֓TZ6@VN�5�g�m��p��G�A�^٥��cp�:�q��b��-)I~6�!�P�!6�0l]��~kI�_fα'��|�ѹᾂR��p@��&�^�I��Zσ��WR}� kwr���pV=<<���;̜V�%R�����YC�9��0�"��qw򨌳�|�	Q��Rq�]@P�J�` k��Ac���D�/7���!��1�'De R�����$�~��#�i��:��A�V����]��{l���_���nȟ]�0�5�PS�8u�﷧j�:��rݛKZ&e�u�ѳ2Y��ga�Xjp��;�!��q7���c����(�=���P��pt�^?"(�r�ĉ�PW�����O7��Z��m�	V�^V�M�-&\}�L���~����54����7��p��?�i�osjv�Yy*Q*.&]���'�m�J����[PPC�~��E�/da_�
_��T0rطoiGC��Ƒ3i�)V��{�����9��A�O�������{x(���9%�R�w�qO��-�4�G��S���9:��o�/;faߎ��+x��]|��Vۀ�^�l� ����R�*G��F#�\[�ڌ1wEr������i���)�8��+,S���Fao��uW�&mS*�IE�&韕#Cf��߱�cŊs.��������E�O3�H�]E 3���$''�LZ����EUKK�(��=%2��j�,G�2�"I�Ѷ<�z��w�����������j��𠡝�`���ܻ��5�ܿX,gde�>}���-�'w�v;�/.(P��F�%��כ�0�F��%��"Z�sK7gXl���v\qA�p�fr7����]�O�{	� ȴ���KJ�H���L�I�P��_���e`�M�2�^�s�8�v,^S@!��7�?��_(ݣ=��ӵ���kjD�����~9@�u�^^w�ϻS��AbAk��e�v��F�I8S��\���+;98,�82�:�go+�K���ؗQF�[�w�w���
<�
�O�̓M��Eو���5&��|�N�����g�7�2���r�.@Q5���O<���Z�Ǥ"��X���mڍG[�^��� qKϭ���&L�� ��s4��j[Mq�U~N�5j�͉
^�ˢm�2͑w[������j�4kI�m��Gd�8}U��{�����&���=>9e�_�[7T��]z�r�����#A6%7���e��k�������0=�g��1�g��Θ�j�`4��.�Q���l�ƭ�괕e4�#@��C���[�� �g��Bn�9<v"���k㖻������p�IY�g��FR����y�¯)p����D0�DyCE���M�m��Ձ���>�'՝B�P��X�<p��ev���&lx:S���uX��,�����#��]�~=ס,�XČ\�#��3�6ų6�Ed�nV����h˂Ѐ�a���ǩ��!(��}|k�ǯȑqkϢđ ���$�I�6J6Ǭd7�Vם��M~� T�08}�H ����\��6G;qU�s��.�������|����H��gO����xz~�|�U�b���2"{h��\�o+5.E@�Z��Ŕ����y�[n�e������z".�1���4D���`���r��{ 404��M����Qн�s�
ϛ����92<������|]V�g =u��B�I��LmX��O�&��\�S�) �2f)i��H��C}���q�4p�f��s,�ݻw�؜
��R����?<����0�e�i}?.[X�4q����(KbC,������2��E�Ț:y���9�DW��y\D:P��vE`l���?���e�6]䞱�;ĆkC�"��Oy�+�s}$5����꿂�!��m�\2e��V����_��7��1�ys�8�zHA��|�`G z��1Wau��td�4�X��zz���mu�VW�����;�2ɍ�xó&�R{vB�Eְ1�D�Nr�7���'�aT���Q�q���*uV�#��~�.��xu��d���qϝ� \�
���8�($�W�z��-�����2��"�KѶ�����a
p��Cì0�d�E1eU3�u=�^e������B���6b�En��tWhv��G����l�vuy0S� u��a]��G(	}���~H�����Y�g'%%��H�?�Z=/�����17��G������Þ�h�L�4�B��� ��9*��׶@���֚�p{����25I�ڳ����V�u4�+��љW����;�Y��;�=8���P���8	�!I�ҋ�������C��͗Ew'm^�cVYD;�f���$φG�e�Xuؽb�ix�;`M���`K(�K� �V�@�?!Wy��9	��>>���PCJN�#��zs����
�+�O]*��c�DKuhGa�bϘ9󄩬��l�ۇ�V���Ӆ �	�j�hQ������eE�]2]�x9<��
AA�v݉8�hI
���Gڟ
��ٕ�����R�5��ŕP�A�'�w�Z麉��+x#>��1կ4���~�����d6΢'��a�tY68��M~�*s�����d+���i�+u��5�Z6��:(V�ϛ]��n��!�x�	ѹ�q%��TU�v�NduzV��/�� EFkC	M���9��	6{�h�%o0��CľUYGfUB�B!ۀ�-h?2���@g��ۺ��Ya��v}��R�|����d�5]a۔�%��l/��P$�����/C��a6��8������B��f֏w���7�)�U�R��k��{�g9~"�!��5^�������Z}WXgN����?�%��}?%���$���w>^�:m����&,�Cr��0t�TE�5"Ϭ4�}}����Y�=��٦ T"�敆�,|�s��3�FqP;:}����% ��Wx�+�݋{-~|�s�I<�܈D���q�ф��Q��ѝ�q
y�� �y�}�xVO_��!QL�=�u�[u���8�@�2��0d�J�U�xN��6�T�������F�m;�l)��^�P�1�^�����vg P#Da�<������
�D��cE�:�[��/u"�*^�N��S!��;$J@OV%���
�g�+��%T�/wk�*v*e�x;AQd3mx�Հ�(�7/����l�w�p�L���g����kA췞�Ij��Z�zJ����ȍ�B>�K�C�R%@x����A�@����cm7��I�ȁ�?5DL	1��1I�?�)CC�ŔlL���ؔ����M9EtІ^F�S-O����8��"��q}�v�u��u�}<�x��8]��)F����i2�~�ɭ�j-O��``=w$����V��Zqd����֬��.x�q+Il�{�^��-ud̪��H�;/���'K��������?,<�hu�Ĺ}>����{본<�֮���\��
��#�uG��`s*~���T�~H,�H�f�c�62�>Rh��j��+��Kh?�h�O&gԚ|� �!N��߉�\���{���@����P L�����x(�P�j��o݁���.
�5������kE:�U�y�׷����*��N�N�[!V=y־�
��P�8��mZV �|��b�
#b�Z� Q�8�8N�=�B�S��Ʌ��Cu�.R�Nlq�$���2�P����A4��B�
�H�j�Q۵���ׂ�-�����˗GC/F�Xy�&_�8��JUU8����I���M�]�����lJ0��-��?�ta97h�^��X�V'	�\ח�����q�)�@�9�VDo�����H���8���K3ߴl��ܚaQ���W��VX���ΐ��$ޙBW����Ɏj�.�$��?�5��
�)&e�+��P��)��9t\uE˯���^儿S��wV��Z�����qn7��y���/��0�Ӝ�o]����$�{g@�*�)c�kx�b�kDE�ԆNN���%���MIlҋSH��wK��7+ ���6��A��^�����5<l=v�o���2��kq�C;g��ld���%�SG'���s~P��|DP� �4�ᩱ�U��Q�2(3�Yۘ�M$\�*v����Oؤ�k�l)��]����<<�KiRQ�+����1CU�ii�j��b��������$�?���7�īk��	��z�q,݉��?m����@�������f��+:Lxs��<��[3M0J���g�م��D��GEb�G[Qc���P;��������a�ut���G}iXE�7��m2���OxFHҙR�X��#���Z�.�ox��U�&���lnj�nuo�D&���Hv����H�嬬��N%�H����%�IR��XU���f�������B/yh���܃���j����gE�����A�.���b�.�ʱ��T3Qǅ���LL<E�򛪶�\d�����>�/@�Lg/߃����`�%�,i�x����#��}�ȲI 8v�{s"VWqy�Hy���ȩa��d��oP��i��c^헎�5�κD�Sq4���
\U���W�~\!q �п�U�w�3�xrժ`��}e�ڮ0+���]5I�.�[�L�i�4�4��r#ɪ�k��g��,�S-/�k�&�~Nk	]w`�� u���x����tS�<Gҽ��X��e8��.|��ن���@ed�^9E���7E!�<mZ4�T����Y��7��|sm��������׃+7 �VOT�5�?����߿}��Aҍ�)����17���|l,��bɗ{��ū5�Ll�aݒ_����Mn��f5��$�>tR�lc��x���ă�P�ڃ
(�0"�!V�6�nx:|s̵�p��ت�A�o�����x�_x����s��?��%#���#�_�I ]��:z��K㍖а�tt~B�
-6��h��94D&�as��c��Z/ȴ�qx"��#��ǧ���be6�6��t��V��4^o3|��1�:簗�r���N��i%hh��o0��hy��Y��!��;�w$����z�|�C"�R��!�q��7@t*R�i7�����TD@p�9�;�?>Uk6I5M8	B��뇲$�̆�dc�՛�j+��h�3t���J��7�A&@�z��e��D���-���Έ�+�8tNF�Α���p��$`�Z��_���o�?��@g��Sc�
�������_�"�l}{˫<�^3��V:S+y$�ƿ���js���0�t ���CWg�캂t��F�0&��@�@G��)�~���\1`��;;�y�bڪ�m}��-���M")y��)��k�8�:�8����d�n#�QyQ�e����`{�I�5�f����1�x�g��X�-�D���D��+����f�	�����,n<鏿�4��{�#HI^w�q�K�>�;�|p0��͋p+�},?���G�1I�uP��ýY�/����'&a�OA�k�(�U����CƐ0��u�z�������.�o�B4���D�9�]�$���U�-HT+��拂C�A�X|��X#�	}�Ԅӈ{��> P����OI�/�l�~��2��g�i�¨� �#n�����^�|v�[HB;^{x�M�E�g��?{j��I@y��������~��Y�Π7��}���?I��ct�?��_;T�&����/v9�ԡ����-��D�';g��G9Y��aj�l������kaY8i'4�!���}�d�-z���x�p�)�6?'��MZ)�]�iS���eX��9z�5���L�e���4z����b��o ���(����稕�^������X��)����"ڦ:<vbJ����Y�M�m�ZY���y�u�����;v,�ò�y���-� 쯲�	�o%����q6�yh0~�g�������h���8�N��8���Y�YE#��������wOP�,�Ǔ�8�ՆmHd.�͈i�lK�|>ڪ�%�U��;�^r�7H��F.>k��u��D˶։��܋:�s�k��xp����Rd�����x�CP�2�o,}��y�I�m����J�K>��aEy���(�]�tIN��"}�˗gߔ�S�q5�=�(o� [}��kd��:1���*���Z�z���)�D�����b$Zu����  =}W.h��:�6��w�x��<�t]��Z�'���u:�K�{oO����7��4RҌ&I�ml�"[٧	'�m���)cEؑ��2�`jڨ-�(����{]k�]��|~��y�?�W��Z뾯���x�C�@R-���F#�>������毿��G��8e�G�bo)�k�͒�j�d��	r!�N�F,�<�t���e�ö�|�	���d���g������B����a��1p}Zj�S��o��J�+��>��e'��/k�,�}�Kx��$��?�L�	��V!���S@Pe�wj�=NoO��a����?T`%몖cʚ&�~$��p�}�k. x��kY��/�qD��L���l�=�bQ�#~-�p[�Hw���k�O~V�7� �#�"�L\�M~n�00m�1N���Fp��M%�0O~�u%,�^�RQ�w��ݎ�_�V�ۛ~��iJ$�b �`��-����������x9����,��Y���?*�5��W��tO޷M�����<��;�B�JT0���K�6>{���G��M���v]�Q&%e�|ܨ��#{����Y�n�],f��'�ǩ����=F�\��P,���1MX9:t �`��u��>֯~q���"eW�7Wa�&ws]�4L4ݢ�V8�T'^��1w8���!���U�g����$t~�^�ʚ�j��n#n$R�~�� �%;~	yۚ^�:K��p�ݪ֪
_D5�&�p<H3��|Ou�Y�tv��bԹ�â��͊��$��}��F���}I.�P��g�z,����9¤�M�o��-� A)�tT�.U�l���o5�1�!���J+)�h��v��t<�3ޒ����o5�����{8�8AI:���,���(�@Pt{���Ȁ��b�j�2`�GG�]��+U�
b�zKe;�� �I!�Gp�J�
fw�Up��ُv)�]��i�R{Np�/h�*TvP�kd����n}���2�q����1��w�&�&2���}tݶ�U\�M�gO����W�3
�k:�U��;>w�K��J�8?�0�Ӂ�D�YzG�}�����9��3|~�+�gC�蚞���uD����ϩ���Wf�S�f'�G��jC�Jo�0y��mmC�1T�ǯ07F&e�4�3���^��95��Tx���X�Q�����x�ķ��%> ��Z?��_~�i�%�TS�Y0a��<�]����:��c��;�pi+?Z�x���-D�Dx�d,>�Y�MG����e�?s�{oA�ǩ؀��+�,�?�n�$��_ٮ!>��Ҍ	$r��/�NgT;?Z=ah�n����+AP�IЙ�w�&�A]|����?�����|��9�N���c�;ܤ�>� �W&.�V��t�?3��ZC�z���k&�\�5uճj+�DD�	Do��L���?���x�\�I�t>�<�� �[���LT�L§��n�h�:9u�,�D잽o���U.�S�O�x�~K�f_{����l���RG_I����/V�|�J��x���R�D6 $��P���z>:֑Y�3�bv���b=�����k�LTޭ�N�e�v���q�P��}i�cz����E?���R!��˙��:����c�/j��T>�w\�g�Nv���z,�x1_�U�$�x��93j���<���Q|�F�=�b~t�
��ԧH+���9+K[QSP���[$����uU@�xBM��5��8�G����F�c��c�^�
�Gs.�����?��i�E��)�~�vL ?�2�b�H�md/�\�?���m���\�mۛ8�ɮ�*���,���Ұ؛�k���~����������wNp{n�w3|�f��� 3����$��|�c�3Q�Gn�o�6�拧i�ĥ��[X���|Ƌj'�{k�p_+e�YRǠ��#Uj�t+�g�� ��!�Z���?�ȋ��6t�|[i�.Β=�'�tc�e��`c��Ш�	+���'�(�E$����	|�"��1ѡU�d׸��20�����@��Xq]�ʀK�=<�]�~����
�����P2�~���ufv��j[g�ͩt���4�Ç��>������R��Fl٣Tu_�c������ڻ��X���<�ح"�_����]���������ǒ�[����k�Mf���r3ڄ�4x�u�|�Y�.�.���B^�S�q)X�'b�!M���Dy�%5Ŷ��K��jt��� ,��K�:�eJ2Iʴ���a�>URR2{��(��g���(m,a(&�D8�)ءa���:��>��ź3V��c��#�?>� �-k-s�N�;C[8�xr�T�����M���A��5&yL���K��G�Xox�v��-o��K������jO�t*�g�p���O��_S�������:::<�����꛸�ʱ�&���2��_f�l�u���_ǒ
����=��G�����ߣ�{�������%���222s�,kZ�H�t������"�l�"k^���#:>~�����q���¤֮Nm��nS46:��*���a��y �:�/�'�/�N���#c����6uy��u�mQ�Y��yu��|zV����T��Z�d(����'��ڵ!��u�@���Kn׋�{�ɷD��{�ҿ�kǎ{onZ�����M��&&>d����x�����/_o?�KL4]s��p��C�����R�Ro��>�mH�x��%�K��Ĝ[R:+�G+�8p������D�"_Y�?5Wk��|�n�{�R�?f����4�����<���*[�|{46��}S΢(����!/�8<Ǝ�^�t�et�ϗ<=���7`;o�Q��מ�C����F���;+�[|B�uC��͗_.Ƕyl�57{����B���L�%�Zp"����lb�ŷ�O��j��ͷ��~yq=\E�|������ �y� �mז#Sy�E�}#^ܖ����������������lܩz���.����O�ͽ�+�a�����, �+�C[KW���7�;<��FÔ1f�������QQ�M$v����	�>�������@\xL���-q\-������a����id��66�06���bm��p{������"����bwG�<K�X彄>�������R-J��G��}��Lz>������55b؀�RԚ^���y��o���S�����q���^}6[i]^����ReA��'s|����ɰ��R<���Შ�'�6����K�l&�JL�#wE���᳟��l�u���Xm����js�dmjs�H�6���Η&c��]x���)�>G��DE.�;���Kg�m�{�]<��oz��m��ξ���6�|ѵ��}9נCX�	�jy�/���ȳz$�Ó�E�M�N�Ǯֽ%���G:�-�[��f�چ�:�f���1ּ�d�p�s�Hߙ29���yM
�xd�a�և������
�f��R����i)�5e��O���筮?~�K�ɒWf�v�(t��h��~���B�b�ڴ�ˣo�^F9��Ie�U�a�P���f�O�ޓ��s����B#Ǐp��2�s;��Z�P�ֿѲ,j�Ce�B��v/����?��V$�cịG��٣����Q�jT	)�B�lFB�h���������Yv���돿�ܦ�Y ����6���[9xxCS��/�����b׬YS�F[�*�٫���+�{����;����e�P��wY9uΒ2�7A�*Ҹ��޻��7�1(��EzS�]ׁ.���������իW�d�c>��g�����6b��d��Ip�����H�O�%�5��W�zl'5��|�\������VL������UU�����w���#�5��&�y�'Nxo9�� ǩ[/a_<(d2>T�P$j�{{Ǖx���#�Hs����+W˹�+Ə��9c�i[Mf���s
��	���~�5�����
�� o�"�����E�'ؾl�.������R���Y�f��1	�vq�?C��U2��#��)--� =��Ν;�Y;��C����Z����&�,h:�t� ��)���]�#q����
.�� 5�<8�M`�2���6}qM��h��S��#��io��,s��wJJ��D(�yb�I��jW�,�v�b%������n���ج,Z�U�>��s��dq��X7����RXL��������{{{_fr�k �.g*͋"�� 1� �HP߹� �iq��O���5i�w����X���]�-n=1�Q�.�%<��^���9��-\i��`���s��+�>OI>~��Q��[*F�	G�ɭd�)�1h1�Ҋ"F??��8p�T8�/�522�{�W�q(�#���%d5.ݯ�Z��� �3Д�%��W�o�~YN�mxM����IFA/��g׍Zc��9C�MUU(�eI����4�w�����74�M�:Z�-��yj>�Ц**SR��zr�P�YYY\��.��A;�9o�^B��`I]:��B�����6��,8�*).�a���w�0dU�io�R�.������i8Xƹ���/�$%�l[�p�O.��;ٴR��x��U�.���������ȑ���WU��<��]��=�R�;	��~���y����!������'����b��jl��9��~=�LeL4��]c	�m3x��W�������_������7�W����d��e�;R��}9�l���̩�P�\y�j���OsR����~�iQ�}B]Dg�+wHn���\�GV^� 3�Z�$&&��~�U#1j9�nD I�	����fo<-��ʲ�6�psc��T���"7{x��Ea[Nև�E�F���$G�?:UmZq�@ʉ����Ho�3B(��[�p����`��x?.:���-��I))�|���ڝ�`���[��[�Q�C��kp�P���2��s�L;�^����✢�sT�_�^�u�g`8|8t��1�ݻx������;/J�,ů+9��ƒ�G����@LtT���v�����O�:ՉE)�t�b��7!��$և�;3��e-���������̕�KH[���~n�BM
�g���ђ9ja[$z�ԝ��5����tc��b�"`؇)���_9,QPG)v_^4���e]�d�Z��!�m"�3���J�|~��5�rd���͛ ڊ�.��#t�Uh�@6�Y\I��G��~��	��T��Vp4�h�.q��<�!�;.
�Θ����v��]$�޽�����d�A��}�ә2�u#_����b�9r�[d}�[����x�����w�˥���@	;)�P�*��|F]�U��֟]W��9֓s��z&}uڣGE��f
o�1qS�7Ҿ�׷���Y�d��Y����B����冸�ꇾ'��O���\śX�3P �:/���I�Y���WDw�Vh�r�~��$���?��n�]ztt�r�V�@Q��O����Zx%�v�hy��tld0���>`�l���Yk�Ssc�I?ů�T]݋d���ݥjj �A�]X�@�����w��q5�`Mv9p�]�33�*�\�H�/Aɾ�i�HK�w���Q�W���o�r����囶	"���!%�6ߙ2�b�"��~c�!M���|E������$�T���ǅk���u�U�$��EJ+�u꿨�+${��W$�m�)ҿԵ�k���2�����>�����ZB��+�zs�����|Oh�������u����,��:%�)Cx@r������P%�����^9�@D�Z�e�Iܐ��f�O`Ɲ�im �|�8��ڲY��	a��\o�`%np��Ngl�����Z�c�Upi�uX��,�e9��DG�	M$y���ް��L���Mݶ����ї��� F}��yP���`3ν�"|xnC�Umֶ��"r�g+6pE>���]2�J�m�2Rn�,��nwڌ�ٰ���F������\q�G�8,%�'��R�K�s�S�}�%[N��T%Wey4�	�2Oϥ^��c2b*�Pu^��z)��������o�ws�d��3���b)UJ���1�[ȍ6�t(��t3,z�nܸ1���i1u�F8�:�yv�+=EDC���~���;l�4�(�u�����d\>��odĢ��v�ȴ}�>���rS�=����UL�'�<F��
�M̩*��&��+9|}� s�����OK+**
��5V�]m���P�8�v�Ѫ��z�o���lƌ� m�ュ	���'O6x����*_���X��_o4:S�����&-��D�6����a[�!|�f�%�)Q&�ɖk�LME� �೟D���/�a�?���~2�1W:��@�AD(�\�)[Лze�L�hm�p��,�ϳ�`�鹪���V����.>|z[N߇�l��a�����=������BB`�>�N�j߽�A�i���1JD�ʄ���g��Ĕ.� |U(�?PX��>��6 T2̩F���'s��v�<S�AXR�;8�m��D<��R����MN���2sa,=j&�0�����Ms�e��]�^����k�n /o���M�+������%��#��veu�c�C��Aa��x`�\x�����9C�D8�h�|8I�t|lXb9�DŦ �EnYY �v���jӍH��c"�'��)�>ʸ�!a<�2[n�1����4X,*ʐ<��t��lf�
2���"?qQ��t�pZ̟7A��jn#�<t��T�OL�0wO����]�vj���GrR��3�	����o�hFC`�����z��{r�*S���[�v4�e�IN�B�������-	,pd�kid$,�,�@m^����G�����F<�
�ioM{Ld�L0+�����N�T�|R�B��o�z����3���+p����\A��]%�fV���<X2��i�f�s�����r��r��O���^F�E��J��R��\�a-���t��iR_�ۗ��P�ܼ�T��w��G, �[�x���� |3�������Ye��
�Դe�T���؉� ��SW���Jcm�z�+«���%�}`�w�o�����n�/��4�g�qiR���R��)�`��a |\x���|�>_DkN�a+ɴ9/��c̆z�[Ճ}*�8�+h�P6�]���ti<�jrsU(US6�Z�&��������"RS��Q�^^�)�Ie����Ç�xC���J�i��)�X�۲e�j���|�Z���t����70���:u5r�| �{��P��[)i�CW$^7�r)�JT�:;r,�{ QOR���G���JΚ"`�r199�L�m8�9ɵ���%�đ��}q�;=G��WB8>]�����^N���D�����2������|�$�h<��VV�ڠ��j4
�	�U�_�P ��Mm𹮞d��O2${B�;?�,/�+o%�xgsԬLM���"���.��ʿ�F���U���FW�f~�C�#��'���Γ�t��G��Q�S�S�c�	[pF}�����p�3_�L#�M���m8A�����Y̓h�`![6o��/]����=l�����d�w��UZT����Z��â{ ��қS�����T���ܽ�E�>����|(WPWY�.�>o:[c����24�=U%�+�s���{?md��B�����+~�� �;Ý��������O��9���}����Qm~��ܫ��M��[��N�hq��)z�2�oYÜ4�b���q���M�3�e
_C��q�
�����m<�6��j��'If���sd`����y��;M�;}:?8bb��)-V�z�@>����j,F��p?��f,;����O�ggc�n<}�d�W�6[@�ي�9ΎK,�����[�pY�``�����U^�:ZÐv���V�}o�W�k��Wz��ύ^�J;<��ю)O~W��V���oGſ��2�vxi�`�g�qR��#1G���q�Y!��nU�s}{Y��'N�Г�|s&UJ�Er�Ʃ��t]���/^��C�\�����/_�L=��x��:N~: G���p�HR�n�/��8���f0$v��.ڑ���߮fn��-\cDV{<%Յ�=oo�B*�`7n_��~�Z����N���|�L����3L����4��&P�Ǡ:_��Π���'Ԛ��x���P���81�wI�ا[tP#�nrEtL��̖-[؂���1�2�:�W�= s�3#��a柟��__�>,�p�M�Io�����V�:����
!ˡ5�v2&g�އ-X"��� �n �CO$*�ɂ�Ӥ!��^�or��0�|�ɴ�m~T{���M���pz�F�^k����w��0��W�
�im2�$�&��X�i�eO}H�erv��Z����H���ß�\���]y�T��=����W{����ݖ��,`�=��^��S���&��s���Oy�9F4����D(��]o�
�>�,:''� ���Y�^wN�3q|���bR�b��$�T~|Ԁ<����7�y}{�P���Zw�q�S]cj�uWf����܌�*�c6���f��j{x��gW�A�8wQJ�O�Iyy����j|.�w|�`��Zr��3`���7s¢�{�3v��+�Se��X���MLdHn~&�H�]&���9��#�U�7�<[|1Pp��0 �v�e��p�?q%M�/2�&f�.�����A����K�?4���p��Ƒ�UjiiE�� ��8A����=�uj�/�.�3�Fr_�W�cn?��>������3���=��J�T��Ӈ8I6콬m}�,���/k�Ê1;�:i�ĩ�l��@9xٷ�t�3m5� f���#dS��2LN"��t�d3J�C���F�zyc=��3Dp���E�(R=�[3XYG�����:���4[�[�"�?4�K�$Q�D@���?�S�����19���Ƙw)�w�6o�9Ɖ�IȒMd�Ԅ{��~�.N���ƨ0��m�}S3l���.bƅ=<q�f��װ:��P'���%�u��un��U}b��p+CҼ9�v������-��㏟95��VVi� �?B,R���ST��� ۮ����-t?��7h�#��L����D�Ϟ��U�e�vn}X	`��m1����O�*G__c��z��l�-��A�t��6�\�YX�]�|9T�ݍ/_?�Q� ^TT���o4�"���@>ѩ�6�O�ۗ�����Jy���MA�0�yӵ�3Jö��PB�
ޖ]?����C��*"��-��BU��$r◒ζe6�6��a�f��$G�.�	)i�����M��IuX��,}�ǕfiZ������3�-)���oiF|鳲n}��,���r&7׹_��l�¼p�e�1��߃T��P��Y���G�VP���	�����̩��C�]]]XY�ooH�L����WP�=RtUT��+pΜ���4�v��^=hb"�DI���=�:���>�.�)�V���K�*��ݻ���sd�ZH���6�-A��|�2�k��:�������=�\Cތ�Q���ڶd�x}�A�l:]*#����zk��X��z�d�\0� <b�1�G'\~�����c3�΂�-'M����	�#��:�����Y�"��0�Y��bY}l܉� ��?�2���{W3����k�c9R�***��Ǯ�S#ws/�
,dI������iE7�E�I�L{�k�D�}Gg��4 ���������6y��6o�leGv�Y���6��6>�I& �m�
ˡ���w�<���A��Xg���~1R����1X{QԶ���:���v�Z�P�X�ϫE9�Gߢ��c�� 1�N�����������Sl���H<lm![1_�{������^��;|8�0�&$O�cS���9ͱMкYKF��h^_g�D��L�"��������d;�z�E�$5P�1E�u�຾�A�w��WD#�����Տsu#U�Sv. m���a��a�r��*�r��Œ��2��za=[�=Q#�>���t�T�#ۆ�[5�1	�:���{C7.cj�Od����V�{��5w�T�>U�/���w���˦9�,�x?�i�<	��#�]�����wYQ�%;`;��n�K0� �&NT���b6D�ЫA�혿J����*�{{�R��`d\���X,:��l�����.�Cv M�ۙ'S�&N��HƮ�^j�����a�c4��ML�J+�� �7��h
H�漿�^�j��
}UfX"cnb1y��t�y��=uQ74���O0p�8�_ȫH�p}z�&p�C�G^�5���ӛ��4̋�-+^�lz�MЍT�y�P]7�)L����}|������7�<.��ݺ�C���j���Mvg�b���#�;<�|�%�b�{Ř���E[�|@�+��1Z���1[��o"�!
b��蕔�n(���&�����g3��q<8���!�,o�u|RKU�3TΣ���29�̸��J-4���P�t� �ʃ�-��D�g��<o8?qPh����֛h�B: �y���,�{���BU]��-\ЉS8��[:O�0�K�.&���5yV�d4G����_o�I����eUlq	 <`V,��ד]
3Tt[�~6۶��HT�d�>2��.��؉�t�J�>_���8��� E�.z6W$�zS�H"����k�ǭK�>g�>��"�u+B��\xm�&�?�����ɘ���@��Vn<��|��!rd�W`ح���sEF�&�8�kcI �όo��ZJ�`S��k�uk�OMmZE�r�������tص��v^�-�����{�ZӚ�У\���N��BE{G����V9��	�Yfx��)e0�o#�6g1�ߠM��{ x���]��ͻ�d���^��zRGA�V�{=��.X��Yi$�t�{�5�[Fj���:�m#h��JW �a��;q�����ı��ƶX<ޑ�y����G��4,�����P���P�c�ַ�H���iR�nx�S��_��n��>H{�מ����o�Vݝ��e*���ۆB��+��Ԁ�c ՀdW��H�;3w���9�σ%�1Q%N;c��K��ց�Z�5���A��?���q(G�)����@����}��b=�c'%���� j�s�4�Es�J6��s��@c��@�w-�w&	kʺj�I�;�N ���9~�����}����3���|<�~$�C�k���1�v\.��lM����]��!��ӴH�W��<`袼�6Q�W����G�����G>�e,Ĵ8���>%qqq�C���pv�tG:!�Q�I��C���h�`�%��MC�:02V1�k�@�����g.\Wu��(|Zκi�{�+�`c�45�`�C��O��E%Yg�����8�Ĳ����ö��ࠠ߹��Rn�Ȗ-[lA��<J-M.�6�y����;�®//�):�� ��07^'�0&Uf�WO��g���V�Ȕ���\i�{�>�fa�D���0���|2[u��"���W�X��D�w��)l��"���[��>�k&&�<k�$�3Ʒ�Z���d��Zr|�B�b�1�&�iY���7�;SF #�={��bs"HP���Tx�'O��e3j�6\�}4������Q��$]�Oɠ �>�;�xb���ٚ��U��#]��`!x������w�ߧ�&8ݎ�]��[����j�r!�'�L���d��<��&�{˃�R 3o�n1�)"�CυHU1��CĠ�&�閃�s�o�W���~�Nk�a5�>����C���[���/g��g�v@=b�=��}-\i�K�U-�:�-�6���a֒����p\!u4#T��=tp����U�߈Bϴ~��<�#oTj�����Q�ݻk���!:�;J1�b|N�\w�=V=u���W��J�7f�%7�iy/7��MPŹϷ6׹���� [�X�$�DW�s�E
��i3�~{ve�.��.�%��&���PU)�
c�m5�x�d�> ��X�]g�-X{� �̊�>+�����s-�1�׺u��k��p��A��n�q��Σe��!"����fO/M����ĊiʀD5S%�I��D�z�}K�Y���J֖�w�h��ů�u��t�(c��%�,��r~4��&�pB�t����%;��FJ`z QsF�p��K�ɇ|a�mYߣ]��:��FV��W/_���u�o��&���0Wn���'N�X�<��0.-m���zo���g���멏_?�<v������� ��k
XE�}����f+w<�J�j����>�ݜ�s��R9�����	Jz���@��P2�Be��l{�o2ʸ9qlt8��t���(�� ..j��b�c�f�}�,�����&9����C���t�s�A-���Ũۚ&c���bz,LF�����4��!ʒ�+Pgȓ{Y��0�Wi�|
�{�L�� ��ś�wv��B����ȅ���}D7�o��.��Cs���]���B�b́5��l<%ι��v�5}W�ŧzE�ZB����E�X���N����.w��cW07�ees���a�h�A�	��ۜS�F�� ��\� +�Z����	&v�'�[�����{ �o�\+G�4qw�g(��a�K��f�j]��&��@ȥ�95,,�;]�f�N��5t����3^�ǹ���� �<���>]؎OOd�4�a��s+=����&���bl1��I��bl��_c�u�8��N�����ʀ��D���6�W@v>�)S@8�y��+-�<Ob]������O=z,���!�c�
�ts��8�[F�^�e�����TE���Զ�T��A�V�/�Zo���Gr�9��z�8;(�4���}���7cߺ���;��W{qEEQE�y�춬�i�i�G_2���}E��*g7Rc^=VƉx@`����f&X��<'�r8��ƾ�u0���}������ �e���w\!
��[�[k�l0ғ|$��
�ۆ�Z�����D=�����eO���j�Y[k����.�x�2�E6ax�8	�
�EV��X+Rh@���_U�uZ��"Ѥ�� ���S:�Os�iF0+�
���sT���U`��kR�C>V���su�*�a�(��t��T�qI{��o�|,c��M��zy�j�;v��=w��m�s)�53���<���%,�ؐ7PO����~t*Ƭ؏-�����������A�l��l/uc��	sQ�?6�Tv�7� ��7"'�����8����݇�FF�F���]�k�pѥ��XʌE1��ka�)�n �#
S\��o��/��a]�r��l���@�y���/M^���Df�$C���޻�����ŋ�1O�%(Y�� :;�$��cV!-��h�)98> �p�&&�6���r�w�w�{_\6�El�,I9��)�X1H�W�c��U�^�M�4ԡ��n�S����Hw7�ś�����_���P��[�E����m��f����ؼƽ��L�>�V9��-�K�/�o�:�e4]ATp<�����(��7ZK޺���ۍ=�2@������D"��=-w9�ME@�'�$�0:ŋ�I�s."�Q�]
�~~*Rܡj����D�jN7�'�u8�n*��i� p!�7 �/Ĺzx�So6U!,��4m�'�b$FK"�����ǎ|��/�(�	a�h��ݳ9pf�8��B�q-Q�8�XT�� ��yz��
�&Z��륌.5�&�B�j�M`���Akj��^z��!4���$Z1k�Vi{Cg�v�U�b�<h�-�o��`�@�~^�u��TmG���ǜ����pA[V�;^� p�����NT�aj깃p����U�	w�`�]|���k������d~�f9�� ����W��#�>�I�{FS������ ���(J�)w��IL�f1��?,"l|�:8~�&�^�r��(�"OZ�t�6	�>䁭�xM"b�r�r�{F&a� �`H|q��g��{�M���h{x�uC�R_�Sq�C�l����cl��`a��Â����l��SSO ��l(.ޚ?����h?l�B1�㚹��v:�A�m
��[	$ߝD�dC��Dب?>�L�Jd�f��  t�\�k<�K�tO���+�Y��nwiR��.��״2�cѶi������A��oQZ��4�%*4�Vy����1�)���XÊ�8���D`�Z�%yk�Br¢:��LQ�9:ܯ�R�;������_�2Ɔ�� 4`�{�Ú1��>8m[,0��$'��q�>����_֬��b)K�Lth��O�V�ÏA7��]����eM��b��h4Nl��j���1G,�kO��<���^Mf�~��f��x�QV�΋��è�2Lp�|0J��EiWt6c����|��R]֛$�BX����u�������bu|�M�"�ɻFK���%^� ���%��j`�g�6��7G]�Ǳ��r��lq�^�CƼ���Y�0'M'�&pװ�9�5��`j��&c9xBv���sj��W�5^pg;�Y�@Ҹę�k��;���g������0A'v涻�X����J7�����b
���� �4���%�}9B��آnY B�2��k�Y_�vk��L����*�H�]�3[���1��3�P���Y~�(�(�}����և��k�601�Sc�YN�T���*4K�輈���H�|7��F{O�S�k)ݐ �=�z� Hp�:A
�NY	��m#���~x_=��L�����4����蟃����1&�n��q=2f�Ó��3>_Vh���'��".I�e��r�h�[�=�]Z�-!rI�@��=��Ӥ1P���xB�IS-��-G?�H�$�b�
����Jo��Bg��*�E�������C��⠕S@a �_���	����Pv�ƍ"��D'!l�ZD�%)�)ih�M��2��������+�3���H��1��_�Ҥ,X�����au;nE��{��#N;3��?�Wm�`��o<ag.�P^���i���F�S�5aIɇ���:/1���?�v�y.渮]�Ko�W̱����znn
���7�]V�q�G׉�h�6��	��U�.^�w=k�'	2y���ݽj������h��
S��i�ر���xClO�x<�)w�,@��{��Zf�ڵ��_��KU��E�wma2 ݥE��� �XԪq?%E6���^�lǌ1��X!�BETK>�Rj``���P����7�Nd��R5	\ޘ�y������(�@� ���q�;}�0s�痗!ŀH�hq���uX��}3s�ӟ �����~x��x���L�xo젆F!P+��VZ~C�d	U���*b��>2+K�s���ǚut�c��
+������|�qT�X�2U`���s�'�|-Z �닷Y�j������f�&��A��G��������	Ѓa��ξ�����W|¸�#�#��}!�˗�$�[g��?��Fn�ņ���v���*S��XD3���(+������7��F���$��"��+8��B߄E0���Ǭ��5�Mv���=�+bv�+|�6m�J)��r��|{'�.��`�a������bUG�ũ��A�5�b��S���i{���b�<H[e�q�*f�Q���j��Om��L��^��ВZ��� z}}}���t��X�l9(�^������Jpz[�u��;� �@p%���N�����_"6�W�>��:�Cf�~��/��8���t8ao��h�8��HX��ԇ4dF��=�פ�����o� ��z�G;�X��/�)j�V;[�tU���Y4����Q1a�0����R�����lmFc��i�뭺� .v�bO@~[���h��Zѩ�r$6��UBX���̘P������ԠHh�$U`X�	�F>�?OX�nN�2f5pb�����7E,"�s��b��^]w�����<�Eޝ�z"`6�q���	e ׃I?2�X؆��j#��ǋ0'z�7[�7d�������ʖ�;�MՒv]�'i3���җ����`�9#@� �-���b�9��j�*�F�\�psB��V�s[&Z_����YY�9O�"�K�pp', �Pt	�zE1V�M�$6iAl2�B?/�6�D���GC�8%7�بRi'j�JW�)�TrlF؁��^�~H���M)�W�|2f�ʔ����l�f������G��f-ڸ*pٙ]/�2$1�D��N%��_�_��`#K�6'�,�.b�	ND{����XN���M꫻�ڡ �f�!�v�������
��h�Z�������Dw�
IԈԆ����`��`S����:,���?�=��/_����+n$�{���Ue��3lp�6&JϏ/lb9exS�L6��x�Iked��N�,U���2�."�^G��f��xpCW��F<J7d�Q�[HS*�Q6qD�b�O�Y�f��+��K4���Ө*~�Z�nb=޳�
�?U��*Vk�
%q�;�X���Z���B��_��@�LT^� ��%�1?f,�Sr�t����T��Jj �SP+��B�y;����Ǐ�(�<��6-�>n����G =,j{"T��R�~�m�p�F[��rH�E	,���[�u�R�H���'F�ݫx54��M���#ɺ�K/���C��=8KBU�,]S�����q���M������� �͚����g��[0,�+ N�@�G�u��.�K����K��]���N#�h"P�듮�J~��=�|U��h��@�?#���tɈO/d�_�Nt��n�8��x���$���\�[h)R@
�S��f��>p%5/sJޫ�8259�
cz(o$*����Bԕ2R�0<�2�-�	!�~�J�	���ن%Q����)�8��T��`=��>y��{�v<�	Gs���J!Q��m�$�m� ~�K�n��N����a=�
��Y�Z���|d� w`:�H���oG��Ó{W,�նP�D�#��
����IVt��b�ř��~{K� UO��V؝9����ޒ���c��x��:P��5�sޯ�I3ftyc�b�͘śn��������ё&5]V�$��1���y#����U���H
ܲ�,;,��������u�GG]ք�x+J���5(�o�<Rlr������c�eMm{�ݞN[vr��[05��=����Ʌ)����'&���x��:X�%��1��,b���Vp+�<�f|���@g��맦�ս�T}<�mz.�H�x�"Q�F�4�������r^<���jZX��`�BR�i��6b�ż$����8�@���`���_^�`kJ��7qs�W>0�G������T��P������/!������'ʳ�U��Pb���@�S����8�57~������xz�]!NWߎ�°��;QO�>^�[i"sǧ��͗qߞ��R ���'�E|	�����l S<&Ft#A��s?�����ӓ��m?x�a�A8���̛C�CZ�|9��,���!����䩕�܉Г�3Xq��dN�m�˫��-0$2O궝w��Gs���[D	�|�(cG'���v�N�C���8Vf�A*��0&tj�u*?����ćO_�?�;�c���ly��K^��R{���V�o3
�h~���U�h�|:�f�/�ɴG�D�"LP�?��cST���)�iUVV6� k��7(sT�u�u��DWɲ�5��_�G/	#|�_�DՌ��/�#��%���>+�8<J	dy)���oK�o�����;(eC7�����o�3M"|��-���%��'{�Iku:.z���5f���M�ue���{�m��"O�=�>>���t�Pe�Xq]�:�I��\��T��gO�%�gtfx�����)ʧn�_����W�!t톛^�^�k|<=��*n��컱zt8&X߁���fi���/[$��o�\�^��}�e�U�\���X�ʤt,)<s�� !�e��x�����#ɑ���&B�v�a0a���}dOR�>R'�^��O�Y�	m����v:�N(���6&tj���!��2�'OR�/��g8�������K��s ��I��Qt�'�_�
7���vK�y��pC��o�{YD�:��"D-h�I�/a�vHз�է ,�
Z����u�ZB�e�>\�M�� l`�%�қ~�~��7!-�mt��S�i�r��Nq�[E��LK��:���������-��	x����0�{�I Q�/��a��W��� ��c�cAm�I~�m�xLR�x��aS����>f'�Kn���� %�5)Z�֐}�b�Q���>'0+�Õ5��>D	՚�&����уs �
Re�Xt71��1�6�}�=g�=��G���T^v�}�dF2V�l�_}���pE1��?,Jo=F?ٸ<բ��m�.�"i۾-��=���ʗ�f.\G�} ym��a�xj}T�溫e�پ ��N�����s����{��q�v`���K���q�kPia�REE�}�b� �v�����C��\�޾K�սT���#�[f;�0���+��H������
�t��_�ä9��և2��D�V<����V��^w�$��z�wuӬWf�L��nb� ���N����+5�ʒs��b�]*f}t-��a�s{�#Yy'5��:�����5k��`��	 UG9��c�������]�m��vb2�v~��u����)��`0~�A�;�L+&�Ff>- p؂R�
7�6;�}�̢�"ؕ��o����"�}]X��R�=���_EO���#bgq���-P"���𓿖�;[��Q�$i�u\�8Go
�ϓ��A�h��k9>V�J7w��Q�e�Y���C'���c���R�v��t�y睝�ĨR�$k 'h����B2���}�y�<�F�ңJfa2w;G�Yݰ���c�F�:���ɹ������X�K�~��Q�#u�0<s�t�L�����Q1��|)�lo�>��&uti����=�HL�*Z��鉓��r�<g�\)�L�g��#�6��y+ή)�^(�Do7�,bs���d%/JL��X����߼wrrj�n/$~�G�˷s0E���hWD�=�_���Ţ���q�b"'>]Ѷ���xz�n�u�9�E��q��!S�>�{A�8\�L��r&���F�+�)-�G��唓&ӢY4�kۼ$׼���B�H��J|+�a�ҋi��І�����m��R�#|��eJ�2��.��ӥ�Ɓ��$�����/���X�H���'#�a4.�c&a��?_GF��|��ܔ{g?|x��%g�DV��d����B��&��`�XI�����*�|���к��V�b��W_+�M Z��ް���&vZ���-�! '!������&L~�j�vbe)�E/�h����&P�����\?��p�$Ґ<2�A�P����`ڈ���|��v#++�l�խ�$�4rǆ�%,X �g>�:<xP���%y�����Lp��wB��%jn.D���yP�B��������������@9,/��;s�fkw@}��_Iq���J8$b�ƾ߈��8�'����wP_9]/�-y� �y��er�c?�<�3AmT��OcJ�k��.)[�d�|��TìH�����y�������C�T��Q�*Y�r�m<Q��wR�p�DU���=V�i���ϊ���
a�,�#ȰT�9V�0�NIz�`	��n,��"{��T8a�@ بz����m���%�v_�5��V�2M�������R�(�r��O9%^�<��(��HV�F5�|�u�.#���'���|��|C2���8l�I8w.֓b���)<b�X�Q��e�$k):rRKUEI���lJ�A�8NԄV�����Z ��p�#B����F����ʋ�Ұ�Q8m��?��p"���RopZPhA�a�p�����==�������(�cw�9U/���(���A��Qo�S(/�2��!���s}-g�qۃ�V<_y����y�����6C�%xb6U��u`����%��D̈����e��
x֦�C�\6�=�e/�o�'��2pN�+�bP���1�[�w��c)P�ȹ��f�� [��q��dC�=g�t�ﷷ		K`|,�Rg�_&M1nM��I�3��A�_���ڏ8M�N��e������(�8��Ƣ�H�1D���+v}�6��x�\�@8��B��;t��n�RLf�"�/(v0��W�����T=���GN$�4�E�V4��ߠ�6B�*��!����_Ýޘ	
Na�1��^��Ҍx���)�@������J1t�iL)u�*��x�yǎ�oY��a%z@�ÄP,�w�nX����j	������TQO�*R:�����.C8�dE�>ߨၖr|iBgڃv�'bӭǈ�v�A�U�o��r�궦׹a�fv��JM�+1�ȝ�����J �K�:��$k��ڀY����/q�x~���\�/�x��R���͂���`*`K��,L��U�x<�p�V$ 8o�2tuX�n��������?�V.y�*|���u ��,�x]�0��ܖi���A�_�n�{�����N��hF��>�}��j^]]]\iŭL7H̛����� �Mr%���-ė�}x-_�&^)'�o%�C���9թ�q\��K�>|���T���^�>�+�q�����^��J�>:T���VR�?Iq�3�Kir\Q� (�s���*O�A��#��q��J��%����صPu�8�m�arhu �����4j����QA�a�f��HwN犬�����h8Nꪫ�{��-��([w�Nt��F��U�S�cltC�H-&�\����+�[==Q 薂XA#�DY�9�+���Mxq,}��&T�nh*O/.r��Dn��=�߻ZP���h���+�_=�4����el;f���ž]`n�t�Lbl#��}x��g8�Q�+N?&��� ��-Ҽ����E8�3Z����T=i���#���8���L�I){W�)Qd����(Z�ӂ�g�MSn*�B��Wv*%�U�e��\����'���?���嗙���|<�����<�<f��f� �]�&?���q�%S�!�������ΛW6QO�}�d�زH�.0	}]v>J�����8K�37>5���d���6-Xj��U���bR ��b;�<��{�GZŦW���Ͷ�7��S���� ��I�t<��.��Kc�Ѷ��b,n!O��`%2�w���թ�s�/�Q�xp2����v2� �?R�w��y�3Z�Y%^q���Y�HM-Xq���,}"ݎ��{�s����0XM��C�!��K�@_���&�=���E�vy�q ��P�r
?v��̸���F�ȟ���f���lN:��x��l��2�0�r?���c|�g^��H�aJ�f(�����yO#�#N�OO��tƺS۬�;��챸t � &��ͳ��j�a������7K͐�l�j�c/X2��/^̧�\2�+H�KD��`�O掫����`��V�K�L|�P�5�h��svg���M��vh!��f���#�H=�w��a&k=�|�1XG�W�v\�f�.��M��S����\݄iH�kx�C&fN��ag�3�l9�x�l3��E"ny]%&��������-�B��X���꩏1�0��a���n��L�l��/�1���cS�M~��V��F�:�"�(�$����K̛{�:�r���7��\�z�bti)�|��&0��ܮb)�L����P�4�����1�WW���d��l�?���,�H%%&��*yx��v\��`��Wgv?#�Ջ����O�U�����jt�c��u�w($ke1�T�-=�i����?1]=۹�6ż�"���&31{��'Z�/5*��H�{#��8����C������v��1k�0��,�{�!kߜOvN'�;}��Gd�<�ۙ���kP+[�=�/�}�w�Ԗ{��L���r`!r�o�aal��e)z��a��~{N�:/p[G�uҗ|P���j����Ǒ��b&<Y��IW��Ӓ��7�N���ra��wb�`���%��a�����
��������x��6�r-���-����	@z]!�x��g���V,���M^ï=z��J��x��L_�	� 8���ݱwVl/f �O}���8�{���F@k�ٛ��=�7��n��������U�6� 30'��u2#=��~2��7ؙ#޾�>��C�퀱d���u\����CR�Sl�c�8�X��W�\��y$Lm�^҆�m��֣R�&p�����y{�Uuw�޽o"l��#��|���E�����0�g�M�Q,d���<��z "CL�%������t��f#�gl�G�k|���a���]��G(-�+�wjls�?Z暻�.o�e�,�½@"��D���1=�di�����>Ea�SX+�I���l	~SoU�P�:U�!�}-v��/>Q3���M��}�(�V�#���W��9���U�ܮ)���i��A]05Z�Yˍ[v,����W[4����^#5C��-�̪#���L�a��϶Y56�?�$G�D�������ia��Aof��eBd�ݠ[�ؘ#�?�b����A.X�����I_ͩ������xt�D��`�R�x[t0�`����L�������vWr�ҥ�1݄���=O��1a.���R�.8�r$-3S{]c*�nlп� "��qz��'�ߵ���ȉ�Հ/n(F5���\�%��yO���3�J�s!��V��Z�X�ا��2��E�f0>i/FgZ͸�,eK&�bo�60g�zk^�I�(k�cX!ע�I�°�誦�Yal��<T�z6���}ŇU3 �;g�q��X� ��8�}2�� 9� X$kK����&,�=���u�!�Y�ݬ���w�Zg�C;Z�d�5��:knCnŐ�l�-���E�d���#�ؑ��Q�O���/a�xڊW`I�Ԁ�yk��k�twg*�̨�m-����/d9��ꌜ�����@�E�Ы�.4X���n���?|�/��������[YYڿ����x.`�{��a�]�4
��!;��V�;���jo~���yyyy�D���&�jtY���u�<����`��:a�lX��ˮ4ļ�:���O�#��y�:;G=�QǤa���`?;�����V,C�T_2}%�x�Ҍ%/�v�Y�7P��A-���TGZ'WU�9�=^ٙ�ob~��>DI6��}Q@ݜd�7���}��p$���n}?��J�����T�xӦM��D^z�p�^��Y��ꄽ'���U�>�}���#�Y5��0��Ě��(���W�Gٟ0��� }i��`�+Ϟ}P�o�7T��%�����V�i�^�^�p�>�w����>��$,((h&e�f=\	�w*v����C���Ξ={�iȫ��rn+nH�_�r�ɳ�����	�iŝ��ET �QX��������!�i?S̿k8O�ĉ�ؗ�|�l��}���_������}u�a�E,v,y{Wk��ϫ+6y�fr7O�s��wS/��uUۂ���d�[��N��?�L {��:�0ky�{T��@y ��?���O���l}$^��:+�ݱ�i��Vɖ<Lʟ���1��d�w!dy�W�`�v�W�eox� ����C�ox�y�v�Y�s��;������W�M�@0,*H���)��蹭�s�@ueX:j�|���S���ѵ�-1�+��[B�] ��hS�@�s�C�x[V�`�@�wR��
����f��!Dn���:;w��i~�'�UOtŀJ&�zcg�C���S����([�xk�:D���pP^;��mX�.)}��9� xO��� �)�t®}`��� 	�o_���Vt��D�����d�7����>JC�̴iK��%s��`�It����� l�EZ�u�9`1�
�	��k�PG'��z�"/�^���$E�ca�Y�1�;`{Ĩ^�E����ֶ������f����[A��C�o}��Q�_<��}8#�?�^��U�;��o��x�>��M��v3-2��R��=�r��?�㶏(�{���s���$�0����}́8�l���Z��|��8j���Z�sη�v������B��,�m�=��z�lt�����G�^6d�6kx��YY�	�Y����Tj��D�/7#F��U��N|Λ4x���`�REY�ʀ��5�ZNO��6� �~I&�x��iܼ
�X��k����X��je2>Sm�O���:����?�r�%���/�!�̋��>��#VVV`k 2�@w֏bA��B��>9��[�U�tb~y�g�+xD�b��jߌ$&�OO��g��B���F�FX�-��	9+v%�$��Gtz�e|�I����C�M#��5�W]�ױ�������Q
�i�E~���R�a��sm�����t:�>�<�[���u=9��*�cmI<,ƛA���d�M|T�|���7͇����u4=X�p�zlE���r����΋������u�5�O�bhLa�ś����c�U� ��yQ� q^�Av��(�"�U�N��[=���Za
ɥS%G�=���踯#ܖ������N��Gβ��������I��7���Z��dѭu��n��Fkk��I=�k*�ZBuul�>�-��?�?&`�
��n,�>VGlא\o�;i��l��R�	�ǙZʨ�x�N6�����@DOBT�WH���aC<|��MXVl
 (<���s<�]U��Q�+^%i���߅�����'i�o�.���KHH�8ΰ�T&��0�E͸�ll��Т��cAicN�F<����h���e�MͰ�;,�>]��	m�)����c?>l2M��Ɗ����ck�����$$x�8��;x��ql�]�]`�i��_.�Ī:G���.�}�dK��7]3����~�`cղ0��â���b��UsN/�A��{��c������$��^��<��qo{��N�/�	myB�_�+��Ri�g��B@���+�nA�L�������k�)�A�	�5���uZx%�o�q�=FWbbb�d��69~�O�Ѡh�F`�D��b���@�/"��K~�!V.��B��G<���+�BgF�S�b�럨?|�@���O�9��$O��ɯ)�ȍG��k
��J�L�Xqs�� �t9��޳�Ռ0��`'����-W���d29~]y��E��ז`ٱ:�L���Ǟ�X6Ӝ�.����̄q����Q���yl�gz��n[1`g�؊7�K�cĔٕD�������w��G5�I�'�p���+z��ܶ��=���nW�������I�6��N�����Βv^d���������_>k�6���p��4����to��L�Y��"䵖΋~����>S�A؇4.�� 6�$�F���>0����{�,���^F����i��U�Xe���WW����ZyRހrW�ҿh�[�I�c�%���g�A�P?��:oj��t!����>�٫�6� �_j>~E[�G:$Q/�Zk��p^䎍-0iǊ��JP�^.d'&����h!0T~X��T���h�>D�����w��I�/ބ����o��5��5�3�M�[�F�Z[�;,�P��LĂ�p�����E)�Q�I_t��7�߰T*��yK�Xr�F���L�[g��J�e;PfZ)�B6��
�拼��h�a���<e֬��Ơ�������^x�N�d����t�����q�S&�6���}�"̨�8�B\o��+��>�#Eu�`i<�&}��=��`�N����J��E5�\3@Ǔ���)�ȉxS &+�����7�"Vk�W�����V�f��+����0�ŷ����!�ƪ9<l�$��Q�)5�j�q� L^�̻�qF����ۊg���E�+�N84��������5�(zL����sn!"ZNO.ԙ�$y,;��4��d�9�~AV��_};1:@6)�� �<�.:^Z;U������E�y�1��$�����M(ƱƧ���'���ܝ���7���7�b��
D����`Ðw}y��]}���0-y� >��D� Y_�Zj��=�4��v<���Au5:�3A/� ��j��E-}�����zߣ{_�.�L�OAL�}���gΜў��y@��(��<�y�C��ςź�	����Bx��L���Hly�R �����5渑@s���w�ז�!�%��Qύy$y��*��{���a���H���R!�Gek�lj����
Dy�k�W��8��(�1
���wɮ�K�g��e��E�48AMr�p�w"j��2�����ǒ��$ZJ*Enl:p� �&^���Ps��;����ţ�CG�Y_ԭ���׋���oR���<Ȟ�c	/`�?�Gg�D�k��o߾a�Q�?�b*�Z��#��ի3% o/}��̴��'Fd�"`�G{���
@��(++[��f]�.)�Q
;���Cş<`�.����L_��]tم�Gಓ�Jj!�1�ؿ?^J��v���C��O�gܗ �L]�sU�o��9D��޽@G��h����������O��gz;�b���㗗
�4->�mJ]6\����N��>=����o. ��E.��DX������x^��"EbO�%�U�W�:����R����c�A�KXK����0,�&-�����s�^}���FĂm�Y�DP��$�X�Wm~0��� �1l���/�h�G�������F@}�^[v����.Z�O/��-S�.d���~�8٬�����<�䓯o�v^�	��!u�|�?<��a�x)y�z�J��Z�g�7��?�c[#�΍�q����&���S��p�6��s�4�������A�R�<Ӱ(s����_v���a&�Y��i���<y�y�h�Λ���W�}��W�ϓj��voY���9�	|b��vm��M����7*�T�Un��I����jk6�֔���S������1�h	��Do}�&�݄�T�M'���jZ?��P�s��\U�.�&������pjpm���x�/8���俇�@�l�����7��j��%��`\�y_厃˰!:�x�E�����Aؘ����~�Ov���%�Ԉ����0�yͯ�(����S�} Cv䪃o�
�̈́K�b@V�c�����Ѻ��/'�Is/�XT �,Ƌ;//Y}K1�"ę�ޒ�Oy���+�������SW�w˅��k+��u�� 饢�#��C�X���ټd�K��O��~!o0����z:*+0�FC�}-y�ݯW?h+u�ÿO�{�f��:�b��O T�ٽ/���Ubg�%��rF�3x ��(Xd1�x'+!T�zc~"��\�M���a^�E����н"�HV�yvDŦ��/���x�u���7o�=�d���Q�5>����_?�����S�Ɗ���zȝ9`te L�=�m�1����nX�9�=`� Y����5���o����N���=^��D��A���Z�Pa]�fJ^{[k�G��Ï����{t��@�狧Q�_\~g����*W�G/�+������͠d����7X�u�,l��!�͵1�=�X��8��;=`DNaS��|���C�`H_�Suu!��S�}k��rj���{3@b� =� ^��vc���w[�*e�����"����i�E���߯���V�|6l�L|����k-�^��}&��Z������+�hr�0s]���{rl7���ly��q�'|���yo��>Sn`�Nb� ���*]o�1��gI����X9A���+z�*V߱'VC�z��{�:^V��Y~�珁�ؕ��QƉW�����Zf�2�lC���f��+���ٙwL�mC���HϗW��+��p2���o
X Sb�Rd�P���)���dF��I��VUO܇[���Y�yƳ7f���vLY�5���zK��-�*���K����?��"O�1�B\�����x�86���Oث�7��l�����Gp�Ǜ�B�J6���7t���Ĥi�d��~�\��Ñ&�;x؊���dg�2� ����x�Poq����$�shӟ��'�%_�A!U%�C�2Izp{�a䡠h^bD�ֺj�
b�OͶ2~܈<v�\sO��Ʌ2
�-�;0p�~Ye��e�mv&X�lq���~�/��ƅ�ov�lg�2�`=�Q+R!x�{�?�c��j�{z�Ym��=X��(����[��\��;�}�[E���ԏ�����r���6�h�a9Z@1x��[��NS���ռE���㬽Y_���Z'D��{?����=ɿ����l�es��.
J����V�~�,�� y��_��o`%����Ś2?�K: ��R�E�w�����]�o~�K�PrB��)��qJ���@��F�^���SY�_��y��JYˁ|u�����I��|��<a����,=�ܓ7a�E������6[(Ob2`Mh����D���G���˚/��,�s�!�(	0�ߩa�X`�7��r2����rnk�\�эL.SG�ɥ��V��n�c�z�p���\������_�f�R��D����lDG�9Ա����g϶=/f�}���$�W��������ԇ�y����N�z׉T���>�y��I)ӻ���C�O\5���BVE���2�B����r���F̎�����o,��p���ˮF�w�-��κOۥMc�(��{$Ӫ��(�y�߻��|�����,�Y�[�������,��1z�!��� ��n��#�����%�]��xa��kc��~&���L_�\H�"%x�ǧ)�E��1��iic��W�Mc��,*�J�)����̋؊V񘕗bkj�7�Z�����
�֫63_ {���f�����y��j���Z{Yܗ~yr�KiSd2�2���E �MQ�G�p�G2�R_g�z)9!�U��5�	������G��i�wa�/���aŶ��x|Eؔ��1�f8 ��+�.~U@���(�+��^�U�au����z�4|�.�0]�4�Y��>Tk.@��d+���5G����reccc����r����H�H:�W�Ӑu�� pb����$��<?����%,ҩv6�g&�k�L���o��q-Ҷ��3h.`ftJdP�W�����
4���3g�<՟�fIQ�>�U�R"���$2C�Z�����w��j� 3�����{xx�iZ`*����f3h����W�O�@0��R@���|�����_:	�>p��u�e�LܵL�ŭp�v�t�6��e����\�k%���������YDQ7����&A��/b����VJ?�!t{� �O]��kN����Y�@�X&������5y���w �u5[��0'F�4R`�"X&��0@�7�@
B����)m���k�=?���E��I�8G��p�K��ž�s�VHF�gIF:��?f!(�Y^����T$��ǖ%Rs���#�%s�ܴy��'v�+�-Rǀ�i�<�3k�̖��� �ul}��_	S	Y@z�!�?�Y"�i:|���]Ai�� �W�1:�:�]-�"��B@�gՏj��Q/�3g3�V-7��#�-��J'�g��v�໭�j���)�999g�׮��WRR��S�͡��3aD8l]
��$!��*�Čc�"rAP��7�YRh���_a	��hfA!�߱D�ѳ@3Y�Y�#x�SꝜ��&^�#5�nR>���-T��3&��C<�˴ix�-�6�����d�f|=#�?Q�88��=KIfK�̚X���AV��t��bJ�^$��|C���G��J|k˂$d��r�]0�P���M���v���zr[�7����A�� �gTUWK������~oS9/��B�I���=���>7k�N��U��Ο��^g�b����6�Q�>�MNIP��r̹,:��B��.�È�xJ���_XĹ����@��~6E+�����<�@(h@��/��,)����@�7
����˗��'"8�x�W�HG�5�7Tt���C�	�����B��s�����-�b�߃-�
��yq����V������3k�uzI���Z:��B�-�y�kJ6�c#/��}
���G��&���'����~p�_����?��:Ʊ�j]�QＦ&PuoA�;i&~�]�~ܗ ��&�-)-�1���	9z��4�dŶ����sS���t�U�޺jIk�ע�,���~>���n n�8|ӏ�fy1!G��ł$�;v�$�ixs��8�"�J����{x<B}�&K�H0�:
q)�/$6����SI���cTٙɳ�8qs���s�@+?�US��'���8���E�'II&%��[$�ݦQ֣�P)� �6�5s��,�pS&��fPh��u��E �!{#�y5uu����- 욇+����na�cm<�[
��Q6�v�D���I+O7����P�5�b6=��UW-A�-�%����ӧw��p6~"Sr�2x�0���-}�
P=����k��J�-�)<EF��>l?d�ڞ ��N�����V9J m@;�X�vh�?���O��s��4�����7w_���<a/:�����Ab�K;����vw�~|�$��K�_��{�t����}��u�c����%�	��F���@��{��j΢�uTsT�������r� O��?�}�%U�nGv>_����a��uXsTW��)l{�+��L����3�y�rܮ�v�F�G��c3�~{Dȅ�'��^P�w|Bbڎ��y=����O_�����?:������K���yfxw���2�x����`�EX?^����X������?s��`��{y5�~7�m�۷o���Y�Cȓ�=�O�gZr�nͨ��?�]�N$�`����h/=��WSS��~�{�p��E�=��f����Օo�����/Wrݩ4/R����A���V9���"�ᓨj���۝��IF_�S�	������_�n�S0�!2)�[���'Yc�U����spghQ!�o^ ��"����M5��/3\���WO�nt���A�҃��Z.�j�A��G��u6�ڶ���B���"\�8�x���A��Z{�j��,��+�Oۗ�\<�޳�gMɈ"[��w N� �?����ͪ��+dK���W�����=��v;�D�5z����}��y|,�J��j�,�z�}In�7宠�s���@����m0{�����CԖD���~�\�DD�����ʢJ�sd���������� �/�ĦM�4
.�	�o�1���%�79������B���Lsqq��p�5�0--M��7��[�~J��������+���+#/�j�B;�P�4�Q%�+�����7�psLO���F%�'�:��ܣ��C����6��^Y�+J���M��
¨L-�X��;*o�G�ٲd���-/a!O��8�Nw�xxz�z�1Puo�EL�A�t��2���̪�0�4p_�@�o�~O	�Y�/������_�}W�yn�z��eM�d�`f{5!`V��Hї���v��X"�%$Yw5��ƭ���[zL�� '���9�^��hi$��e�؀����Q�g�8�d����S�@�����'�986�([�H(�},Ҕ|��v�����]�rL�ki�>ʗ��[F��� �=�:��:�wt�K�l���.0�F�ɬcT)I���@����+X:��T��Ȫ�6�W�\I96�����F�;���������2��������>��eUYd$�Dd�>4-������̐�͡��y���$D1�@~�P���w��-��Br'u�A����*���0�Jq��Fk���/���4:�;��=:H����T���הw��;%����o�)kh yFVUu:T�`�k���os�I�*���nޏEPq@��� ]~�,���tBsԖK��A�a*.7�*�k<���m���hC" 4��'�S�8�T�i#��g�� �B_�E���ɵ���M=>*T���=Li-��D����b�2���N
�G  �:��&�ԭ�&@�����UK6���/���h��goʩ����`��-�l��?e������w9L𾥥E���>�FG4�}��om�nuuuy�P��=5̻�(�'�U�R�502R�D��x��;�\Ww�P�ˌ�Y�1VJ�{(�@�x#%�Y$�����֤^����];�Q�h�� ��:D�&Ꝝ�554�H(ͣ��җ���_��걂빍��x��8�[7eo�N���vM���sϵ0G<J�0�):lL��l�b2�� y�e DC�J�7���T�%�������̳=��'�*݇���V��y���e>Q�6��ل�"k���	�a>�PDR��8�F�0������+T��.K����@�o�\\]�"D�������}�-���	���nZ1����]�j�����T����s�l�#'N�+S�K9F�&$$0�Ftzx��f-��Rk�4<����u��x,���T�B6:���*Jw <-�h�P<8���wvvz� )BAeT$)�.������@�v@V�0���5MM>�$����i���9�%*�����:'F��iZ�I��gjb���W�iލ��qU7d;a��r��=ea����,n\�ti�������j�W��
 �V�����'�(�<�����TP@@�_��KpLp a����Z���=�#����\z'Y�xO���
�߅�FF[���9��-�V:��H�
a}����^��ƫ����I�i/�������9ɶ.��	Uc�$;̌�>{����9�9�h�����]�szP�`d�6 k�aH�H;��t���_}I|��FVB@�#D�������AReN 6��BPp�>��A�A������s#�3�9���_jk��@�������D���某4}���t@�i?�T�Q՘?=�[��z3�7�ir�}����p7�!���O���򽠤����t2�������[ʬ�|�@|ܝ9.��$U��d�,�#��_����)��ˬ����f`u�`XD��*!����ǖ?�	
@�اV��	�l���'����:E0�3cj���$8��x����t�1f�+�-�!���ϴa���� W�t���f�d����p�G���*,Խcp�x�A+/6���QOB�@���r�{��d �:˽V-�DH����0��ֲ��=��P�ĥ���tƔ�����p�;i���U3s�p�5��(���:�����)�FH�#R��(�)I�T��R���;������>g��0Ǹg��ܠ&
���Q�r����&�� efܞ�WՉs�K._�(�������c-�ؑM����������M�F	�|�h�c��u���(���w޴���0{Df|P�ڨߴ�	@�a+�H�%/����Q@��`P��Y,�k���Y#Z.D
D�����@s6�Yy�צ�� �2�j���	�67ņ�P�D�\P"(��=�?�۱uz䤦d%@a	�����R��3�K�H�"<�2��|���5��:EK������T�O���0�n�s���g6wXD?�C+	<V�D~D�[_�gj�{C	�5���3q��$︕��[EA�Q(Y�r�@�h	!G���=���U�)++��6�-���UZ���h{<�+�N��}��I�-�	I*����0˽�"4+`1�!�U"o�n��m���l�Ҫό1T��Z&C<�{��{�a
����7��3���Ԣ�;kS�Ae���_����\�sD)�_�C�p�(�9�����HR'�-�[���Z�dIY��<��𨅵ݻ.��oĚ��7�\/l��(��1��a�l�����a;�$��,8�;%��-���vj�]�ςN��cj��vR����m<���;�5l-b�^9�e�8k4�ǏOb�J�!�dTU���L��k)��R��>ۨ�l`�������ԋ�����v@@�;޹��mm�� Z������1>:�9�Ƿ�	l�PSS.r�
lH!�>�J߇"���f*3�1�u Y{�*azx龬Y֖U�O[� л��O�<ټ�@�}����d�v���X��A���x����He ������b1�j,U�Xy��ko)/Wd8�����ۅ-=�\��̪���A#���M�P�z�R��-�6�t��+�_Q�SŤ�q��dւ9
\�i��D7�f��74T�S�q�1
t�C:Ɓ�|wA  �t��W_z�x)��`yy�t;�m=[<�k;����q��9�a�G�fKο�}�ԩSہ1�e�ۧ��N睏p�*l����x��[�� �E�̅����Y�y�^��h���_��)޲���j�?^'#�����֪���Y��Ȃ*%|E��ͰM�#�Ǧ�V'w���{�,��WnN�x�X@^�`�a�@.o�Д�ࢨ>csҡ�{���N
Q�P��!3�3�e���&֫%8�13�R@�{��&���0}jh5y��E��'�A���>}�X��Q��J���E0��{��Z��h^�� <uh4{ `��� � ���h�{r0:���	�!��ԟ��Aû�KY����դ|!��@����u�<��Ev��������E�������=�)�yծ2���(9aޞw�\���YJ*<�Ѹ�b��|nLIz�m]۫�ؤ�rL�k���ZǬ�I@�5�<ⵦ25&��=�t{��1;`*�gD��a����j���v�����,	�T9v�T�/�t����Yjn��'��ٙ��=~��l�N�>��!1cP�
0S�aJ�����|�	�����������r�R���X�蚄GD�퀠v����z.�b �Ʉ��l��un��r&��%i f^|1�[������$>�W��U��W����-�����$�03��a�`	{��}��Օ�?<���_�&������_"�%���	�/q���9�D�u8FD�)�h>�5�>b��w�s��y�SE�W�-��!�"�N��L��I���ϵ��?WW/�73n�_TeL]}b�H���)�A;l���ݔ�s|Rgw�41�GyhD�7!��(�}�W�ҧ�Xԋ%>y�Y 1q��0��D��DK|��� A�ߩ����|�%��z��-�l6�}�hT�ͻ�2���:� T[�+���9�U"�r��(�N�{��N]U��W��B��J�4tevg��s���x�9��U���5��C 2��GiT��(��]�a"3��sPS*S=\��bDϛكnE�M��<=�E+[�ɣ)�s��i���P:����_�~����s�覯b3j�z����A�T�Z��`g�����<�˽���������ݖ,����Zb�e�E��������1��@�@�n�=��8��L�_D��S����`�2B�-��]z���4p�*�%�����:�G43�e�٠����LTs���tnRS�_x��Q�!�5�Uc�`<�a�K\�
d���>.�ǌFUA��wq͋�fx\�k�jHq�l�<�� ����YԓA,7SE"@򷐒o��rޗO��*}x�z�2k�_���n�:�� ��Z߇�!��;�=]M���96�m ��\�Ah[�H��)@!�F�� T�#�sE��)Ha�+�!��W����Xį�����
�g�����n��t�Sڟ�jhԶ��7���[�؃e=z�RUV��`�$��羾5��p�6
%:H	\���pnv4��IOsT��s�oR ��� �G���R.�[���*^��-��T:-%��É��E,�J�
���� P�"��&�T@�~�ص9��XN�����!ʓ�U��t�D��t%�e�[J����h��q��k��P YPg~��19qb�6[A�Ŕ����D(}����W�u�����yg�^f
�z��nT���q��Tm�_Z��!���Xj�D���\Z������O:*��ǀ�j�z�c�SQF��@����%JX/Q�U �L�]���I�]9j���(�;� FPk����w^���:6�B��'ʤD;\V�))[�:Ŷ�2'4%#�������Q�yh��+�_�?ݛ�ɉ�I�Y먙@�} �=��N�ߣE(&l�D�g�QuNke���9��tm��׷7���L��0��YT��3��;��z�M@ܖ��L���x$Hy�'J�P !B ��G<��1a@�VT�� [�"��������+j,��<�˗7<��zGwj��7�}��G۞�!-^�6,Ƭ��	���������Òo��M��9�!����x��iu@m��k\^�־���)��P�1D��ROJ�~jS�d�:X\\|q{ p��W����ܘ��2A>)1�{.+����O��D��E�9W����g���z�cx����3�����`�h�G"��j�w�a�e��J�QPW2�L��������T]�{{��߾}K�F��3�k�<P���>SO�c�n+�j4|�wGe\,8����ӹ�W�o"3�<�9O400ohkk�N7]��E�t�t����?��f�b�{������XOi#�����D_�fii1`�+pl�<���?Ք��dM�����%��U�H�h`�n |ظ�k�:�=*���ŝ{����ܔ��é��J�,��B�vM�L˄�����$�Z��Z�renVP�=�{�Yݙ��k~����L�)Ũ����EW������G_��W.���������{����{����{����{�����?�>X��cv��IM��E\��]�qM/jJ�����Y"
Q��L�̐�{���S�	"T��U�H�� h�_����Ƀ�\�4��3�x���~���vv?�	Iō�?�q�m~!as��Ο=�	-�^�<���(w���k7N��t���!����-�N��ԗf�wK�=�'�倔��ʣ_���s�M�*ך��1y�9L�W�7��GXS���t��͞ˈ�H�}Na�Y�/rtf��K����/.*�1��b�ۋ٘��q����O�bQ�p{�T����-��'#3q��s)A|� �v��K��}?��,�2aZ����d}��T�w��W�|ݰ��_O��fk�ũ-���=�J$�. �D�"��L�(����>��zA�\,�&t>�1�-PJf)	��t�\|�����k>Q3��1zBmK��v����� ���� �M�˧ܛ/�����X\��N,�s��G��l{8r��p ���I_Ds����^a�#���q�_��g$��Yx<p�c���g��|"-0����&�)��3�{������[�Tf�8&��3��0~@F�� z06���e���7M�jsB����R/1�;"�׮�h�3ϻ�k[:��IA�F@��2r�87F&��\���Of5j��-WH�D��C���z��������c�S}={
�`�t�!��B���Y�/89-mh9%Y���C�c���@u���7��F���s;�W?�qjr<O�D!�T����[�)}��1�;2�7�����������	]�_��>U~_�G����)�ᖿn1���x��vs#w�ǘ��9@9�l.E~y�7o��$8E6}r|8/�j,��Fz_V���\�Idv/��4�/���׮];�an��h^�ԍ���;_2�/���h�*,��$qZ���B��^����PgG�YQ���>r���:��������pGeyQ��=�����ӏqA�ڻ���l��wD��}���;,t�y'�7�!v������6�������`wFO�x��BI���q�b����"J.Z(+Q�R23� �sR�O�xO����{.����Q�P{f%=���9x�o�t	9���s?��(;{v����ӧ�H8}*H�Y�&㾫�5%�XsjJ�	 -S��J��x��`/�1"�xr��C222"����ηK����/��u���u�HQ�>Ǉ�2��6�F8w���d����g��	b�TY__/�� �M+�щ��m��<+� j-8�),���=�X�x1h�a��t�.i�d�Y&�W��	���ܲCX�%g��d���1Y�O�4�i�a��^�ڬ���̲�#�=H���?�����C�]/���O����ej>|�R+=����eG�/�ͣ��|���5�_���,�}�����?���h��1]�ۇ�G��F'�5n�*{>�������7���R�GmI�D�\ض���MZ׶UK�W�u�w��kD~�������/�7��V����L���<����_p|p�ޟ�m���%�\���O�`�m�E1�M��a�g�
����<�-�4�o����;��	I��g2��y��.�P�$����YU��E݄�[/j������݄u�n����pB;;�ҥK�{
D0GU��3ed�n�΅�7�3��~��U�)~��ݭ�<Em� "bS��nd��ӳ�%�������}%����$�����ÓBm3,'�S�c2�(��Ú�_��[��	�,��v�����~ʅ�`Ƅ��7cI��/ӓ�f���ٹarrl#U�(�Gl9%���� ��J�Y��߿_ے[���-���/R��ĉV	Θ�V?p���j#�p+/�
�t���XΌ=~<}3�;�[A��v����)��*#�����Q�
k��4p��a�J��+�a���^���L/���o��LX3��!������X�Ѳ��S�	�f���E�p;�3Y��v%L��HI�>�+�g- v���Uɦ��uw�o ��m�㘤CK q��{�C��?O}ɶ��v�����J}���d�Գ�>�y>�*�0�p6�����1d��F�Jo�1��9�/��x5M��r=`�l����O?'����I̔>�&�&�a��W��J��RHHH'��q��n�vk^J|�0�a��.�"���Zy�}y�ۃY#OO ��}"��=�e�I�;�ֶ���sjl������o�}~b>���yY%���\@���ڐ�%�Bt���h���jrRǯoo�TWW�HS�Jm�h)�ɳ/�J�r�$[&x}N��=d�ʌ1�U��|e�M�LfՄ��c�P��� ]c���N�Dد����������4���%=��־	`|{��s�[�@^0�TC���}��Xt������X!�9k�(�e��B��҇���eژ#��.s�v���6�#6|�4�ri"��A��4�M-�H!��b���E�A�-�g��=�ZI�NNŔ4b�������L�R^.B�`U�L�o�'���w�k��OM�Ht?��E轎 ��a3�OWn�}X��'��-Փ���n1_OMr�0c~�j}Ճ]��5��@ ?�aP�ΌF��=�D|�	�7���I��E(X�u?�^|�������gD��O��yd��U�.RAnqtP0��#5` ^w������O�voj����(����[|�iM�� G/�efj�)Dz9-]x��,4�y�R��ku���/sm1�M�Dt7c��Ε�愊�Դ��I�F*/��df6 �M�FY��[2��R�S`Em��w���Z��Cf���wZ��_m��8���4�S��c�.k*}��&���狘�3��U5�jj�Ȭ�bJ_�Z�f����!R���گ)��D	m�$Y��Q��i�}�����{�Y��rsX��P�	`���>��,#�I_����M@/����]�SGG����f�yR�9��Umtn�tZ9^f�脑�d?��&��ɮDɭᙢJ�������ɶ�D�(V���
�]}o�Tf*��0x�V�xzw��� %���G�H9��"�}|*��.���`�gTm��4��
M�ϝe�O�F��2V�U��I��y���. b��	w��Ɲ�ङ�ȴ��/_6�(�H��	$Yvрe�p-�L:wt�c��}ճc`l���:�3;�|���&Y?��č7b����ĝ��Ʋ�qW+��L��� ��C��@d��% �p�ya�{���Z?��My�Q���H�Q�h�ff!ft���9��/���ԩ�?(��c5'E�Qf�3ο����ۓ'z<D��Nf��Me��ԠRH1 L��
[�I�����O���;�
z���� `RzVR�&>��%Zx@M��=��'�Ȓ��*U��KA yLEL|Fz�d!�������$O�����Yɨ�S����ɭL+��H��"Vj�ƾ	���?8�w��D�c����<�S���K���`|H2�R�8����h�=�j��!���Df�o������d�Cx���&B6���>v6o��9�$Lѐx:N��"uʖ,�6��1m�8Y�<*�L�%��S÷��&��!�o�mdV�h�	w;0�k*���p�w87�/�H�+�#�a���^�w��a6��W5�����'�=�6��9܅�����A�S/����J̉��K!�V�o��a����!4̶�̃* �VU��5�MJ_���������o@���2�%��'r(�'�b�.m��Κ����'�����,S� �� �>}��0�2D9���!y�P�7@�6��Q��gN���&Y��N��ɕ�i1ÔW{��\OɶjP���&>�+L\#��xaKK��9h��#UBv�}������!X>�/	K�Z&耜�~�?P�:�m�EU�)b����b�m�س���D����\D�-`�����^�y�
6�����qn�w_�(���~1��@5��d�������ݺAN�'u��u�q Zb{ݣǎ��Q|�Q^UCւ%`�J��Y�������qZ���:]�\�G�q�v��4Cx�G��zYn�r8�oa1�ݻ�hp!�R�p%5���
����|��XF�5#�Ç��1h��㫪�ʮ�����`յ�G+x�s:��Z1���� ��һ��~DIM�}�c�7��\$���?f����������1�Vو�!=k�{fg�s�T���v�ya�uh�ٷ�(��m��eB3�������(��-`����B�r�u���k5N���� �?MI��;��v�����V��QU�����G�p��e���z��=�F�/�G5�[����Rv�"4F�
����VRT#@p�^&��b�y`�?OB���9��Q���t0G�$��pF)MI��H����y��Fn�o��"r	���M�:�ѷ@���OD�xt�6KI�(Q����1�[���jeK���
�D����#0��㣪�Τ�)���U笧>Q�>4g�0��1�=Q��hE��8>af�l�Ɩ?�uA��wZO����r�H<݂�ZĒ�˝���R5]Z��L��X��M(83���"�M�;ι�����vV=f�ut�s��#�^�C9�$�h��ۿR�h�� �E��+8���\}w\�W�~,-؊`j[P��#*��B��F�DC��@�����Z� Z��@���=,(dh��1@DD6�������W�Wι����{]gžu#�v��! H����2*�ǣi�D�*�
]��~���PY�\�.��W!��21�ǫZG��'��2��HSg�V�Wz�n#�:΃�⾭����2�w��E}ۊ�-g��Q��g�H� �N��O�nR��P~z���E�po*�
�������_�:f�=�ɞ<�jW��e���G��Pr p�W���i�=�e�r@�	4HO�^��ҋ��aߝ�Ϗ#R��)�P����-煋�PR�!Ϯ�qD�_|s�.�,0��QP�;xJV[�j���Ml������U &��[u�/�'�\`�E��?C1��`��aP�}�pno�Q�#��pv��SJ�;ЛSu�o�X>�D0ܔ
��Q��� Ů%��z�a�Pt��"��$p�!��V�,�I ��u���������ЫT	��Ϗm��1�P�/<Fz�gp/�PI�6�EC@.���a�Cna)�v���Xs-�ԃXU�#�'�X;��PBg$z�}�ȭ���O���vw�L��aBQ��x�9�waP܂�XQ-~�;Qo=��Tb�@�\��hF�-ɳ�"�Ց��qV�:�Nl�+u6�?��U5%�]���}p|��AU�%��<�J]�f���ȯ5�T��4zv������`kI; ��QJ~.�8T��x�]�D�����t>xZ,!<@��B�s��Y����o��6*��fý��$Q'7��x��lo?t���n@�~��1G�Ԏ�]�r�:؛�ga�ʄ�mH�$? x�V)�2�
����I����i����˾���NwHj`�Vxy���}'�)�^��D%7�ѧڳ��M�d�Y�S��R���zS����G(o�:t��� �w��R�fM.*ľ|��V����$j8c�=� ���$��.>���[��<dǜw���2Uѭ����3(�WAE���O�Ą(�i}�	��HR������
��1��zN�hÙ��:P�Q٬1A�[��H
1�'���.R���9�i�TMTn)�ڠ(��3e��]���2 ����t����Q��D�H6Q�x�A$ᗰ,�W��Ӻ��fh6�U>v�<腀=|ly�dC�,�=[kbf�m��L ���(P�y�_K�[,q�]]�$�D�>��;��:��k�ѻ �VՐH=� Y��f���y�)�Z��;y�=��|����1<w�_�QZ���uX@����1��Q����oUx�; �'��r������*�AKW�4�7����]�}�s�5���4tEfh�͹%5F�����8ׁ:�yq���t��^��"��"���k� �h��~�N�Xu���頬@?j�5�P���L�Qc�N"�~࿸��lڣC��'1�3�m�635qv0�&CpH����Jidg�gT�J�F�e�+(�����aB~�a����+�߻6��D~�[z�u�Q��o����<��]>H`|�П��N$@�2�W����jg`�$�n�e^�e!���F�����Q�N �%)���ہ^0������N��x�]·W�N��]�.>1?�)ͼ$�� t�s�*��]����Ê1I4�+
E����;XΓ���u�uc�:q]~?i��|�m� c۩�kIU����O���*v��a[��P*�{��_�8�̄ң�Z�����5���Mk@��͟����~�q��Y�!�^sq:;���u��ڪ��U@LM( �C�J���kbu��b����ͨW�������۷�,��=/��e{� �(bO>���hsɺ���2�^Z`��l*y�x`�7��8��$��ĉ�������u��51��z;��B�:�nWe�H���w�Keu+��������x��ط�8O1qE�drCAI�FJ���?H
j�m
��
Z�'�T\��i*+�?�bk�`I��9U�'�ʂ�pdo�B��R�����d^s�"�U«��_�jI|sI����#"a&[Kڅ6y@�:�dl�YP5�G��~�.C��<�ߌ��X�zĕP��R�L63���
�3PS���v%�#Bΰ�İ0��Y�No�����(�;�u�:k�%ꌀ��_ݬ�¥w���pk\����f~�@$G��d�ݻĞ.�f�%�h��VW	߂h{�gR���j5��.�|����#Ǧ�`����%~��]�����ʖB��Q��ITo�2#��3���=e=�:�bÕ���k�$���W%BrN�͒��>]Q@�ś�>'����]O��n{0�q�&wC���܊�}�~j5���]G�����ߔ �����xǫ9�8z�$]$�4ںa���u�ڲ	j��/G�"��薂myܥ���2�c-�iQ�7V3��̀��"f�~�_V>�P�ׅ�<Ztk����k�&|�ߣ�r��(�������C#�@}г[}��j���Ib��A�%��>+Ѿ_���P��n�R.��. D�[���) ㎿�x�g�y`M-C��Z�q���a�
F�^���|&*��iŗwL�M$5���ckJ�ï���[	Kes%�Θ�
8�M�f�[���&	}��C_2
��)i��_���P�\�x����x�����%liB��ؾ��w���6��rY��,q}�9)@޲�d�+�H��ُ&����DsU	�-�W=��P��?R�y[<ݷ�)���A�aɯ��,��Q�w
�M���CF+�����Ft��7�����[�"�z�<]s8��OJ���&��a��M��Æ:�\/i�x��ߙ�E���6Lj�#J;������q���.Ȁo���@�#:�?`�{rɵ*�9����vb.KP�+����}�@��'����B������$J�r�A	�&��d5����Zt�D�k��=�ڕ��S�+��N��@��A�;	a
������v~�2����i�7Ua:�=|
�
�mF�`
-�q�B�]z�`�Ҳ����ӧO;v6�u�x�#���61�j��]ؽ8��<��o�u��qqq��kgݾ�ʊ1T.���f$N��Ils���gL���w��"��� ��*�Fv� Js,+���U�c_�k��Q��O'hpUB�p��W���5�NLL���A(�h9_6����+���_�p�w�4������0i #��
m?;���[^Q1�'�7h룺>A�w5�g%1��݋������m/�7%ar�FY+� <�w�
mƥcW�������y�dU���}7w��M��w����bq51�$���"�� h�k`������;� &�����ӧ���;V ���%��+��j��v���!C�K��s����=�q���g��")2h�$�]���j0q"���h
�����(��ᮋtq������,<���^�)�� �1Y�����-�a{�l8�B0X]���G�>�
=6������,ܾwb��m+z���i��d3j 8(
���+���!��xI{�x��R�� S4�p�p3�8��4���R��T��@��ɳf����o��F�#hlh��^�Lv���}{�J̿g����r��}��0 �c�d�^��*�h��q8���R"Q�[2���?K������q�Lv8z��`�`���)DW�w��������[�6��v�$�hL���ZB�=A��*�rBۊ���^x����fj�k��	r�v����q��Ս��xpEv�-��Ką��� ۺ`ʓ�Qsu��|��O�nj�u��<����O��\��D�NHsug��- q���ޛK]Z
,\h'�����gn��\t�o���m����k�N��\@`<������@�;V9�AW��t�S�p����;���@��apg�T]��'���O�P�?O��f:�?z������q�;U5kDڄ��WvxHGHm*�X�x#J���aT��&�>���C�7c�<u�T*u��I=~��;���b�L�B��yCZ�s��f+���9� ���~�.�RR�����F��y�\v�4�C7롸6�4����q}�':`��'$��tM}dO�#[�D��Ae�իW`�&c�n�}~�=���K����X�����֦A��ja6ݖ�vz�N0}}��tW�M�P�X������=��\��<�7I$ �WDĔ>�.C�K�S�V��Sh�Xx��Lw�� ���x��@�KR�)���F55�8]�~x�2a�I����!�ܿ��o���	&s��ܹs26[��%{w%�{U�qM���|r� :#s:�?�6� Yh�v՝;�L�H��w��§�6ZU��!Y�� �������B��������3GC���-,��]�Gz�@�I�8-b3�-�kd]Fφ��bP����O�1�J�얨���(c���*��H�_A�nq nS�)_Ie��i��UgN޴�8��`z��j�Z���]�?zl�D�A놶 �8�ކ`H��l%����H��'����E���ﭐZ������X/�[1�ᶕ�5h�ͶAe�q�d�
�؛*���}�+_��i5�s"S8�+j���1D����*�Xy���v�;���'�1B�8<DrN�g�y�g��|>s��ÇK��m^��Ks�/�.s��D�B��v%tZ�Mi��V��T-콤�{�=��ža�������J����.�\�F+߈����n�>h%��ފ^qlR�+���m��DE'Z�6hU晋��M��3w���U� �R�����H*�x��?�� �?۬��XK���_3{����N��	R�M� 㪢�Z4����,r�V�0Rt��<���_�n��WU�r�e���W`�U2��ۭ�d�k�xb�YX���Λ8q���\��Ӵ���D�ϡ�l牘�X4w�7}��kkk��^S
���Zɮ.V��7���,8�_A)cw�v�{�������#��> � W��yMh�n��J���d�TN1��"O6sy�=�F��ּKo�r�M]�?�����\]9�_$a��q���htT/j���c���,`	���M��XIE�%��U��%ZV��a�"74��[%��!����2����PV�Ƿ�O�r%���$m���I��oÇ��2gww��T_�kcP�Z�֪�E���_,#���СN�2�h�C�%�<��O˟ �kp �����?@��C���Rh;+~?ZK�?�D6��|j��T�,���;wF}���X�W{i0Y.$� z㕅V�Oݯ$�~B߶��>r�u �|쩟:�����������z�2J��%d��,b$AM��.��9���ȵ1}u'k�S }h��GߡZ�o��N��z�:�	᧽���B���Zv�X���@��"��p!�	�=��w��XF_������V ��q>���ж��؉������
2�xǰ�}�����a��vttW��A�<B�ۀ� !��h��v�L��c<����`ojz=/u��6��,��JF�6	xTn6ͤ�oBP��`�o�	]'��t��ÿ,	�Ln,��{7 �� ���p�ɷB��@\`dc��a���Ƶ_+:U�lν�Ю{r�@6�zwR�8j��v0b�Q}���Я�@����X�y_�tÈ��1f�Z4�:@J]��*Z����βU��mF�֞�ON� �Ԩ�Pߡ�V�a�
a�+�)>�y��V�:~nɈ���U�ԧa�D;���V���������[�掘�.iS��®iOuT�f��{f,;�V=���B��E�L<C��P��g�f}�A$�xJ���s�{��2�*8YX�ވ�(K��[��C�lq�bXz�:LS%�P�7k��&b� R���o5�]CrG��7��Ѷ�6�/��A�(����T��MB��D!�W-՞(k��;A���-	$�ơ*W~O}t�8Lw�;�Zf՛�k�E�"N��/UI��~���/V��K���/�R��h����S�D���\�rv|����Q�yCb�O{��l�O�ʄ�\�5����Wʻ<�+kۺ��璘Ign���8W���Kv��o��J�����n��W���$qo��D��W[7��>}%=�r�xV���~�����1����{��Ky�x
>io��i����=�۹��0��?*:P��:�S���g�f&z�����ioʉ�#����[,��:H7�����:qa?�wg�v$ �TȏaH�vgB�)^d�qS������N�85���vP y�E�u9��̓�f}�H�����k�,9EeQ� D�滋	�U	SXz��i=D����;���c��(�	$Q)���t늪�BK|-z ��z�u/�U�cR�>�*RAm���ćL?�]R���ek��zSĥm!`� �v��?WXs�K��>��hc�!h~U�s�C)�^�61�Vi�����n/��OA˾Ѓ�8�@:(����+Ո�{��}������S-�bJY��}
h�GlV�Ը*��&�̶� F��ߩ(���gG]�M^x:=7�c�a�A�n������߾�p���:ZX6p�vĭ�x3�u�V�1��G�B�0��W�#�<{��h�����M0����:�n�Ӌ�/���9��{J��戁�Lr�K�2���:Rs
�Nc�Ys3������ɍ��	]�����[4U^�X�����񅣹��#�|5U��`���;h�|f���=�zSͤ�R�U>fA�E�;�2��&f�g	V������n�����J��p�
��d�g���j����P�e��������Fa�Yݳ����ׄ�{�ȼsi�h�ށ�t�.��.�&�^sQ������"^x)��F����]6��=Q�	�8@#���*�%`������F�ʞ=�FV�-�,|x��J����X�H��q�<=3������L!9'��0�x�l����U&�XC��؟��Z%�J���@	��Ѷ���r]�K�_��]Ƞ�� �kk!#��HG�������c���,u��b��b�?PE�:�Lm�īI�	6���-r������uQ����A�����l��~4�Ъ��\��X�g���E�d鎜(M}F��vIeQ��E�[ZZb�j����Q��5�@���oS�_�[7�D�-z���1I�s�n��#_Wch����� xÅ�,!�����tHcj��0Hwvrҡ��� ��L�#��p��w�O��!ԓ��[�7���Q���M��¯͔B)�@�|���\\{��� ?�^��� ��ݽ�;F�@���1U���C&��I`����?^�I֮��&|����s�Uh��z�s8#�e
[��en16�ŝ�O9cL��T��J���v!�
@��(��c���B~�n��w�[���:�ǔ�㱱�x%WV<�{���Q�K�E���:w����3 �כB�J�2�YA܅���Rq�����XjtQ��.#�M���dY�3���6��u��(ט�>vbSmA�x5����qF�O�0ƚ:k�Y�Z:=2B���PIؖJ����蛴�)}(i
�A����n ��-�t*�j�t�n`a�8@��|��we��B�w�r�-�pA��l�0�r^3Am�ƍ�U� �89]�n8	��ؿU�l`BC�e���HP��;���!��S�9�)-�x_���9M�Y�Q*kj�$�@Q]��E�(Hܫ���\��w���&*:á�s8�����+���{��R�[s��zf��~ '�a)�w�����_v]bw�I����Otz4���z�p2�Q��8Rv�)��m��v� I͢'߻B�؃r0�������x{�Y�l"n��k>��Bd�#�ϏL,..�%��P&9��������55\F\�A�|gݐ)s@@������:�����@JuE6e��ɡ��xM�oz���E���1w�\�w�����]c������(�����<P��8Hм9�D�5s32�}e=�a �E���I�ŪYOqB6���fnn-�Ǆ�'�5i�j>��צ,!��1b�<t��~��9x	K��L�r�[g���/^�GRg��,���+�`��1�_�#JNEA��5�%���ׯ\�R�G@�J�=q�w��A��?�C�M��S��V�$}���\z6�]���[Y,V)+��mt���q�Ά2�<ivkd����l��P�����⡡! &�3��G��!�g�p��J��{U����ڒ�nK#�C�� ��6@�)�X�b��Ɛ���(ۀ�χ�&�*E������N��1�i�Lh}X����]�|�_��}�d����\����d��XWtE���˗/��/�υ���0�W�:����ds
�3X���yF�*�S�v��ӧ�$7ؓx緯�$�� vu� ���̬+��������\�j�~'�Y$=v�P�k�(/���L�5rR��w���هln�n��xd�:y���aT*J#����p�����۽G�R���{ͯը�,ۖD�Hnr��[ت�[�]��ܽ{��vY����<>�j�A�=N�{R�vel���W�7��yx�i	0�B�ͱi������W�@��= |�u2/8��u0.E�-��V�j�8�.�D�Ȉy�x�M�ط��!Q��D"V��[�ƞ<����/��3Q���~��(����1�$��u�S�cc�#]� sTR#�(m+�3��͵����/r�Ӭ�ԕ�o�f�K����b�P>�]`��a��֛�: ,ޖ7�U��܌�a�����\�F����w��ʟ�s�u |ۿ�
����슴!��oy�Y�y����P�9���k�KB�K��$��QU���ρMJ��߀HrZ���uB�O=��
%��83C�1��8���t/���M֒��˧7aG�.,�"�l�0�����߂�r�,�d~+I�*�܈��rs��P���2R�>�F� �E�����D���p���EN�!4�/o~<77�E��@tjOd+0�5�\Z#��6�0F=Z�6Nn|=��!���
N��qa85r��G=�s@
+�G��^IU������=@�><�3�|����.�p���f���=��H����y���:\V	��_�����`�6b`/�C=^pwSS��G�<��&F.�ã��G�����2�L��' ���@a@� �F&3������ե���c��}Y���}�1�a8]Ț���&�.�m�f{�n+��$n�ܝ36y�ѷ��a�1掝�޶?Zh��q���_��kA�v	nHQ�T�j@H��41�!�K��g�P$�6xkc(z��Q�N�[���bH�l��8��E��j� ���8NG�AC�:��8:R0�t�p��sRA�3l�sT�Ǹi��|�}ƞ�x]�g�#�m�5#ȿ���*�)��$]>ifІ A"�e��#�N;:X�Oᵙ�=�.�XY����?�~<������q�O�.�����`ӎ9�^Yqj�CZzz%O	߭P[��I��XD�[�o߾�j�ޚ̈2��D��@�cV���`�������J-�/��	9���z�\�np�M�;t9��@�y�s��j���c��e]y<�I'f
��#�]9s�Ӳ���vB_닀(ȫ[�q����<��"���a�W�q�ޙ���8^.�(4��o���,场2�MՑV��fbS��$�������5¤je��ʬ�W��l���L�a�*���ax�b➮k;*���y�{1s����-�#X�E�З�.��u�>lZ��f��z
aWo��LdE��*�ٰs�)Ռ�i��
��F�k)�9�"��ѺA��;L��w��/�6@��������eg�Yd�*�P-��㶌:;�5�G��=��Ff
?���7���oTt�����G5�#���&����A�(`����ߊ��ܱ.�/����w���&�CJ�"�Vc_��j~�FHjf���!���n1u2|xc��L ��io�i:l��>6� ������!*��r,� �#^�[��$��6
���O���'�B�.F���<g��T}/U":-��CtƊ�*T��t�q���> 1�;�|�y���F�й��]:>�Cm�@FXOD��Y��c�6�Ǩ�le
c=$�R(w���Z2i7�� �ssS���c�?n���]@�H}��X:�$�������c]��>��W�E��C:�	B7��"��΀������4������^\����簉����S�ҷ�����U���-�~��Ɏ4�Dv �ߐ $!�n���C�

�ZP�j5���\��4�&�՝�\>��^Y�I�̽���4�JWz:���O�޸fN�%b`(�	�$vhW+������B�� "z;�;��q#�pD��c��}��Ff��BH���7��-y�3��=ˉ�Nb,�Ya(�����\�=����}b S.DLg� 
pZ4�G}��c�������>M�s�OE���p��z�`t��-��H5%XQǜ�j��c�����E�Pg3�!+H�	�'�@�p�p$��g6K�M��wcY��i1k6y}��c�#����k������s�1��)��6��kpcwL(�@!�j erF��NIHUqa�{�E��Ř�^�	::B��D� 2��*g���R`y�7@��Y�WáY ���nwyjj�v$�TLm¾:�i��f��A�HU����bq�=ׯ����t�o۠��%r�������H�VB�ie�N� �4���h����ij�Ӭ�c���5ca�|R~ 7O�cŤ�t��i�X�V�f( ��,[@s��X����(:Ϧ�6/Y�DG���2��=�L�U��� ���Y@Z�d�a;wn$\��G��bn���ίN�O��Kݳ]���G����5W��D�έ�����ٷ(��ര�r+���7���-�-E�A{Di���3-+
���p�@K�bӠ�h�� �����|X���b�� ~\hYm��J& ��2����2-`��!i�
��;��p�S���uN���
^tHfKQt~$�H~�.D���t,�j5�2�N��!N�U�=?�:��{�S�˶%���>�nZ|~M��QO�7�Qm���Ȉ���K"�eG!P]7�m��J#_�A���5y������O��7��iS,G$ �Z�3���d.h�X�@rm�{r��S7�C��+��L�i�ѡ���@�l :;�L���9�]*��b���h�욞���0m��e�� ��V�H$���D��l>S�,[�ߎ@�$�l��i���C��mz#[��9L��L�ge�i�S)H��͞��6��??����w��^�N����G]�u��+v��I~(�<��i����>$�C+�|��e�;,!��@)=���s�83����?[��s��}@+;%���� Ϛ���tI�H4^��o��bڎ�����w�d��[{����W¬+��<i滹���G�������F���<�b��f����?��X�	E�Ⱦ�
��0�^V���{��Kс�������lX�����<1�ss�#"�� �^"�X�]Z�IB/7D���Xѱ9�$''7w܏}|��s�;(ȯ� &׫��V��]��tV��V4&iE�Q�1X�-H0��blqBՕ[ۛ��@�{Y<�;�1�L������~�kVb:�b�3P������A����ئ�������t�
��ԚK�ᗕM�u�M��5�����=5B� л#��
b`��?��Qb�aA1������+�rxn�+W<��&�_߰a���3�U�RXe�OJJʈ����G��n���i��c��`_��W:����&��sZ)kI�ؿ�Xi'�K�+!%|�Pm�RQ��l:��x�j�����]:
D�������˔�'�x�3�2���Z�R�+~�'M�G܌�$�L�Q_�-e�!�)Z���I�ؓ阩�7���[��44`���Y���D�|���� �1s��
��Q'��bG�w*�kf��l�&�/�a��HO�;u��P�dA���߼�/)�����?��ٓ3�|� �a/�ZRTѥ𔒓��)��	I��/�CM3�*'ԧ�c�6�γ�� �1��u�kx۳�3]a&0��P�]�A_ƺ�`�������\?$QT��H�`e�hh}y�ɊL�؝�J�r��?�OhoeL>��+u����N=��_�-�tr
�a���%�������tgyyy�n�=����&8Ғك��AnS8r��	n�`#A�,���Ƞu�M�E��M:n��������R�R�[W��ji�M��C�>��^*�;�P���P�*�N&a���G��9��R��B[�ܯԮ��|SuH|ᶠ���Jj��A�Tv���ن�9@����kr�1�L�8��6衄�=�X���~ғ�h��ȕ�����d?6aG���~���7S� ����[I~�^|�YQU5��? �E��O QFFyoO�m ��h�hj��'���r��	$Tw�9{����m���D>��0n*ݾ���Urp9��	�r�6�`��b�#nY��M�q�؋�� o�&�����qn�Ѱ�:��kbf��#vX7(�qpRX5�I�۹������?����$���XErLB?����G�h7X����s��E�=��'�����rs-�~;6�wXE�%�톐��������S�0��}�%̈��7Mr�]�­���O6����H�_N���c�Tˈ�16��1Ǎ�S w�Ȫύ�%[7��H�\�;�M�] ��r"H��
�^�>`����i"�g�����=��0.Y�i��]sZ�s�B%pJM�I���u����.�l��x^���=�/3�Y�������0�zَ�`:�4IIt�Ǳ�E]�:�%[Օ���V��˅�����ᬆBغR7�(_���Mk�ɚʊ:d�-�����D��xD�8�1��Xqdխ���\������8���IV�1KOu�,W �VVbJ���v0��v!0�VGZ�62����_[7,�l��$* �&�̙��bj���ˑ���ñ���+N����V����H�����_��+��_�f����*��,]�m��_�% rX�խ��<�bZiݾ�ǗH�2�jo��[��|p�����0�m���se�m���ndo%�}���pv| ��R��!���@{(]_�9lH�
s��!�����/h�N�tZBZv]��s=�}"��2�d���r.m�����p�{/����B��B��Q�?!�ĳ��y��\1nп5���io�a,�`O�v�g�<N���ř�j: ��N�I���Ts+�lbu|v8K�o L�r���l1�L���1yT��Y�1s\�|�A'�§�_���*(�c���[~,: y��%=�!���j�*^pY����v�@8�fsK�����h�N��P�y�Oe��ָ��\l�8����$8��C�7����^ق'�\�3&�i�q�F��&�O�q���~
!ީDpǙ���#��X^�n���nJd��ax���>�0x��ő �oހ����b�R�Ց�Z��&���؊/qtj�X�!��`ɸj�+�(� �m�B��"���G�M7Uȃ,�Ҫ
��`�%�Nm�(�b���V��/d�.�g�yfC��9�������n�\g�E������ܫ�ϱ�!��E��
�uZ�42N�i&�'i��i��iqA�>�qB� ��۵��=VW�I�8=�E�g_��^���څ�Ѽ�`*ّ�U���?�#o�1���s�rW�В���O�!Φ_l��,[8���v� ��3𧥩NN:ivk�v�n��@ �i�����gO�'
=0���4?,,ͪ.**��7�K6�YLi/�^s�#���1c}�O�TW̵��|�����I�v1�$���.i
�����	,�Ae���I�N�EkyT���x�f~��;&+�}{���[x)&����������8�2�V6��տ-:�K[N����.��q������d�6Ԇ����?=��Vy��/��L�����!�G՗�\���8�
D��<^�C��@�Y�@�;�U���|�m�<��px��<�;�?5[���ZM���ͳ���Wx\��4 F��3�Yg�`	��[6�a���V��:˰�Y=���d6[5E>���1�����T<Z�����p������A�g;�u�c[���R����x�R��2�c�>�-	HM;	��		���������.`_�������S���'������8�>AJ�ѳv8��N68�V�թM�z��*	�+W"~�I2p����z�e�aZ�2���<β���rdh�oA��<�.t�\#�`�;b@��6Z���򣁞r�˻���;�acN��dҝ.)}���9���D�}�2�q�4%�<�Βe���#��Bܚ6Ч���tJ�3��M�Uʃ��)���b1��1��>��oEY��=��ӲsX�_��h �S�h�:h��<M/�s�
w��؞*Y��1L��zAԐ�G��6���N���F�;���!(@����m��a�+�c.�����:�l��fueK����z:��P|c�\�Vu�Eo�o��]B�R�''C���M��s�F���z���+˞N�5G�]�z��!Ǐ�i�+�9����E�XG2��!�M�������)P���Ic����(^|{�Bض�l���-W�$�`z	RX�zt��@�yj��
e�:��}�0���	��g|�����`	�7+#U-��?�,�$����]�u ������2}̵kѡ�yH;��b2zԟ&� ����׾����O����h���=����yi��0��>0SDAp׳'��U���!t��sCY!��:�l�����Ua0K`:zN� ��8-���	����nva��~�]���^)bOc��i7�yw�vS9���`4+��?E�G�cR2���_�V�H5�I�v�����`��o���s�q�N�u�~�/�;i����?�N�$���U!��NN�����	_�d<��	ٽ�����k� ��A�����lh��1f&��aO�E�A�[�H*��u.���&�455�&����R*�;���҄�8
} ��H�2=�/�o��5w��٩�3�l�G�6l�ZN�_�y(�V��ރ�w�M�;�9���U�� ���q}lKu�e܂U����)�����[�#˲5�/�[�6������3��e�׋��V]]��z|�d:��B��,�ڴ<56���gds_�"d�׹R��|�7A����u�?�k�ZX%f�_(��ٔ�����Sɉ����XK~�-�𢓓��� ��a�~���9�>��P���W���	���$�_!n�W��?�OB�t�(:��:�����Q�` A�I��b(Z,�~wl�����������1��'�GX&�"���0�\���.���n��>%�4�4��uF�MUAd�!�q�Ȟe��XO���bjY�_���3PW&�$%��}WQ$�/�'��`8֒䇡Ϳ͟"�O�t��V�n���w"ޡ�e��ah�k���m�s:u�k�f��O��np��e�xf}v�e������h-�g��c�Z�����O)��%��� І�e&$˽���n��ҩ�����c}�N�ČU*=[�����L����f����v�g	�=s���/��G�{�?�v�� �a �uE�����
��LfL\��Z��N�C/\��4�&�b'4Ns�V&���M��/殿~��>`>��}|��t�/�?��̈́��X���U�oM���s _�������m+Yf���y����L�G��a�vE� ��}��C�ñ[ĳrZd�Z�ӄ�~��HMM��
aw�8dǍ"}���2ԉ�'�<?���lo�W]]�G�%�Q�rB})z'�L��؇��g9��y� ��ϖlq�@z��+��펢SdR,�6��c/T�X���2tgy��������J�D�@r5�!���S����z�L�t�C�P���L}�Y�1���	�d���x8���ɷ��!!�ß�y��}q
=ҏz� w�d�M�6:2��B�Y� �|�hf����v���&On�����Pg*�S��vg��Zn�/zm�Ν;W�-Q�o�B�ڷo����]�B����XM��y6^g����͐c+����q�M�l���f@@�|N,in�t5z���x/U�S�_��)w��ۿB��r2���1�_�`%�6�I5м ՝�@�PIw
˲RڥB�͏�c����9��������WT	�� Ų$�]��p聳l��zZB�I�ʂ��6q�ʪ��K^�; �̍�B�����
TG�!��.�m�m:����G-�u���e�mUWH�MV�ޠ��ͥ���5�ҟ��`}ě�+��ܱ��QWl/A�Bn_R9
�֧���VO<��s���xM�urj�o#�(��d\w����>W�i�O�ܓ��5
a����;���'�Cb����tӳ#B���q��6�s8Tu�[�� z:_f��ر
i��F���45���m����Ճ�m��p��ne�f�7�Lb�zm�4�D'T��L�v}x�g��J\���J�bA3z��:��"{��e�UU�o2��9��(!H��<��	��I��,����yA5ڝ;�*̿{�nF~2� �+�p��q���	\<<j+�����2������w"�}|���Đ�|/�й¾uv/��j�n�(�%�Ԣդch` }�Ǜ��nxů.��EQqE���jB�I���W���Z�J�o]�;$�*{����CI;Tb�6�Y����n|t�&���e���	6�rR��]8D��tr��Mlٌ��Ȟ�̉[���>X�]8��0���h��Ƈ�6)l�h�c��N�4:;�[�(u��ӧ���eg�<��J {Ž�87ɲ�'̈́wH�t(b������$m��R9o"�����V$�N!](Lb����vU/nm��(���y%����� ��:^p�[G�~�,��}@]߾�6���q-��o�Z*	���P����[��xG��U�l�|g���w�yD��S��g����h����g��O���y�M���xJ�y������� �^�OP�+��֠����?8d1�̫{e:���4�GwO�R�K�kwے��J�;J���ı��N3Tc=(\�`��*i�A�60� &����>l
�Y��H�sr=F�zGv�ܩUhӭNŖ8z�>#�'ɲ5Y'�r��B�%K�c_J�4�ׁ���p��{�Eyy�9�`!�4�=���dގT_�n��M�l��GW�E60;�J����"�5'��}��IN3E�M��P��{�!�vIp����-bN�۝��ww猵s.�ki�i�ȟ��:>w�����&8c;U���� QÙm����p�
a�w	�a��w��m�
g�Y������� ����y��
%#2�<vvrC� �E0�K�����sl���UUj�W@)�vg���X�c	�"l�P������F^@�讀�#��LK�&�*
���jଐDچ�#����if.'e�qW��� b�UW� B�*}u�v$�����>�J}���H�:�H�&=0 �ҹw㑪J�,�v��k �pj�/�<!OL���b�U��/�4Sj�ru�/�x�.CZ���4{?��A����O���F��/����o��C@�>Za6�%d�pIG�1ɲ�X��:�lp%�F��ٞ�h�f
�h�x�S�@-b���΋ؓ�X�H2ͧ� nǲM0 Q>e�4�$ڍ
�Y� ��M�t��<�GDLC��l�P�8G��D���o��0��0��=�Q�l�T�P|>;�h�����&��[Ԕ��s؝،wh�'�f[�����w�IȈP��ِD�!J�������b,�>�j�P)w��H�������D"��Cd^:W[��#�o�-�n��vܤl�$�����)A}�xd�^��G����837Cm(�i�ng0?	�&�����߿�XJ��	t���~p��CL@��e�c%�?����ʠ�
e���_�̝�3m����ܰ7��dv-�G�&��W��&X*wy����aO>DM�d^p0�5��������nn1�������j�E@`���S$���.���l�A��˙�?��0�X�j^������-�Y�xJ�Ib���5߼�x������*����3)+rL�.�I~�B:�	��L]Y���ə��&fT?�*R�d�L����~����1c.���g{gj�^{��}EHU�
4&iR>��&�I99s�eg��4wLJ:��y�G=X����N*oH�luEᘋ>�2v��544���~�(� >����O#������,Cp��gL����I0�+2D����J���6g�߷��B~���x-���5�����!�����i�S���uC"�I���}Uw7��P����vA$}��� /����4�s�_�wƆ���<0���9 ��;֏9p��[�+��(�h����B.�z�����ǆ�Q���(�4�[Q�PN� �T�Rv��ٷʗS	��	*Z��$����y}l�݂�:ʊ���w�| �	*䎥�aح�K"z�a�gv�ڪ(�[G*��}��%V�p�rގN-��\��ԡ+������>�1.�L��r���2ϋ����CR	ް��)2S��y�[Eڴ��J�3��"B55y�%���䤯�h��f?C����ȁr{5Xɬ�.���:�(�谎�m�ȵ������ޫ���vS�w��0�������S��,�!zoA�[�}߽��$d
U��xbw
���8�=�TH���$К�ן��O�L�M�ٔ������������H��npz�g��@�c�6�����pYi��3��2젍��٢47w���u)	�g�u���ű���;�`��=x� KO��  �[ &}6[�n���gO��e^.�	���H�]�o�[�K�y�GK�N�|���c9�Y1= ��'�ڽ�yV�����%��9�؈�ޅ��}�&���C܌I��l}�Id��gH18�
<�t��(@�]Q��*Y�O>9�%��M��W������b���a�y����)�7k�C�0��&�G|Ua�X�q�����4I"�/5c��;�Q�
�h����%,R�c�g�b�*N과��XW���n36ց������H�j'Z�w6d�l4q#����m��Z� ^H�k֒ڱ;s�\VMn�ԋό��������F`1ѥd�����{�&�.l��i�V��ZEh��b�VT�jP0� �ZE�wd	`m5*�c"�H�"��Q$�f�5��v�g����������=�̜9s�u��9#�@�9�v���f�%}��)Df#��Hrr� cΜ�3U7�̈^����q� ط�=��]��w�0����������o_b�;�`���3(���b�;�'$�!��m~8�o9�_**`�*�&j+��v Ӕ�&Վ�Ĩ"�!ܵ�$�'��6�8��ޣ�����e����0N��0�3��Uށh#�\&����I0�6!���/h��nh<��'������l'���K�ХE�΂%�������5^[��x��ң��޷��e<�R_8GO�E|�&EJ�H�����\��]8���`�G@|c�A����hFrr��y6��W�--%��dJ}�c�XQ7�����(P
m���JB��@1�Py{��vrBlu�%��*"{�`�~��k���Ϛ�,��N���5^��3����
P�"��*i
{Qjo������2��g�I�n�u�}3���V��sk���˪ox����������r$EJ��N�P	*n��+S�V��@_�.�����F�s�:$/ �I�<�&��"U�ª()ciN��%;�l�#�&]�n��#�'���'���v�i4�gnT5�#�5.�)09��.�s)Jp|?�sW����מ�?&W��/OϾ	UM�{23X3�n�����F3��'��1$��OЈ���&�SH��A�m�P$i6���(i�!��!�H$��fS�MU>����~��:i'�dP{��Q�;xgiZ�F������ �q� �,G�Scig��<e��ʂ�(d�P���c���Rv���s�hт��N��3���L¡I΃Ѥ�i9}�gm+�������Q[�9a�=�g89"��r�����a+#U�t!��
�]���kd��>3�.��b��mB\��2�R�Wi'�H:O��!z���5yL6t�PD/�R��ђq����Qڦc�A����ZM��}� º�����r,��࿲���_�EhB�4ىft��R�g���V�����$\��L�P(��s�����顙0А��A��Z�s�x�_;,}�p�#�Ng�d0R�<��G�L
u����L��4��Q�(~������5,c����3�.I���Y�W^U���DJ�!�Ti�M0����qW�(���Gz�Ǝ!T�������H6��>}褱	� �f��$������k.�&Q�`ux��)�I�N0��76��ji����(�k�nE���6h�����a�M89�v���[�=[�L6,�:�.�_��ρe��ϋ�wf�v�{���S:v3M�^���@��[Q�i4zmMvv��ׅ�U�}����G���6����Ȕ�i�F3���&�lP�d5�hB���1Q���@��|�_�>-�>��i�
��4�K�+g�0�={rBՊ8u�i�p{��>���ٽ�`:~�Z��0�d�Z$}~�z�_�V�15��G���$�3ډc 'V�
g����3��6�'�\*aG��=��6����?�Q�-���Ԟ��(狒r r���#&2���srD��-.qw��2�?J�]��y�\
S�w��?�ZwH�H�pwt��I_6�B�W���/�O�|�N���� e����F�Ψ���Y�/p��`?g�[�u�J��f���F�8����+��-T^$�]����7\�/ٽ�"��˷(4�wTY��l���\�#	:�$����'��
�׷���W�[�$%ŕ��e,�	����N�KRS�|M&�rX�DY� �ګg@0V����T*P���7>2��R�%l���u�JC�b����"�nڔ��f�v���=@���[И�;Ś�mK���y�t�K�hI�#���Zle�S'��c����b����e�'}��ͣ/�o��i6>�1�2�`y�9�-�]1��'ڡׯ�٩�.���͠�W�� JDV|���]濷����)8<T,m���P�Oh>��T�v�b�u��^���
 �v�^��"�G�;�^=L�ܹ'ΟۅXd�<�L�.�)�)� �FAC�|10�P}[�f�C��o�4H��@��bT@;�k�A�Zy��Lz����jm���$�G0�[Az8�x=���7~��hl���Xj�����9s�oV/�@mt���*?���8�������Nm"�|hvE���ʌ���k��i��]�����wQGm�溞-����Ў!_`lB%�,��+�f�WO��w�P1��^pa�
�'�&��,̸�ͷ!�0��6���T�����E�eg�&���c1�Z�Y�5���`�C��
z�A ��UF�@S1���vts�,
��x599y�6z�D����+{��W=s��Ɠ� ���'��9~��$�_F�HY�7wE��q�&c�n������o��So����V#)�j�6X�����OB��e�����C���_�ĩ+��%�f�yF�U�2:�7L>{��
�.�N���E��'�)�IЙ�OORV�A_{܋|�n�z��ҳ�1���
"��j���opb�u���ޤ�|$9j /�н:e�r����g^�5�j�x�)\�P|R-��)(zA^Y��z�=���=�(Fn���y�F���@!R�1���;c���s�z&�A{7хW+]I��|t�&�B����ȉk�0����G���F�m	zf�l�b:�'n��������?5��%;cGJ}��
C�2���w�R��c�zc��<�\q��˝
/��EϑH=� ��>��$_��b��U��"��=�%u� zK�r�����|���#7ZVD"��h�e7'�	[��&δ����F��{�7ZL��w�S�W�Yc���v�$���eŶ�[F2���-��v�$�j��;/hK�Qq����T�d��1T�|������S}��G2�s�`��	�2�>h1p�6��q��\怊�}v��m����w��kvƹ,V�l�c\�f�֚	8��6�ǁ_���Q�|�4�	�����1�4�G��1�x��B���XT�#Fu�mnvvkqP���~�t��pQ���:�<|�����J�aQt1(�F#�|�Ntz=�l���ME`�W,c[V�]��jYAE*w	��k��7�k����,���%�����f"�,c���ٮ�U&�В�~3�d=��S�0ǝd(��=;++r4PG,Y����5�����$�
N�o,��Y�]�Z
>�j7ٻw�YiA�Hc�IR���o�@�O���:�8�<z?o��?��ӹ�Bq�E�Q��;��;b�zS�p7m����-�Q�n������Ro����jI��4��`�M���e�/��d�[��P:J�� ^��KO���|�FјP�Vw�/����M�+S�-a�K4Cd�ʾxp�j�4ש�(C�v�9�{{�N'�Zf��J�����P���o��%c��̪�\����)a	r����J�$/��>xj?H�"N{e5�����5�n���������[TtI���g��dtS�v�q$m6�f��y�1d���M���GGTӝ��!���Ior��`x�e�O�y�˚WVZ����P��;�D�w��6�	������AE�S(��fy4&�-�s+~0i賋v�$,D���9W�i ��~cr&I`@��2H�]���W�2��$'����3�l0�g���qⱱ���(���6i�-�J�ߌ�����9����tA]��|J�r�ʃ?*A������'���ׅ���k��5�զ���V�f����V���I�lC��l�z4�Y�b�4(�7�%�����!������8:��P��6[^z�&}-�I����j� ��2.nu* ���l���ǣ��Ue����,�7_f�ay�b�����,/���?�D�K�Jp>>����[��آ�b��Ng�w6>7��{�ԗq�X���N��4p���rמ�֟p₂&�6EPb�6���!s�X�.�J�C�܃�<�I�N�kZco��" �@�of�PW�Ůx~�D�ќkX�|�r�O�w4n��3��R��y�^���Pr��k|�A՛v�e{��0I~�.� Ѝ)�$�����[ڏ ce���nJ}��ݑe�-O�4��\M��쬃A�w[����A�܅���j,@���dM��d  �7��<���pIد��*���1��4�9��4���>~U�I��,a�&E��C�F`���Z�sK�L	e(V�b�W`YPp����ha6��|m��Zx�ϾS�B�aM'���-�<"�D���_��|k,Sf���t�hl�e�;��#�×fK��z�H��9���Dv�(���a���!�V���&6um"�]U���O�w�:���v��w�|�h7]�����}"��{:t_�B�}��a[���&RZYYr��I�=C����������kRc�{�ћǳ����h���SȯPk��Z��t%M�B��o������dsFU3ܖ�Y�І���'
&�g�.]�4u�SV���6���.׏~�Vs�������l��S�'�X��d��ԯ\��[�#��K�2�z<4�J.q��0t:F+�N��+��ܞs��z�;���=;-:�� �)���ɔ�m�@3�/C�3��#�z���a��E&~�5�]��	|@�iY��U�����=CX^2�0�0yP6�4vj�QF-��phh�N���F8x�����Ռlc V��#�NI��s����=���810�\��(3�. (K�q#J�[f�b�kj$���6:Z�ň�L����oR}	�\?�͋����\X3T�?{�æA�7�=���It�/���y�q��uw
H��E�|��N`T�٣x6��_�	���^����-�հ'�m{`��u�itd{	Zᶼ ��ǵ�_�R�]�&�Q"�y����d\8�����~0Mea���+%AzD����R����wNz�#����l2�{�C�+;�w5��3���z��@G��O�\4�^��uB�'=����Ğ���VٓU�&�<���D��m��B�>cZ�<젊+݋tmK5���i9}>=�d��qb�9����|QR����Wͼ�i�HX�-�kc���t����֑���c����Zg͵�gt�q�[�p�'����B��?�^����I���6.v��	�������:����l��c�e���J�Ϗ|����w����믵�߷R"�j��������R�r�;i���	��l[�����W�~���s4I�N��?���	�iW��J�넁�����[W�����
��(I/�;�������/��6[�Я�{���L}�y*{�g�4G7�^v0ב�g��dd�p�������u$��P��(�R��٘#xǈ� ǯm�QK��]��\Z�(�j� �k�Х�uw7A����hWϰ+ʞwzD���D��I���a[T!U�qo�H�l���Ku�KI�#kTqڃ���i�8�"D�j�I�ه��pk���9i�F�tE--)���vbR�� �@�B��p�w��e�$6~��x<�2)�?�1��ޣ�;�d%R��q�+k���81'G�H�Y��(N���/r��O�{N���\����)���
ԟ���]3��F� ��xa�Y,O9��oG������u�*_M�,ҿ�6���Ɉ"���V����5�"���.N�95GJ2~�'��%����5M�a�)Btu�1xug�YC��8��=:�T?����/�9'���ᰗK͝)�'�"d��r�ѣ��5 ��`	*w-lA+�k����XZ�y�6�M�l���Df	��s���qR�j�oܶ���H�����O�`��c�/��S\2E*A)�_��=��}��� ~�̈́��_]���{t!�ڵt�i~P�V��jM����C]�8�&2�)F{ʋT�}E!M�
i�e]/�o3�eܹ�������Ao#�R����S(�9���R#??��5�P�o��!����T���ݏ���[�2�g�]�K�2y�t
\�ՁT!B��Y{�i���Z���b��1TIބaɉ�eכ�xL��s���7��(e@�q�F�L��G�S�<j�F)�qX�^+�Rf/wNN΍�(��r���̠��8-;NW�9��C�{g0.�tdw|��΍�r_=��<�8H] /�h�'={�,�ʲš��ăS*����+��}��di�����%�}�H+��;"���MԻ���eO{�[����Q�*aMlz����-:+�!ﲲ/�朳g�j� N��A�G�c/^����S�j�����kϓ[ՠr{rbUuu�Mn1�?~�NkkS"A��)���C娠M��4;1K�8=_��ò��C��^~%����K��K�^�c>�Ӝx_���"���{(�_OHH��o+��/����)���վ�oBH�!��'(����}��J|jY��� 1�3̨�gQ�1��N�f֏{�װ�#=���?��is1��j�PoM����`0J~���*����NlH�*�@�
๢�fU>B�g��q�&��\�LE���d�NKI�9
]P�b�-����$qR�D�����Ν�N�byGS=���Է+����I�"KFd5�����l�gK,=�2�3L�؊3K�,1s�����:����	)W�8�xf�F�e�K��pb��;���y�y���kkku��Q��b�F�K3Dx{ߥL$�ޏ'U[4.<�]��s;lG-n�X�v�4E�J�J�_��wh��`��Pڡ�ە*�ʧ���x��8j�$uF��k��7��,n����Mz�\��w��^fy''L�-C��&��'���=7�)��zm9;p��꽀��,Au�ͣ3���q���п�y��{���:/��2#��(M�`�I�V;��K�)�wPϳ����9[���R_��)	���87֝*ڥ�v5M� s8�1sz�l�I���4Z#:�^���&��4��	4��1��ǩjX�:"�k��ÞX��"��Wi�;0T~G�L��8�L�E�<`~�]�a�Ϳ�4;�X�q����z�#v�)�R�eo��j��@�?~r.)�g�C[��1+W�^��P�����U*a]U��.�H�a*X^��`�,P�[�(B���WJP�ӉN�LT�?*Sm)��!�k5ˣN|Z�z�\�\�5�W��35�� E�~��cn�.R�-���c`�Y5�6�����rS�q�@Pn�n��[�	n�;F�����������T�h<���)���1����&;;�p�u��.KB�]D��z�h�2�+��l#�=7_)&xt�n��-Y..�ArU����h�,5x�����gT�w�*������07*̇z
�{����&X�J�j�
dm��Qsl�i���)�a
8k�9Ok8� 2,�>�Un���OE���-�a������
��]��e9ob����#��FiV^1R���FuG&�JQk����e�6�B=��W��K��)R{�PC�w|���j�IH��Iډ�r����
&�)�R�4+(|��
̜L�n&=%
�p��j��T�w8L0����,�Ȥ�����æ����&����j�/����4vI��gX�����r�����+�~�LRv��'	T���3��o��M��b6DT�ߤ;��GmK9�Z.2�=F�x��1�����;��j���0��W��øW�F�?~$ع�^.�q�y������i�/��w���n�f[�ɉ��Z���sy8������>��PU�]K�,�yn4c��GyH�7����ן��Ŗa8�?��rM�z�Ldf�����Q������t#(�=��ۋ̓��]KG�:��h��K����!:�y����|��/��j�Q�Pߢ�qp�)C��8C-��՘�5l�=���ť7���؆Ov�o����a�~�P)~к�p>fX����Wn�ԗ@w�C�J�᷵�����`M�-S�x�P]���{9f�]%��C*�����4��E����䞻.��ˉ�bi�m����=G۔��@|*Df�9����Dp��8W�39�%x~��j'� NS�3��P?�n^� ��]�n�Å��[&s{zz*����=l��M���ua�H������b��������Ä�1��jPxc��|��keeU^Тmz�K�G�*�6n�3?�CG����C	��2b��ݬi�%K���:fpp�F
������2��_}����2���܌����6�D�Ʈ�������u)��p�ۣ����TbS�C�w`HJ4������҅,����.�
ޜ� /�|T��&�ʬ��=�׷UG]+P��v�FR�Ě&!�Ѥ�~�<�N<_'�6'!�
��۹��D�&���Y�%�ۂ�}E��jh�3��wU����а�̅�y����շ�3R��TD��^�	<|�l����-�H-�F�U�ɘ�Ga��D�L���ǔ��բ�/Ӵ��''�o;��?��i�h�KwN�U4A3���J�9�H~���D1�������;l��8G�vvt�M1�K���
��k�q�8��f'����\�ɥꨥ+�zY�^SE]- �4y(q/w����Σ��Ē%�&j���<@������.V���N�^_��m�����џ�S���6�/�qٕF����LyMU/^���B��Ǭ�PQwQ5����b�B;rt�Ƿ���P�PĒ2lS��i�t�>�P�&����gYq+��J̺о�������b�����;�TFB�Iӳ�>�[G���i�·�'�Wr{A�����ёÔ�P�7�f�{}p��_���[�F�-*
���gi��](�*����Ѧ�(A�&���L�]���g8�q�����d�:�
J�-�ˬ��n�)��{%L��wP{���;h�=ٶ�{;���Pv����4x6V:ՀDrW��ޣG6����0��_�P��p<{�<5%%e�|��Z������?��D���>��ZD�W�ķo�������9v�w}]]]b�\҄e��m��F9Z��x��+��z`�k*��j�L�tmѢE����mkg����5	��*Bg���ۛ�
'�&;����袋���ۓ��+��"��Z�>�I��G+�cnX��m^�F0�ǅ�u+%�`��>m�cv�F �� �s�_g�����P��/$ͳ�yS(�r#Н}~-���4���W�v�Ƒ��Ѿ�*jHi�,A'�e�nhiiy�S���L�+D��(0G��)��ç����_���L���uǣ��B���M`�a<c���h.�1��|�u�A0�"�x���l�K�@���k��?�b�Bᙆj?v/����]��=!�{���k�O���
}������O�-Ɖi��0�a�6������v���P4iIQ�P<�Bn���CGe�m��,���跽��pr���=���pGTc�Ytx���*�q����@{AX�i��	�6�a���x�G뀹 q���NW�T��[�λL&�I1���Y���3!'��6���R��5�����V �6�L�j�`6y+���oVo<�Z��=�X�*����Y+���ݐ+���i+�ş���?/5}��ZX��y$�dDz;�����t@x8������=�fK�v��'��3;�T �X���`r���0[n˽����Ѹ9���PG�Q'��pb���	j�i3�F���^{2�|�*_���}�����h|�<ɥ�ܝ9G{ui���
<�Y1�5/=
�L������G�����D�Ip�&�8,}s����|Ƹ�{�⅁=Y�6Hns��EY�N�k�-�8i��"=<<z��
���k6��X�^ؠ�T��/�@�#�gͦ�*�Ha:bo=~����2�*И���w�;����9������0�#���0�'���)+o�rz�>�Wm��t�x
��t�g1���j}�|go����B
E��<�ϱ'{�ǻ���J}EުX,]��V�~uv�#Ϊ�)Y���q�Wc��ms_���G�Nha�@&�6���/�-�cy�׬��?#׋�=ϛ_8T��df]]��.��&:�1��|bMW_|�,n����z��YV��`G�d����C����@#���b[����ڛO���&���b������b�w�!�o`J%����-h*J�Ԗ����F��+��Vvdpr���z�Oj,��^ۊ&pL�9����LF`Y���t�l�3b�ŭ�Ǌ��� ,��7gԴ��R;��Č|Б�:̠�V��Rm����4�h�'���O�X!M\��EI����m<=�lVTT�g|�E(��� ���Z��'���/��%K�?���P�`���y��J`��P9���9�����s��|;�?�;�����=�� ���f"��b-ŭQ�R89����ϖx-p��ĝ���Y��ܟ����xo�n�I�/;��sŘ���6:�*6R�Ȏ>���
��&��  �iȉ�s��Z�ٸ�yI;���ϸ[K�5{M{�ex��Q4{gʰ`���џb��n�6��/c�`
��k�8���k魖Ԁ�V��%u���;wN��3ρPZ{�$/�l�>L�9I�oK.��E-Lݠ�ad��<L��l��<|�T67��$��Q�y#���§���+	Zi�a�i�`n�ɲ�8�E�Xe4����1������b�l����f��+��9o�Im%�t�;��sV霞�>�C;b��J#���R�V,���FN߀����0^k�*6��|<4���D9Ys�O��׌ˣ�LJJr�ǡ��;�`[\K� 0��)1.(��*���l�x�7ʻ�m D{{	֝��woK��[r�x�B�}�?��ݔ�27��o���u�eRɱ�2��^�T�P��I���9zͻ��]=�6�KsuqBqD����`�\�}U��3񋮈�K���2V��l�)6b�8���`���=A:`���u_�ፍ)ԕ��`���Z�����F�C_��O�Yl%�l����o�x�I%hI��e�����~�H��������c'm-�5�̀��+o��~%.c���q������)l���,��;� �@y������*Q�x<�� ��g���+]�M ��D�ں���궽Z��S�zl�C��<b4fG>4\�_��(����]�3K(��%^����䈈��_ P�Q0��C"�����Ntp���3��;��޹{t��2?K�t�W��ȼ�d�z?�W��o�]2w�#	7��/�%E^�emO�=�B��l�g�e���)�K�����!Ul������@Ƀ%�����*�ջ	%Y�X�u��[�=�gke(��T������/F��6��c�N|�Nu<8�t{�o'ձ}��Z+t��;E��ݐ_����=O=t�sk��1�����3���Ǐ�,*P�]���)v?Cc���K�<d��������$Hr�2v��bq�3�iJ1��%<L��h?3rE����p�JTn�@�;��./�k�IA�ԏ��'�3��"�l��yT$�Z^C�i�y�8`cY1��#������P��Qzu��='��4B�y�t�����B�^�0M���F�@�'mR�L�s5�I�Tu��+�u^E�؉y� ��%��G�`n=���c
)��U�s�]'��H�s}�"fNF��W��s����H1�����r=ˊ3����V�t�r��4�zk�RΣ �X(�H�={�����G���1�	hid;o�
:�n������|��U�bp�<x�jϷ�P��'�)�����|��X�599���ܤ^���Q�.����@�-}���~!��"]��x�,��w]�D��ǯ
P�A�9��\��o��q).�y胋9dG��7}\��E��� �������6�h6�q�$q�2�u�v'*4ŝ���Pf�����^r[��������s0Al>
��k3�+��5"�t��qc"�A����w���GЭ�&���8���I[���M�'��ryoAy���(jr�gZ�-`���Өi�^e�9��
x��h�`��M�g��?���Fr����XUU�}�>}�	oJE(�V��	�����Ɂ����զ���*q�%�EK�`�t�K+�t�l��է��ES�8����B~!�ϟ]������_Yi$pP��c���)��mR����3�"V�I��xp�>0њ�1��ah���ϡ�-�`nE��Uل�<����$�#y�)�a>�~'*�+/
��k�(Ut*�&���Ln(��W��e���0�fZ��3��=���ς2]�ɕ� j���\!��g�c*�IoNA%S��5lE�Kn<f���_�C�?O�����光�:��U$^TԏGנ�K���	���4Cg�Fv4!Ŋ�9�hB�d)Ȟ�(��(�+���T,nĴy,d�$Q��@��CI�L5�6�/��8�.^Ψ	���#���F�t���A]`H��~ؖB�YO�F`�����]8�GF���j��c�����9�5y��ц�W�Z#&��T�)����S�U>R��KD�;�Ӌ�8�v|@Q���Τ��H@�A@֕F��>>>
?��ʇ�'�vɟ�Al5]�np\����$�@j�����?��PLe߃�ܢע����[f$��*87��V	�҄~x=��d���=?�1YG+�����i&�ŉ#��1w��F�I�����+�K�Ĝڟ'_���������ׇ��޶�qD����EƗFk���F�c�yz?Q���/���ԑ�yU�9f�),��	�S&^�%�V��G��xc`�g?�k�&z��*�A����O]�3�6C�jb�A����U�ip]���I�hXz%�7���L#</+�7��	~d_ҕ+��s^���ٳ�խ�&��{��S��)�y܃���bH=ѥ�
-�x�'�`�WQ�3�C&
�֟�#o�샹�9��+�a�Z)D� �?x�-ԭ^��\���ӂ #!���'�x&;HL����cHC|�(g�����
�]9����4v:R�!21�T��1����7�o�p�O�,5]�cH�CF����+D����݃��l��r�"�����F�"o��#q>7*�T�\�j���>���M������<��p�3��>��P�(}�OԞ�Ss���鋘#b��� �15n�'��f?N�k~�y����g�'��e�&S�2H��\���Fg�ũ�F9?�>�)Zh���~����C�F������מ�v��ݮߎW�~��M����J�1�vd��K)��b��J{�.h+V�"F{;T_<96>}��u-��zf[���RAR�cG��Us@�|�=ƺ5���ظk��eL���M	_�E�J�
�Ƕ�~���L�>�עd�7k�.��~����S���C����:���΄+c��R�E�}|�h����䪢�M�m�#�W���w�u��T�e�o�q;�̎hL��1ǛB=�kL�������7��"D/3�b�>�T�����o�Y~A۲��ի��״Y8�5�tn��ez�O�_a��ϷscmV��zj��έѐ4��V4�1,��6����J�~'�AOӬ�:J���A�����N�MD��K�0����yO��j$.�9Dl��I��s��H_�q�����o��[�߂�����-�o��W�(#E�/�>��&b� ��ض�^��l�?JVXǗ��{̛�܌�u�:P>��?�%�Ss���?�Z0��*����|9わ�-�4?�S֊���,��IN�/�~/�\�Tzkjk|��� ���I^Ôյ�V�,�q�ȻK��f�2 ���I�J��>���d�" ߒ:� ��'�qs���~����"�-���B3Y�Z��d58d9�ø����x�x�{�d���/W��≀}�OѴ4��v�{�bɃ�͘<(�Y�)}WY__/�	������)nm��ƺ|��r�ѡ�ݒ�w�Ļٿ=��������+��3^RJ�Fe���>n]7|�#��BM�;^�,-i����ۧ����&{��,9���Fʋ��UC���Ii+^$����ٱ�بe�]P��-V��J�jvh�z�,��l~2547Hn����K R��fk���ō�o���8�m� |��E�ր�����*�l(�`�#�~��G��\;w{��E.�]\���e��5�^^�@����D�<1�.���\�^D̀C��rڬK�=f����=��`�&��H�G1��YUq��W�VWWo�e�}��Bf����^4�}r>p`t�$KBd룏����0�$<"��R���䫇�ۥ�?�J�*W������p�_|)����1�އ}�?���|����E���}�c�)����?PK   �n�X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   �m�X�,͓�u  sx  /   images/aced3900-1e1c-42d2-9dab-094da686c0f5.jpg��uT���9��@���w�%�Cpww'@pw	������=��|g���޻�o��WU���tu���m�m�^VRF 0�wޖ_ ���i��_CBEBBDDBGAAF�D���@�����}��������=�<|||�w�DxD�x�x�y¿{�А���0�������
Gg� G�ǁC��{�P  pHp���-�����߀�� x8xD����_��~ "�G1�*�(T�x���<Tj�|�?4\&NAh��D�$�t���yx���|������U�������cjfnaiem���������=$4�GxD|BbRrJjZ����¢��_�u��M�-��}��C�#��3�s��K�ͭ�ݽ��ã˫�7�w����@����?���<"""�|����g "�Gd\1c�T���x�м�4j.�|�?�4ܛ�����_�����r���?|� �p�^@��3���Y�V z��G��O�9����>c,}�,v}!�����^���O����^���
l5Um/�*gFͮL$O%�ƈ�f�h2)�#9��B#��C� �B,���dl*���9�?���1rR�+�:������>�@��S�~T>�ӯ�{�}�9�;���H�e��S���>��
\ݯd-�<�@�zꏚ�]{��x�
?�g����g�K�W��>���^1rI���wi���Q�L�N,���S~�(_b6�f���?�k���MG�0wc8ń��ȩb|in�u��X��*^=2�vp�*B{�k�=/I�z�׬IB��2�f��t�������0����$�vl�v(�� ��|����Tf��C�\��#�}��S�|6�4!N�ġ���y�<.L�c��M��kW�����G�3���Շ 2A2�ٙ�pVo �
�y2���eJ�/2��a��q�x�RtT��'6m�gx"S�6̞Z���,��.k��b���m��t')7r��|/ip�Ɨ;��y�z�}��$Kw�_rE�-g� m�!M�t��v��a�RLv�@�¦L���q+���/L�l!��|턘	tEţ,�i�b�1�1�F��+L1EY�~�d.�n�/��G���|j�\�#8SK�Aj�S?���[�fݳ��x��r�Hx*��j@PӮ�U���I��TpYk�h���{�_�����Nr�Cc��a��n.��g!��������1���J��8k������c<�7�k��f��>�e���m[��RM׈̸&:bi�M]�޻�{R������=h��-��9��!�;���F���mw�Gf/ׂ&��lM�Z��az���"rVO������F��:q����Z(��t�=���KF^�y@�k����4��	��X��@�B�AA�dU'/����� 2ﾦ��h�8m����_��� �R=#D���kI[�|:<�VM��C�H�M�&-���ߝk��x�F�>�>Iq�m��ݦH_����P��͗�F}��]�$����aއ��-����-�gXR9]$����q�I�0!��p7\θ:ә;���uY��v��V&ؒJ<=�jV�����b7Iw�g�?���/5��
���re�(R�c,m�+��eX������a��!�H�y���ڡN��f�j��s:�����aX���H�	F���.բ�Ck0�,�̉��S>;ۇ�����5��y+�2u%a�%�lD���1��ދ�����̨�Mv6��(���ֶ?IK��iۓ�1����v�������
�OS�^��Uw�=ɫ�cĹfb�\�_Y�B6�hO4���i�@Qu����Aиn�8��2SR�b��Ah�T�����,�J� G���>4&�/_�?l{�N��u��sJa>+'S#
���56�@v�I�iq��ҩ�p�d�2��%��؎�f��QE�k\|O�H��Wr>YfӼ;�}� �S��j�}�{��ߓH���8��d/�l��+�	�b��B�_�nٷ�걼 ��G<T�wI��R��]�7��g��̈́ٽ��DG?�;FC�J�'Ӂ��7@�Pd'Y���R��:�Ll��kN	�8��?�6F����vąR�H�~�/S�b��]�74��ള&3D&|�]��n���dnWJ��^�!���3�Y�15e:^�/���!��_~�fn��|yG����NO7%=i�A�J�i~��Cn����߇���K���K�}g���/��(U�Y9�ݾ6���"]=miT�dA�c��Z�,�2-�Q����C�]����B#�:G�d�$+�Q
>�~�8fE��5�.1��D�Owkg�����6��>�f�*�F�6M���V#�E<k���[T���Uzײe�)B]����y�-M��M>����0M#�hO>�j]�bbO��6l�:ϰ�H\����j�1�V�R��������k�7�}����̟
������ɕ0q�}��*۵mg2��z|h��lu�m�.��.p�K'Eqڌv��m�W�+.(϶3�/�>.͹���N��F8M�/������P[=q�k�ʙZ�Eg����3m���Vm=ɿ�N]���]���}���y�b��kU{=�������J0����E��	=!!y*���(ђv�u����N����<z�Q�r�V�CP���8w|�=V��w��2�[l����Y�]��U�=����k�y�e>�ģ�� �}o�����b�����9����=��+Q쪒��Y���͏x��'��v���6w�k��'����8\��E�]��*!�����ڇ�K,{Ʌo ��"�p_
j*�/.Y��D���)�U�~5������[d�\�^�M�4!�6|^�1�9x�.uQ��� 9��nbۿ�6-}�z��H<7'q��NVx��B��{G���mG����JO������*��;�S&͎*��G.
uΚ�@����\z�)Wvϥ�:뱑8��äM�7�-})�|�f�R-PAW�y�#�n?�)6K�@�̩�9K^��p@-aGTb2�GH_N>kP�����Ed��3C�F��N�'QqeBv��dG��O�]&�hf��߭��uf��+�����e�ˠܥ�V���MYV�S��{����.�0�J�<V�v�ř��ŋ��E�+��#���SQ�se�a�a3e<������zt�D�����0t�h;�ڛ�����uhM�8Q�%]^�&`i��\�Ǎ^�h�o{�5���S� �ⴘ����ӓ�����De����Ñ�?�˛��:���W�ܻ"��0��V>�V�V_��(*_��<ý���[G#��q&�ZWk��!�\"2Mզ���@��ZB���m	�~��kKf).b�Q]�3�����N�1� 6J��B�M:m�K�^kv@)�����"�>�=׷6���^1���Y�D�KI�)ꩌ�c��I�֙� ��;!"�w:7�<ų��`W�YV=�w
�����������O��W���	�s�gC_ҥ��(�A���ː����;�U�?�\`S��YK�]g��*}зtbdU�E��12ۋ��7 K%��� C˿��,�B����E�m�H_�	o��Xj�e W���D���DY��\� }��H�]��L��>S/d8ކ�Җ�?���u�!��U���a3�St5�XpQ���3TB��!a��`E�"���Q�ܬ��9�4�
U�'i v���C{e�`�vV��̩!��=���?�E�=����)p$u;﯁?��cd�o���'��?	�[��i?��7�}UJsY���y#�Ҍ%ҿ\���{�3Q�&m֖<�K�kJ��cX)��v��d�+�i�!"�b2�YE#���2��Nijen4��J�[��2^*D��lˋ̶��dA\�9$�)Y.B����q��X#,'M����7V�;>��Y@?�j@W���Fk/���s�8���5��������0�uI�u��d�@�n�8Pt���ڃ�JѺ���~1��Wf�mؖ��M��߶�6��*0?���Z��B�Һ]�$[;���{t��8�"�"��n��}Jsgl��$@	�*�}7�[MR���3��e�&��,�"blPǮ���q�vU��R�?��cm���s�r�Mr�fJk�<��k��i�h�̂�+H �)�7�&��������4��&�)� ��Y^���=j�^f�%�T��^�|�}�Nܡ J��ϵh���w/	%Ø\��NCVD}~�t�yϝ��
�)��gz�$�?
b(�!�~���E���D�M9�1��1�r	Yg�ϭ�~������Ȼ�kV�zG{�3��e�(�R�q�5�f}��:��vB���G��R���QbhQx͟�G��ѷ�  �8�t�g������ѱ����
�b�\��Im�T�T �C�.�b�&�z�ࢲ�t��J'�Ǐ�J,��Uq��~�N6��D��j�~�9Z=�&�I��������9�|RHq�2&�B�7�(3HD��=~op�(�^ф!n��\���}bm�X�=��Wi��&n/n���pK��?B��5��/A�B����E�k�z[�\-^�ϋ��(�[�-@T��Ɂ��̖�U��4`N�w����<�-c�=CK����٠~yaH;�F�&U����ŋ`��2c\�?��M�t�Qi�IG�v�TT��`��m���o�$�b���1��F�P����$��k��%��,��;DpO
�[����Â�!Q����$���g�E�s�/q���h�`�a��T�o+u�W�w���?��L>����|јȧ�����J��	�
uU+\�&����6��<�*��|��̫I(y�������?��V��]�7�7�>��2.Ϥ����=ކ?{CǞ��#�>?�_�Ĵ�X��,�z\F�g�F5�2��O	�?A���j�����G�o�"��6ٖ�6�͍�<���p�����V&��e12+��!-i�QP�Z&�^�oR���P�Jd~�W�<\+��O��P7�e` �N����Z�X�O�����������V�(CS�0TR˄�{f2h9x`L�Ccm��)��������c[��lw(ʮ��T�=ɀ��٤�tXT�� ���3J#w��з��,��կ�u��ȟ�	���
w��
E�]8�%j�,�кĆD8������AC.!AT-��\*���)��y��J�ey6����gM,�ĐyĹ��
����}����2
��;�ma)�W_f'����w��.�I�ޅ� ��'�5����.e�y8���G&4̏�����h㷃���OgS�h�m�1g*X΍��|�<,uE�-|���=)�Z�Üi���d��`�>?��>> P�˪~Tcq�3�h��#V3qRW�lz�`����r��/Rw.<RFs���;�ND	�Y�[�:������Y���,c��F�3x�*��$@k��P�m���#oZȰ����S���T�[7��@]�!l4xoh�7[B��^� ޺�����Tj��Hx�yW&�>B}����LY�䍚m���]�!h�jȉd�I��l 7�#u�}���`��q�;Ye�JY+���
{]j��+[�2����d�w�7m"��:�#M#�\�'1��|���^�I�6��Џ|ެ��Hf�Ԫ��{%:�8hqxx��g��eu�x��)r���|��1��J�.D�#8��wf���	ӑ!�}���[�kt�f��t��J�8�w�A�hc.�L�h���?���N�Y��D&�}H�s��i�s�w��$+AC(Lx�:�P���'3Y Z�����Eh:2��~9I�Z&}4�م���}Yӟ�Q������"�~v�~Gjê�n�M��0Q1���&:[i�;�%ݨ�@o9Xw{G���i�s��6/)�������yju�Co6a�b='[�L�[v�+�h7�����l,��q��I$���O6l.c���~�I����K�Z����_���)�4�4n4O��V�O�#
�.���Xb'��ɑ�#Uf�<ɋ�-���W�L��������<9��:�)��e�[����B�]B]̑�4�%4Fh=#~��u҄��o��!t��
��,QFG�(��crr�|^}�1��1[ ��XL9;��t\�D�
�
�e�� .�,�$���GKNk�>S�*�H����(x�� ��x��GxB7��I+��}�=���]W�1��}���U~��Y�[���p����S�o��m,�G�)4������&'O��+L����f�B3R�A��W�p%��7����*Ũ9���dX���[{�
7����j�4Iд��E��ٶQW
v�oᳬ�X{�m=�7ڣE��[�ݟ�X���G�L����Jl�r�r��/wC��s�i;sJT���\�Y$VRi�(�Zgq�T�ͭb�,��k;�Z&�;��u�����R�n�`�-.�T���(l'��Z����T�,�U�7@�@	��B��c�e/�,<���HJ�>��A4nc�a!�Y�����@�Wa J�d�ˉ&��'�s�LV�\�!ËϷ�D�?,-��n2�X�rCI��4`�y�s��3R-3��
aQ�M��l�gE���#X���dB7���@�d�������U�M�E�ن�g��n x���#�P�xE�]覩t�2?sS�m��Sy�m�w 0�J{T�a�ZV�ML���m���KyU_�,CN��r!
r�`%��u@Va��0����x4B3���@ |��P`X��:��\|C��R�"��\z�""����3sx-����P,���D��P^�S
.c�Q"�\��}�׺��,�;���% XAkgs@��ܨ�H��!��J~�sɓ�P�X���YK��6񚝘6�@	b�@a�I��~�8j`��yb�Q�λ��3������Ex�ı��#���9�������+�K������,S���J���挒Ɔ� f����i���~��j��{��������ǛVT���F�af�MYe�b�����D�r��
4ac)ݼ�1i�'M�����",=#N�ԹD� ��ֳU,�p�$��]dE'���y+"�@���>N#�'?���r�٠���vYi��ؐ�|JӖ���pg�h�g�v��R�*Mmg�f�n�ڿ5*9e��
=�[&�\�ƕGO��~�@�t�?����y��7̻l+���ޘ|�̩՗tg��yK�ү��#�<{�ӑs��'�8C��X�����Aʉ� .¡˴J'A������;��1���(�)\�j�W��#��u�_n��TAL�Z#�������p����q�!��3n������zڻM' a6��k7�[V(���Y�%�0�蛣�2Ee�3���9ȏ䀺c��Nsj>&Пqy��֌�X	F�T��YO$�B�(y�?����Y�����+��`�Igs�<�;A�eS�4���p!��.~F�F�p@��˴�����z��g(�ۍݰ�I��ɴ="�*a���VkM�Q�AUQ�\����|爞�w�n`n[&��� 4�;~�%e�����V"��mB�.]�)��E�".C�0=�eJDj]޽*�"�L��
~8՗A����Chd���j�����H�KGz�&�49/�CMT�;��L��R���h~�o��Q&�N�\����M�P��(�����w�L�6�%[V�.��d��9o7��H�ѽ"yl��������/��#�ۼx���W�Ă�4��ĸd�HHi��p혹p��i� ����Q]�dOK������].E�tD�dӯ�}�0�Ć�,5^�Bh�A#>�2�QI�!��Sؕt���]$�?f��5�	�<^u���団�k%��@�������_���5�a۪i�0��&�oj{�OzG\z��T�(���(�o�`x��s�p�U��i����i6r��W	!��j�:oNh׃��f��zh�$1����K�1�� |N��Z��g�U�^��˽���ڥO�lm򂶟���]��c4_�*���(C�6��RX50�Ό>S�F㖒�շ�a����m��RmuFe ⧎	��[����e�\��a��u͜#��:#1E=���N6��������`�
�&���.��ЪX��MfDwM�|At?����5a�A�S_��~Ǣ���^�t�z��!�Qߣ��Ո.gL|�5����b#�2��~���xw�v�)t�'L��B�Z19zQq\���-&�n��g��R�e�i���b(��s�����q�wL�+��{���u��egWCc�	"���ϗ-r�ĨJup���c,�+�%3� ų<5�����o2���S��W(�)�S�g]���@�O:im��5�.^fg��m#�Ը�Z).�hr�äh$���t���X6�[�cـ�6��c�B��$
M#�������2�b�b7��G�һWS��-1�ޚ)@f�I�g�^O6)��|�SxT�ۥu��<�����'aF5��%�����휩��� �x@���U��R��T�p:�J�������T���du!��at�)�ҏ�k?��F;I1�6�m���GI	n���r��;���0�`���q�b���$ܰY���-_k`.����koܷp�D��VgM+�pP�,�`�*�J�{W��/-�SQl�J00�yJ���f��Ƌ���d"�-0^�72W�<��D�NR�s�t|#�������̤�4��uĥ�kW��D�D��{�~�9H+�0o{,�)����S�~	X��*�NfWP 8K��{�G7� ����v��r�W�3Vւ�0��bW}����i	�n_�Z�ρ��W;&6{e�E�CW���
�*�����K8�P}�ǧc����X�8�,R�����|��y�Y��rr8����?�'�R��kم͸d${`��BF-;�ؕy��L>�+��D��J��1v�Oа��kv�����-F�@���/�
�_�q�M�B�h��M_G���Y;�|����Tq%!��^��Snj+�]n��y�~ �cq�_�ZѶ@�r�I��2H*���)��7'��w���x�0�'�R�a�9�}���H6(���)�oq�T�K+�$��Sd/���]�,l��7@�O���Xq��P�iw5��%4c��d�[Gڹ�z�p٬�wVVw�z���e*��J�a���a6g٤�I K�#��w��D����p���Y�=^�!;ؗTb����`+ئP4��+�ajL�a2t[�q�tC�΁��?:� �7QP�Mqx��|̨X�'ʼD�ȧ��r?���33%Z���l��bLTox��h;P�8��<י���ȟ�J�Е*QحW坕��w`��ԗ@�����o�[7�ߤ^�Fsk�k��� l����@*�WШV�h�!���A%��I�&$�{�J���v������<V�ҿ�����ܑ�h��#+ۣ�-iܭѥ���KQ�yF��'���i��=����&����݂����j��C�S�F�G�z
�&�M��y�,�V�f�`V���>*}��H=V^�G�m�kw��3�����DM��#J�=C�!����\ c*
���}`*�X���29P	_KgU�$-u����@%��  @%0�ր,{��K,zbw�n�q��L|��� i}��a:��s	��8�U=G�����FYOg��&�=�k��$��+R�X�Y"�]U
k�84�����]C�=.~q�z�9IGG�\�*��$rP���k���{�����3r���O�3�o����`M�oU��V�ۃV��y��E��f��{�x��;�w��P'2P&2��������pm��i�Ӈ���Β��&)��S֛��>w<����;\���1���k/3¼����$b���b����ap�J+ލ��̇g+��I^����V �h�DY@�%Y�sR�P�H��?��D���`u�m.�Ȑ�B\Ʋ���!@�&H=<zZl�I��P%nq0�}a��p�V�����R&��	5�-w��T�[�����TXL�6�mƱ��q��m�[<��t����7'@� �AK��T��l}F�ߕ�ӭ��n��e'�F��r���&�ĮX��t�`z�mTB�Gm��H51���*J��7������=�TW�L7ɯ��
�*،03VT��x�j�cr��� o��F��ϟӆ����px����6}l3��<�gf�9/���:n��)[�����q2�J:���jl܎��!�z��c��U�m}^ݪ���1���\j��$��m8:M�  O���uR�
]F��>L�b��fF�n��kɘ���'z$,��ՓϿ�A��2�ki��v�a��<�gܤ�U�胏��S�%��'��3���ʢwo������|
H�˶�W�{���_:�jҮ˘㗞OJ�ƙ2K����1�#K��%��u>l��b��.ּ�W�?��:���s ����2(���5��U�M��{�3�H���+�!~��l�ɫmz�|2��5��V���& �E#`Sfr)�A)Y��avp(@�c�������L	�5�e�1yN�A�HG(� W@�M��l�^Q09�2���7Ӎd03�(2s��g`���m��0�T�շ[Ep�Pt����.U�pʡj!��k䁙�L�3��#M�B�$�cn�#�J2]ܔ����d��,'l���S8N�wm(ug��3��Ͳ��4:�
	EW��|F���]p%Ĭ��*s��+&�^YxI�7_5���~-��yuC��ƨ�Vv<�(�6����o�6׃���:3�&��+W�|-�1 �E��W��w�~��U�`kte�{g�m��V���foNPJ���Y�/䙉T�6(P�)bU^�Ӹ3 �x�����}x�5���������d`d	ww���oڰޅ�b(L�������MA����c���͎�6�*C���Ǳ@^�$^��3��,	�$��*l���8�Y��)Z9r��I�E��*�����}.�"����ٚ�޲�����%��J��xOP��} ���\�~�(
�rF)>�-?h��0�BPX�9���\;�|�W��9?(-��q<(��,�E��ٺ��I_�l.%��ޣ�����O~�p'�h] ?�1 �O���+�h=*�ÙseL޲$Tя����T��b��f��҃<tU�t�DT
�(�c�|
��G���-�A��G_���2�Tz8]˴�~��
/t��sE��<ت�	��Kd!�`f�%al��⩛_4<�Eu}��RI���Q��[��#�2�`<Sa�4W���?��r�9��Q�?��~U�M?�Yp1�)��G�ּ�5�=e]���@�Ҡ�� X"���z=IHK?;pR������9,�vd�A��t��ء�	�<����&�88�����/�-f4�*�1�䆟k^2Jơz�!���JI��K3��� ���.o F��;�N�a��Oa�BX����e��)�ЍR.� ";��!:���_���j��� �F�B{tYO]W�:Z��zr	�Y[m�D��E]m�y0�v'��e��I��_j:�^�P�֮﮼��T�24�^�̎Ԁ�����`�j�!�{��ʼ�U�B�>�֮��]�i��&y$�� ��_��Qd%�6)af-j�j��g{��@>dYZ��	N����T�F ��!G��j�r�H���2^q�YO���u�3lĊb�����m�'�+(���#KҬʪ���mdFhS������s�C!�`��mwh�L%����:����@�ƃ��t�t����֊q,�nm7|��$���>�����i۳��2����P�0_�SeƏ����:)��1�*�d~٬��~�֙QS������R�b����B�ǽ��D�I��P����*�T�0v 5���F�Mq��1�G��j[k!/R'����#x�h�#��ͧ>��$zl4F���d0�b��鸓��4I"���V.ؚ���R|�H����p�M�	�iAL�i�����ڶ�q27�_2F�1 ��j�e��ZN��nsNn�>���NmLܴjl�V$����Ҋ��e��'u1�PW��kcO�7_�d/�b�m+�U�ËV)-f�P���r(Z1��e ����S�zG����s�8�C�񃖺��@��� �x���U$��$<2˘`LA���T���CW��)K���^��N�����D>���5�s�;~{�wPb�4�*��d���b�I�9y��bmR��4)"x�[b�qp�9 �:*D�&��Q��m��&\ن��!���ZR:�˲4�ԑ��0�U(; �9jT�e�:��c7�`o�,�����YnCn+�Q��־��t`�;��Ԝ	�&OWն;��h0{��Z= �S�
6&��>�	�b��+X�r|l�R��ɋ��8NԜ�I�R�?Et�c�yx;�����Y���n T}�I�y$gjp%��B����WL�bD|����N�}����Qü�o�oV/�;����|�m�
9�M	{!��n���ڢ ����|+s������	��EL%,�:eB�;���� ��� ��<h$!��l��#���y�2ֈ�e4G/����s�N��#M\�֛;�(�W����^m��]�>�7���f-�K�,%��!#�lʻ�`��4v����������kBR��=j�,���2���m�s�h��B��ß[M�u*}���R���B���)���ьa˷K����~��馌�.{����R\}��(b���9n��y!�2�����Ͷ �ܔtҔpdٔ��e�>t�[�*bX������W�O�_�rE�=��3Ξɕ��#j C�B6ս��m�Qc���m	���H��g��)fIb>�B��J62�@�9�uh�Q+��4si��c�=�
�l\�Y2�'�i�@��)�L�Rmn��@�^�`>���u㾀q�ֲ"��_��7����i�S�ቂ��¶���q�ЮL���Exs�X�W�&�vS�[Ä��K,ѡ��EE�-~gq*�e�H@�#=��FE��o�}�̷%��*㿉7g�C�Z�<��&eC�(�BO��.��ZHlcY�/��H���icNIU@�!������U�P�i��%2�<���P��l(���=�Lun�i`?mh�S>֢4���!޾�kn�4�Yz|)3���N�0<��d��� ;ZIH�I�"맏Ќ���`Q��L�[4�*�sl<(�v���_
�Ǝ��8����/$A��oƐ�q�&�	0��Ax�$�j��T�zf.hib����!�(�� m�Ϙ�1EA�R��_��PL����cӡ�Z*W�O�����4���)�ʛ]�c��'.e�6οϿ���+��ɷߝ�z��r��i�q��;5.��TE|z|�9/l�S C���ϵ"�Q�3��W�NE�z-���e��8RUǎ
��.�VAhNC�HI�NFd�*� �g�x�d�ч�ςZW��%�B����E�j±�3W�(���zm��>x#�n�_g�N��1N�j{t��~�&V�64c춀�+��`�3�7�S.�Wz?\�t
�kUv�5�s������������23�E���噢�X�ad	��)�%��j���N�]�ٴ�u���Q�o�7�wɐ�ͅ{��98O����;�a7� a��d��i`n�Ð���]&�8:��^v=�$�E�eM�7�Q�Gٷ��4����`��m_���܆G�c�L��{�r�����Ĵ˾�
����x>_A�>9��`i�x���!�z�y�a&�;M#���+���� ����S�S^6��}|���1��΢,�o�����(�1�LZ�l�ƺO�fT����U���qq}x��&aBϱ�/�3� �.�X���U�6&�p�P�9��ZT��8@��c�a���YH���@�I�!�y�ڵԺ���ʆu�~��2�*� ��H�]ՕFӯ�V�V-0�(azL+����%��q!A>����2F��5<���&���m��q6���3o��^�8�C����;x6�>(H(@L7�����ʖ���_#�m��̨q�C����11�컑y����A�S��c̈�佇�g��%k*����e�����%;�:0u~���l��h��v�26����^��ƅ���c$�.��Xv8�4 ��7F^?��3���Gg��������E�򭯸Ga@�  �当SU����-δ���m>�/2&����I~��� ��T �k�uD����[�+��!\�R~O��6�/M��������Nf�L���9"�������*�9~#��(ʩf�UA�{�9�I��i �S��z�9� ~��%WP���fas�I�Ѳ0nQia�Z7YM��K�'m�Þ��
�֕l`��O��z:�/���B	��AG���՟6�l�ڍ�r��r�@�^�&s�2=��0�d��mp�&v9����`ږB����c�S�W��PfM3N#�� xiN,=H�2�5��`��;�K��ZV��qulF��_d�)-�Zc4}	q�I<%}�n�-`���Xi0p����.4h�4�usG�3Ʒ� ��x9���a}g�(�Ir5�m71�Ү�0��W2��߮Xػ]�Ge%,�
�rfO��ԘtM"����Z�F��M�6�K���{]=�lH7��Hjx�q�nq���O��[a�t6&��B���tT��e���ߛ���}���9��-_�� �n Ͽ�pz5ןP�P�@�+���R�C{�._�����n�3�u|o+��9�ˮ�IVǎ�2��&�}t�i���ػ��<J�����N�h�T�{�����M��F,5�G!� !��6Jю<��m��ݳm~Će�F�c�0vtFD�i�J�ԗ����.�ib�fN�#_j�eƞ�]z�hί!\L����7]P=+�R�9Q#�Q#�0Fw`n5�����H�����l���ծ���/u�=>��D'*B2M4��n��H�D����,tG�9�g�l/c��\����4�Rc?F64��I�::z}�+�p�r�@pD�Gge��`�I��:��bT/�]Ǜ�0�$xDO�r#�ek����Eb����TTp:��"Qp���`e�FI��Z��fո]W��(���;��Nr�늤;�1bN���s�=(l�PgL�d�";�
z46�)����q]'�~k�/@�d� 0�e������a(����[f����l�5��1/g��Ƒb�*^E˖$�֋��m���m�Ǌ�H�5߱�S�����4@���9��k� RQ�&Pwl����d�`�/9�ޮp��?F�A���"�Q�P�ׁcy�+�L9L�m3'X��<��/7n���]ӱ3�_���,l
屘;I�������፷ld��#k1��
��0��PѴcaQ�En��Em��V�#թ}���*�UZ�dX�"]�]�쾽�r+5�����Tt��I�Y����X�A�-�/��	�M˕!.�c���v#�����1�4p�F��K*U���)���rƒX�Y1�&��I�ݒ��x!���Et�{��%n�4��9����C0�I�G�f#Q��E͇@G�2�/ZIg�/���1�K⥴�6� ��_�+��A'%n���,{�~V�mm��G:{� �v �x�d�-	3��c��mt8�=o��Nۘ&b�X����6�����-�{��<j��.%�~>M��v�9-�LDE�!Ę���]F����C�!vMX�%�N�&�K����$��T� �\�H��taag������)��F=*�6"�<������lr
�}:?;ʛ4Rnc�X�ƱP�0��y3�%k~{�O�O��$n�7�Z���X�aQ�)6h�i��s����ۦɘ��!����s��|$��y���Y§���r���x�A-��P�Kx#���co v�&k���L��+`I�(n!Ӹ���͠��W�Α|�f�Nb =\�L������_n������7�Tu���:���ZW�A
�sh�� ED�!�w�iW��`)��r\U�3��7 *���L\.M��h�n¶��y�Aݱ��i��A�Jvg�GH>�M��S���K�E��ڐ����&�;�X��~��v�Q7�#0����p�e�@���0L��9�#�rW�̧���n�k���-�%�����l�!N��H�ڟ�̔���l� ��_�,�e�?x&���%�p���v��H��������]_+��u���cxP�����  v�O}���^6���\�g�8���M�1�AQ�L="VS0΅͎�t�HG��pz=�r����o��CqE�a���۸�?����qwrj�6��]�5��'�!ᤇ�-C<�*WGO�|��E���A�qOXp�H����=O��&�[��*��X�� KL��ϒ��4���u�VAq8q�� A�� 	��A�Cp��6�	N�wwww0@p���/[�Wu�w��y����JU��zR_���n-���a9��7:j��,K�:f@U�X��]{��{��ܭQ���
����y�(䮖ޱ�-i��O�7]���塰1��[J��\\�`l��O�i�P��A.����ܒ����AM炞���*C��p���D�l�Jj�w�~�D��̙x�
�9��f9N�Iψ�	��#�,�-�nk:�!_�%s�6�J��%JZ�g[Yy�O���������]���7�>;�@~��͍^�-�!*�d�N�f�LȱӦ1��k����ŮTR���������+���B�s�5�+�d�8nڹ�����@�����?��p��Yu��vx�.���vձع)�s�]ce�B6�QX�G��WVyB"�E��b8s���\�蜇|3̎�7����䞌���%kt�O2@�>|���҃�`�����Z�;N�1^��+��v8����m�X�+e�"ׁ��B����W��c:��s��~�7�'=QӼ3NU��C�X>�!}����m�O��`�M�B%������N;��Q�cOw�M ��ׯ�$�E1����P햞M�j���5����8]�Uy�CX���|�9�� 2�����F}����m3��7}�E
�
~
�.�} G0ʇ,��D�C�?kE*��A��U<��PZ��w��XCR�[_�oW�+�<D������fv����z���6�����H^�ё��U�i�!�e��;��f�g��q�޷�K��~>|�a���DT�K�s���݆L2�+���~��47����͔Ckx�Ge%����l�>�6��2���g3�_��L�ς�o!
��{���8�/�њ�0��c�ݎ�`��c/���%�柙�8�J��Zp�or�Q��x̹	=�bd��cm�g��!��	�C�7iR�W2��l�M=O��6
�?�*����J�Z��#�L�������>��#�����O
�6�C��F�Հ�s8rm"��
wsj�fڴ�)���oOZ��S��j�6����[7�ܨ�]&�7!T��7N�I�b�qw9������c?!َ�y�E�K�$뫻�D�g�������b�����f�Nm_�r�0����i�~�h-������ʏ����u�疛2۶S��rX�2��m95�j�K�
cK����=��h�eʛ�)���ˢ��wp:9���d����en�� 3m���Ճ��랯 LV��L�ިr�q'�Ƈ�R�$���/Cڔ��-����߼����(����/�y�zԇֺ��ۏ�ˣ�J?��@�H���3q�v�Bc��)��Oʹ�=-7=�ǫޱ��$�V�KT'%_ʞ#��T��,�%�z$S�Z����y8��}���]U͑1F#�<G�w���[�!Kx���^l�Q\���L���W@c] �!������@�#`bF��!��YeF�-���<��:��`�mm�n�3���]4[��Ǵ�� �	-T�� E��,ߣ4�AC3%4����s����w���-�}�!�!4�os�,i�4�W�'���<m}��S�-��ʦ�5{b���v��_N��4�#�FGͅ�w��p`L�M�e�[�a�ڽ�4���;��*���[{��z�ж���k	���j5l'}U�5,��|@��������`[���P��1��n���UZ�8��7$*/���[��y_�bC��0L`n�N;�|8.gb�X+;�n����s�Fwi�8�����`����5VE�I�?@ܹDk�вh�ޤ+�`O?w^���n=B�b���w>�`4�5�����V
#��p��1`�qͻ�и�o3�i�,:dݥo{���\�4_���k�:�+�o�\0��	{�	0���K[��~�v4���������1�����6.ܣܻ��G9�iG�_�m���+�T������܅A_'&���m���m���T^k9���t�j���єC��9c���Ƹ���B��cp��"!�`��}�H$���}D��˫��%��G{������b�b'�J�
�چ�C�])�O+��n�� ��u���`�X��Q�1�VdnNR��AC�/mm�W=ܞ,�4���)5ĉF�I��i/���
0 �4��6��Hs���ώ��fN���s.,��<N��md�i�ƹ��(��k�mȟo5�I�M2M*U��ll����"*�D�]0#����IXNU)���q�>����?��t�%���-�IR��)�퐑=�O̶f�J���HJ������$X?;/6�r��
(�웾ڲ�i:m�Q*0�c�({��(�{���շk�0`��B{m��`(_��M��c�Ob�x�Z�
4�GB���w�e/�ԟ^�fW�ڈF�v�D81]��[�p�}t���jt���6E5oR�K�>�Έ�4�}�(ыP��8�Uԡ g���%�� (5mc���l]>��l�Pf?�U�R(���K�CB��nNF��d�K�h�D����J��gꦟ��U����0g�i�Ge�A$���̰�A�Z�c����z�+^#�I����g�eaE�^T�z|9	tS�����u�S|��s��-�z'�WkD���2�n
t^w�/�׿ES��W�=�,�-�+�v}�U�N.o2�`tSPm���8�[�fM4|� k��׫�e�B���\Kn�0�X����w�SYQQY/���=1}:����(�|͘i?�f�|Xgx(��<�&Bv�f�䙴k�h��s2�̵c����y$y���'įΓ�TP�"�Y��v���q��k0R�Gjv�9�"B�"'W�K��)�и�L�W�����^"�����D��T�,�4Am5�;k��'}2|#��K�s��R����9�&b��}�4>!��n�L⹵sq�}�Ye9�.��O��C}n�7�@M��U�>m+Q��2wY��4aS&�!�:n
v�>'�N�M�vch��S�I��S3��u^�E�U?N&(pzN*	�;��3W:�_y4��Oݕ�8þԡ^���|�����
�b3���o��4D\���g��N���O�~2H�ܑr��D��a�����v�|�@,k1kAM9��h=�Ƨ���z���6�ފ^��̹f��$E}ֺ�mf��Ƞ��.}M�,�u��.�+����Ǜ����q�G���'��8�L�� ��%�'��fv��d�+��!�:���,�L,鿩�����^�<?7�����Z�R� +�����d���{�ϖ
u)��ю�4M>��~O��UJ0��$Zɵ�P7��wWv&�� �[��1�}E�;s}�xL^l#�3�+��Bl�o�b�P�Țh�K)Zo}�g�T�������%w�k^��:�<*���؀'������:)s� u��H\A�-%����dC��3�J�86�KDb9tT�.s�`�/,։�h��w����4	�]k�y��.����֚���o+�؜��\��k��n���V���Ӭ_+#���W��,'ߑ`.��^����U(�챂D�1�qy���K�e�D��#��B�,'I��W}(�,�,f�<=�/�0����|��;M��$����]��([4fڈ��ӟ��o�gG�ʦ��k
��7��5�,Z��&�(��3��Jh��Ժ�JP���MR���H88{��K�-]@���;`����o#�w� Z����X��p�	�ל�t[8l�>����9��a����d�{{���c���G��	[h{�Y��'6 .�jPL�p�����~N~!�/H" ҵ�5�m���l��P�̅����#��B�l�t����a����7���܇-2(F�;%{:%eKy�h�z$(�g?�t6O|4Ώ)ʖk�IF[OD�F�y�a�.�*�+�3�*w��Zw�[8_/I�DGF�d#A�eD`Z���Va����;Eǝ���V)���\�+m%+���8�U(.qx� �K�d�EOI������R`!�բ��Tq<H�0L-ԗ�d�c�<��+@ƒ19����9�V�>��z�ܧ���"�l��Ah"���(.f!�H��� ����%�=������*CJN��gv�Z:F7~v%d�����}��~~m�1�Ʊ�)�R�S"A���4)�O�/�q4��g�w�cӲ�U�bŊ��Ⱥu|����4E�b���R$AdKÓ��]�-j+����;���u���4,H�X~A�3]��)���ۯ|��X�y+ �^jք��L<�#�i��M���$1RX_&�_�����P,-����Q���|��w�F��'�+�K+�#D�Yk9i��d�,�'囂����'�9���ߕ����^L��/���.h�g�W�0��+��0�llNT-4����}��1��X�4L̽�/Fe��?]���jz�L~C�Dӏ����L��e��<9���f�:���/�W�I��`%�j�9C��3��.u]~x��/B}P�9h�#�K)R�<ɬ6����g��N�W^��W�U��5ҩ��a ���,���Lf'XI��]�"*�÷����o���������51��;g7��9L���@����0� d�@�������8������䲮��;�
8��N�!ڢ��M��#�rM�_g>-i�a��Q���M��W�q.���D{���E�5w|{�����#ѷ�S��ƕќ�2���F{�K�-{�4���R��� ��M�+�	������ۅL`HJwd���W�&Ns�0��֊̨��6>2�����}X}F�x���`�5�s�Ǝ�"s����߱��CЪI�̌Ɛ'��a��'~}C؎"o[ډ5�bd�=�c$Z��]�˂x9.�~Op�flt�>g�b��n"���K�>1>��!Y�N��^���T�B/��ߑu\b��0V
'��\�J.g����u'�#"���/�h3*�D�֮'HݶnagɷO��v��~��K���J�\q�:V�5Do7ޟGRU����&�t�x�y�)]�7C��[���b��;��Pu�U�>�cy=�X48��n�Nߜ�s���.����_�'?�F�	'���t�Q�_V����A���:�?�*dOmV�n�T$ f�K�$it!����T�(v>pg�h3��wg��� �w��h��1Ⱥ+�i���CĈ�1r�@�Z���lp�B�ͮ�C/�Q&���;9D���%��?%����O��ߕhb��@��eiA�AN���)��B���5���gu��%�������%%�!@#I��J�t_�(���~u�� F�jb��:M�l������G)�%�TEZ����,��\�hts�ڎ�
�z	]�d"�^��rB�u�q��w[�1�*��.y��n ��:.^!���g��b�L#Y��֓����ã��5�$*��_У��������zx���\���>O=��!d0[pkdХLG��_��}�2��$�q�c��;��z �����ᨵ�㦮#<w�L���`��曩%������FsZйrq��T[m��8�m5�2aa0N������8�/�a���)��m�CY�U�\~�׶�ӑVv�������D_���s��ƪ�72�o���P&	��7_��]��*����n��f���E<��,k'���v�{����Q�CJ�D�.-w��
�ۖ�nm�w*����X&_����\�%"zjF-�`O�@�݈�!��k�s�]��gLu�Y�,��6Rlo�l3���%�����䍝и@Ffq��āSύq�>a����P5��<#l�Y��Ç��:�ɿ��o8�� B��lxp+�T�M]>Az�Q2mG�3仹���U%���4���X�[ڂ0�c�����Sp��G�����_��
�z�zn0�K�2`����B7@�;d�du�0d�� ��xqò��Tܒ5&JXa.K�mH�'G���齐�����~o��)��E;~h�ę/~gM������P_�
[?a+�|Q��������ިE[�c��m��N��S�d�
 ��C���%+�)Y
e�v�m�ɑ�w�T 8f���_�Z�bϳ��,ߺ_���Һ��U�҆;
�eFL�6M��?_&w{�A�CR����� ʉ3":��x
��L��2i�6Y:�����m��ޠ w����n�pIq�^��\�n>��׷�m-�c�llTln}4�����4�K� �p�Fu��)f�Dh��)�\�KI�8@��a�QR�e(b{;��ߒ7����$|*��jXBN��&F����I��2�z!�ϟ����J>���l>U��k��gAX��D�����I��-lR[ʾc���IX���7�L�^��7�/�U�5��.0�nS���[rMI�Q���Y�1��������ii�}��3e����u��
�2�,�di|&�n�8���FzO����Ȧ6��j�).�Ϊ�A�(W���}���|����xF��h�.�u�%��b)����C6��!�u�����U�����(�Vow	^�i�G�&E��z���{A`��W0���s��V�9�Ȅ�۾U7~�O>E9����ȌR,� ����΀eB�ɑQ%�%���m��yp���\�c�:�K:��
�Rp�I��L�"<*=Ҿ�F��mM��w&�����;glc��)�/�m��r�z0֭W�-9���Ӗ�)]�bb��-�NaUn}�J`�A��+}���bL�ߡ�I�ˍ/阓��q��7Ըσ�����1e5�3��9gkh�>G�
o5��Q��ω!�I��g��)��������ri�6��n���Q}�|��	��-�Ng���|�a�t��4�ȝ��������K���¯�Ԑ���w��;s�nZ�OU-Ћ��Ѳu�����RZ���\��<�h�=�@�t׀��-���,c����A���"Zp�w�Rf���8PoW"#�,9ޡZ�`���tO�72<��6&Jc������o��E|��5�����KA��@Z�ł�g���qK�e��Il�ݞ�u�cN,�~*lE����0̵�'�����U^���?�G �l���k�gj�Z{�GV��3�A+2�=7�,ߩh#��7|W�zÀ��JH�x�m�,��w�i�o��~7%�sK,t#�L{�MEg!|C5	�`%<�|rI�5����i��E�6,�_;3f��'�	����b%]�७������sz&+�S� �g`8��]z:#��uNE{*���"Da�k����c��򧛑� �(8�Q���i�F�UU@�7�u#�����,�Q;u�B�E ���7Dp�����=��t�p����O��6H��1�c���.�^�����!>����	{�ח3�����OIY<RbG���<�R\P��&���A|ŭI�����_�&]ޒ���j�W�r-�wѧǑ=��0ơ��0��U��+���z��k���/�\��U�)eļ����e�
uP(��7�-�!!�Ve�<���˨xm��P�C}�����ʝ�@���)3|.�iP�v"�NGPR�H���7��d�'k��
ٱ�u`��`������L��ƌ�;N��r��<�{>����>�
J�H�O�kq��i�9���A�J)�AFm��1 I�/1n�]��i�~�9�qr�1X��>9���6!��ȝ/��Rʗd,�m���P��$��w�[�O�~B��x r^J��B��\2q�ZX�B��;1l��O�G���i��)��P�T,����'i����~�}s2�p��%���heHC>od#H�|�&�Rp���Ȧ�~U�L*`z,�Qn��)FyΞ�q����9�3��ԁ��Gub�$�p�cQ���s9�q���,yϢޤV�2��d�mP5^�p�Y���L�
] �����Ɖ(z�_!!�&��^(>�V/1���\������MELwE��l����G(�JA��z����\������/��7	������6��$���?d�b���r^H@����;��Uz��L��P?�G�'B�6�??y�����0�y�-�Ꮵ|�tL+4�k]ƍ�?S��޹��� k��c�I��K%Y9[�/�%P��n���ſ�<�}�76�җ>�NPd�T�/�sld���T�ẴvFV���)y���a8�\�ϿP%�,:l��]���	3���[����!��ce�_)pxs�Vc�e^��K�w��p�U������®��?ʹv�`.b����MX���;�� \L�ێ,i��_忓�s{�j���_�Ô|NM�!D4J�+����z�7{3-៩z�l����y��H�jH�1x)Ͳ����̆�xa���N�ef[�P_��go�!#ղ� �Ok2S�(��<�D��0��H����휭]G��II��)����U[��?�:9�ڗ���������ۊ�G:�E�de>�B���Aչ
BS	4�Ұ��-/']�_��[*���K���_:���q-�t���Gz�ņI��jl-��	����[�wx�bO??��1�q����Az�S��o�q��p����b�5��-I�n����D��W�;�y"�y<֮~1��f2[pޔ����x@��	���w�m�'�!�[Z�b/���b���n'4r$���h���e�WG敜����y1g��#����h6�EL$p�Q�bڄ��@N�蟛�e˷! �M��ܵ��ܵF~�(��]@ �oD�G��=�M��&Wa n\�k�d�/���\��L��DK�z�E`�2����r��	t�M�%Xr�킞���UGp4l(v>	K/����*�it��v�z��fu��;4�SV&7��6�<E�P��w���%�%:�ܧՍ\��@��-ڰ��zPT�g����cr�g�`����=�=�	~��E`������P���8S�&�k��>MA\D�6�>��4'9j�,Թ:gJI�*"I�����d�������-8� ��ѓ�1�Py������e�@�D��q��jL���Gq��J��>�u����Z9O�{�i�p��b��_� �8z?��x���0��P�j��2���Dڧ�j�s��� �5{r^+}��jM9���3E&��%��7z~XL;���.���z�^΃�}&���ey�?ئ�1�T0s��q�K�L�?0�]Y�a���?��������/�}���Pr�A"9+}�jC�oꛝgp���� ��`��n��	�Լ2�:����}�;+��s��������@N���m8�|b�w��O�b������ӗ��-��G�� d,(H��>��۠�s�����F���3ts2� �0�ܠ���-�U�O���XO�s~9$E�����Bw(��X�h)}_x����녓�&g��26s¸�T�n��4/<:fb8#����4V��l) E��%P ���"����O�5�%����o|�G��:�a��!;���%c?�����结G|H�F��W~���ey.}B��b�X��Y�@�b(�s��¶Z�%�M�٩W���4����P��Ri_tgl�����I��[��\������d0��MZi1R+������fi����<Y<�=i!R4|D��m�'��� �T�3\�٨('G�ܤLc��-�?DLϑ{ϣ�<��^Vf|� �bQ"¹G�ũ�s��f[aq}X�Ŏ��,��R 6�%�K�V�ఠ ͻ�LL���B�w��mQ�����B�j?ȼK(xN��b�k5d��'>I4���d�Wq�W��wV�Y��3�:�KD�0H��*Paw i�C��Q8&���>,sX'+�%P�~2��JZ�F��=0F�Kʁ�Σr����s�U�]�+rTqӼ^�M�TԲ�I��T��5=21O�o���Č�{�M<���DS�hq�Ƒ�������<J�����?�M���9òeۉ!w���N^sW8q|�ɂ�;�"w!�5��\��eW��e�Q6��S���Q�Ta̘�H�L}������6$���qǻ+���X�*3�Ckyܙ(h�����1���B��r���/��Z �!����c�ּ>�n�u�<�v��<O�c����I}�i>�;��l>�d�!���dF)��O2�k�^��֞кH[��7J�~�!䷷G\�ċ�N:�^���S���fMÞc���o�Y]�T�m��Z����TÑ�Є���զv�Σ�c�Er�N��뷘���fr�TS��D�+�7/G��Ѩ�]ؘ����j4��~�t��V���Qv]�Z$O4ngR���)�ŕ���Bf���.���T/���+`&
dT� �����v�p2���L�����k���]��#��Om���[�t��-����B6⥹b����$Q$]�����8Ke5�V����yޡ����Bu����+�@��ґ�6��hd��+��.�NNyw!h�<�;]�e��V.�k?�ծvp9s�?
z'f�R
�>A�drM���0��$���Y�Ѩ�D⏦h�KԢ�/8�Ʋ�@�b��;yq&�u��ҡ���+ ۪>�$	��w��,o5��<z�Ձ�^VB�}I�=��Čy�s�@3��괐�ːZ~�,_cd%��i����,e�=xt��N�K����T5�sԻ�-�]4��JHB ?�E��r���rPM���[��n���{SaӤ�)T�o���rl��t,����l��$$3��=�q�j�������jO,�������Um&���ޝ5���V�{	t`ХJ�y	$�0a@�>�������H��(�]+6Nq�,W�'���q���Rا� ^�{P5J(]݅���V��� ]���jw�}��$�d�.���]��F/F�&-B7V*d.�iP�k~��|���r�:Rۧ>~�����ԍ֫��C�=��/՞��	,o�&�]����1���� t-<t��"�#��D�b�a�������oY�[S����/o�7��MD[V�^,ّ8/m5����E����ܥm��ۖɹ�A�B�oN^K��O��P\�z�c=��Af�Tk�~R�5�"Av���;U�O%�\M�`?�	��R�Z��"�L������u�b�n[�f�w�����fG�M��(?x&�9S����p��V��KH��kN.�Q���k��qQY�����ψP4��$q�ġ�l��h���z:X��2�8d̂`�L�O.�wkcIZ>����Wm��I�(t�^�M]q���t�Qc~x���լc���w��d�'͐�5W�%��7N>k����l�����q#ǌ��^Mn����=��HYIR�(/��$����g�Kv-�����(����Z�uAЮ����t�`rZ��z��APr��;�|����%�� �<G��=��Ì���G%tM��?n���Ao�b;�c�)�-��������/�m���s��;�2��P(�{�
0��F�� \�2fF`KV��n0w%��� Z���(��@��xI��#9�k0|��+`V�4�VYqN:5̖@?G�XS X�J��=H7	t+nF+���^�(t��x��࿉u
t�t1b.�>5���/0��ي�;�����ej**�a����7a8�x��m��V���h��l<Vĝ�����|��0�ݽB�y(#8@k��;�"\���$ ���h2�B�i�B����|g?������i�ić��ns���������	w��K�g���WU��t�64��S�]y��쟮�
��f�����=]"#��d~�+�e՛���	2�wG/������:�vĀ)�o��33؎*��V����������C�$A��B�<�h��*=|IJ��2�ޫ�w�����v���'��'G��׬6�-���Eh`W�.��Ü?�}�.E�|Ç�����>��B��&��9D&@�0}�Af��B�����|��1��! pg<J�֘�U6%e�+F�v�7���ݹ~	�i��4�AߍK{�c�ȭߩ�B��5�O�]���1a���k�-w a����_���W@`'��Y�~�}���?�u�C�q>ǆ�(��L�J�
,��O9�D�2��>l�D�:?'>}8�\гlP�3辸f��=�h����|����Pe�IM'�o��Tx�l��𡏨R�S�L���ݵn�M;N�M��?�o:�tyX<�� �+�ܝޏ��:Ďe�f��lw�T�6��4J��BA�fW�w���3{�Ȋ�U�J�I�|s�����ߴ$����g̷�ns�x4ӑ������b9�)�^�Z°|���"�|�eb��F^)�Y�d4r=���9�	����p7y�`s>��SͲ:KK��������x��!�
�g�3@w��v+���v��8��*>�s��X)�w�^Ivo�a}�Y��-9��I����+���P���-��OjB��BA}ѻ%���X�+�\��HA����O�B�%Z�Z0n����ǴQ�xoȖ7�d����{j~��BIlYܝy�T��$`B������W�\�ӈ����:�u����M��H��F�u��~\�;�ԑ�;W�4+��U�xO/1�OrPuS3���S�wu������������)W�+1�P�_Gvp�Z�)���n�.n+Cq��S+��՗��4�!:�k:;wwս����'.�6ʌ��(Y��@�0��d�pH�58�����қ`�~�ڋ$ˌ��)������F]���XU9e��y����^܍���]����#Ԡ�QI(Sɰ��(C>��4�ԉ�4*�̬i�.�o�z��V�J^��IU��MG^��E��)����^��Ib���-X����������)�<�ľ��
z�:���
���ndҋ�W!ب��6����s�vGpʩ�l%�:�'0\��c����1�y�m�c3^>Q�g-+k�y����8�!x"��M��yeHW%Ӗ�v�L��o�xQ�a7���R�剬m;�e^,%�o~+�,)��ŭ�㔭��K��(�n��~�`�ʓ��eܤ�v�-��%[�O3�6Ӈ���L��Z�rV� Q�J��έ�q�54�����Hy���{y��CL�{Q���z!e�M�ޟ��Gq��ݣ�,��Q-�w�h^8vQ.��M������p���v;�.RivJ�]��o"2���8�6��f��z?��[s��NexK��X�V?ɒ�t�e��(����,ٽ�o���&�x���M	���p��85M�0��S	�I�Kx��+��;���() 4t�h��&l�������jp}9w�A沸�$g�ڹ95�Qq�N�W ����ʹ�����G�&*S��o��/7���6I�H��M�]o��
�AT��OLJ�6JF�3ұ�IN"�:8c5�����精t��TQ��9���*�Vɧ����E]�� PK   �n�X�jߩ    /   images/d572cae8-d176-4294-a2fa-ef26b385cc14.png�W�;���XQ#�QE��hK#bWK��j�QEkS3�H���֨]�v�M�ثv���Ei�o>����{����<������(��6#=7=  `���0"[�H��g�V�dC�B�� ���oPt?51&/r�h��?w���r���K=�x�mo��Q깗s��
7 �T���f���I��>��׎��-���e-6[ܕ��I���V�)$J�/L��\ѩ�ZZ��	�\J`N�欬�=�=5f�R��峋�Ѥ5Ǎ���uw/3.u��&�_-���Z\�573�I�����aR����/1��W������6�F�����]�8�?�r�v���m�N��
@����{�����K������#A�����7�*�k�gqb`Bp(���#|���џ�m�Y��v��ľ	ăh�f`�
R�
�$�u��g�$2�+I�AU��WJ���3aм���Ф���o�AI�^�NtN�j/C'+�@�3��J�y��)@#�q�[]ٶP��ɽ��'g"����W��!�WVg�/ӿz�a�c;����`��y��
�n|tt.
v3:,s�\GS��,J5�{���Q�Y�(BB!O�; %��i<5SQ�\cLx�+ �E��!V�˶��ߟC�]�^�^�<��&�f� �y�^0���#��gi�C�VM�? Ml�\I���eP4+9�j��!l��?�lAaW9�@�/w��Q���CG����(M1�#�a{��(sl�)���8�%���Qw�̵�zFA熒����
�t�$k
��L3����ف~���TI��9�hB*� H1*�a�O��B����=�)ll�n��P.�6Õ6��g��6�3����x�my�4IQ�y�q/q��v�vwggQĮ��iζ
s��/(��e�~*o��g�����z��v3"އCۢ���.j��"�[�7��3�q+��׵�����Ëvq��ɾ��w�4�E��<��QZZZy��FMCX���lvN#qGD9�U>_�|�e�[J�'ۊ2aWJps5��A�Y!g��q6����*IBz��a�j�0�zt�'}6�N����Dˆ��'qI�|$��?SQb�1i�)��E>+��D]X�Ѽ�lb|<^JM-�(�]�`���_�)zRF�P�_�(��r�7o,������L�h�B�7)33��+�
�K�\�dE5V��ܴȀj�(���<��?���B�����ۏҵh��}�S%-��W�5���?��Zk�NWtw!���t�dl)/N��Ys>������ ^kӉ�#\�J4�������p0�L��?���.ﶞ��p�m3��=�(�j���Q���Da��|�I[p`�ϖQjH��O���I��?y_���)wp�5�����t��R�^���ٴ>b��[���T4&��}/E\�������	5]���bk,��}�)Eʺm�5������_�ȣ��p����9X�<x�[�(���M�Q���*�&DIALSx�FH�5��Vd��3�0W���5���vP��`Y���ik��UNf�k�N����oL��Wa6��5]Q���AL��;88�l�'G� >@�bǾ�Y�4�=�,�O�����{���Gd|<��֚�v��#[��Yc{vt�*iQ�=^�G�A��C�
�������ው�t�#���Įjl\W���:d�=<U걸���R�H��/��c�k���Y�}�/�r�Rn<����"@[���>[����S#+�_��t��ԥfe�$�)�KIZ�e����6Ӭ5�A�OF�;ӦcO��?n�޹<��f�Qk�����X�Ձj�s�G���$����l�Db�Yg��T�0���c�,f�5��'p���n�\I��.,�	���d�����)�%7dW)�[�M��y����X��g�Ed�<He�nA�JB�m���]�N�������٫ZC/�ڱ�-�N�m��t]�J��JS��@S�t�t ����d���̷"C!Y�NԴ�mu0�
���'H7����J�X�R��:�E��+ �MH$;%�]!�����JB�)���a�ϩҘpj��4OΑ��S��)�PK�F��<GH��_�̍B~NA�;�ҭG�����{������+z��T���c���!�?h��z��e�'{Kֱ=m'�U�Z.ՊϿIh�r���>��xb����s�q�PZhi�y�}~����,F�,ۨ0�===,p%с�lE�i��PZn���W,�P�����HF��.*� ��_Cz+:����E��j��Ҷ�C������$�DA�����澵5���*a.x2��)D�/}�UfM$5�������BY��怉���k��n!lBŲ��x�e2y����歭9D��@J�ՑP	9�IX�m�?��7��Y/@���p�'��RX&3胅�/1�4qJG�"ȗ��2�i]�5�0,\^U��CW�Q���ݮ���DDu3'�ׅe���B�<�mP�~5e �@���=�O|u�J�{Wk���-B�uA���8�8F�4��ګH��a�x�%~6�̷�GfC|�-�@\yenO�n�oɜ�9ܴ�ԡ�^�͙��������m�Wr���}�Oqz��+��/p<:����+
*]<�"��CǇ	6iE��r{�TU�����5�)�* M��!��h�:)��S"����2�n�<B�U#�_��Y�����(_D�;�&
�t����0��?EDD����Ɓ_-�N����m�����|�g$�	��ހ��>/bEcI��<��.���՘9~H>�U�:�ۑ����n�u��B��M���ԓ,��r��f�`�9���!El�8�2c#���OT4Wο�xV��k�����l_l�-�Ǝ���yu�����	]7�ZC;Wן�h�pIi�|RRR��k�D��P�g4�&� `"W�=���U����*111��8���W�~�7p�n��[�|	�������^_���i����#Vݍ߻4v9�_����i�ɜ��V��ަ渔'B�E��Z�t�>�h�`��k�����b?Ĉ�+�I�fi{�s;�m���O�Ss��Q�hIQys���:c*%`�#Z����WP�� /$��u�a�`g��0+{]�Pl���CH�ܩ^����L�o������F�t5��}�+:���A��E�~j��H�Q)A�%n��A��,O?,)s&��b<����m�PP�`_��8}V�AD�?��s�CF���	�[����2u�fi0� ��GBA-�ݥ�a�窹�Y��
c�S�����Vj�p�'ڟ�y]XH�k�1��C���\��T���Ь,x�����	���52Zm��9[8�ĥ2�uߘ�w���v��U��5:�GPN_BQ�Bk|Ԙ��D��2L��!:rj�m�Y�X�Ay��sp�&��vM
Z���o�xQy�ݏq��˔�f��
Z|�^/$Tu�ĩ��!�Y%�����N�!��_�ջ}ucǔ�-b۫�h�֓�ժcJQ$a/L"���G�5�88%>	�����1������sj7��o�r(�:޴�B;j�4��R펯Ft�Ƃ�����U��0�8�Ƽ^�+ǔ�O��N�4
���K�F�ZA�ͬ��sd����u��"����p6.$E�<�z����sc���(<~1'��Y��������1���Ag%r}u��[}��]dj2��\�ZRL��/w���u[��HW�����'��$�D���������p��*;O����)�кa����0\��9��Qٺ,���8Wz��a�s��ܹ���uw�%�I�Lw�@�s�[׌��5����
��y��l;6	8�H�в얨-��8^��<��&S_�/�R7��9�R�(s"m�+KW��i⵭2�r�G\�l:SLY"'��+1?�Q@�Qh�������L�_��K#�5c:z���Z�VO�7(k R!�G�lWRh�����iE���l�KN\yM�rK����ʪ_k-�g^ Te��֌�)��^7�q>;���bKh��A�Q<�;n$}z���fdm��niZ��2E~6f������|�J��D��Jg�'������H�� PK   Jm�XrQ$0 ?4 /   images/d821bf6f-d33d-4ee8-8367-12c4d0b7d041.png�ys%L�v�d�gc۶m�ضm{col��ضms�o��_|U�TMM�TW�L���uMG*�K ������ JI�*���i��Q0`�V��j����� 5�xg�&�BrB  ��🆐���Z�  H��u��2��b)Q!U�˿�>����3���[",�ӊ�%<[g���xf���F�����$et���{�	On����O���{�L�/�_23O��A;��D�!�HD�����"	0(���sdbR�r7wL���j�O�����T{�\k~��amkioigme�����'ݶ]���9D&��ҭ��3p9�����`J�u������}��}k�w��P�뫗C����[��o˧��?���f{y�ha��?�
O��fv��7N�~� �fL|�M���o[�7��ߡ�vB�I7�3��N�|�j�s�iOm>�u9��8f/���_@�~��������W��K �𚼭<����\���΅C&Wr��P]�wq���Ҷ��ۻ��#�w��ZۻԱ:���4��xvݹD 6�A�O]�A���m�-߱Q�ޟm;v�;:?��G�?�~��T��m݄�(�a,f�:�C�*�Ms�%]U8�*�~,�����<�v��G&B!�e��ojn�\YO=ND+��}��&�0�)�@a�)۴Q� 5e!J��4f�McՂM�V�d��.�^:g�����o�A�v���B�k�	_;l��%G��b�܀�qia���1�9r�Ƴ��z��yq}��O�M��^�G�#g�����p�b�ޡwCq����E����M�-�ѣ�m���C2F���hm4=���"���y�25eo;,��^��a��\W�K��i j_�c�^8VŦ�|���g��fȆ�@�!ǍO��@y�� �)��pX~i��fm�/���_���-�/�/���#n� ����5ϲ�3#������JNW#����KV�K�A���d�/Rg��?y>�$�������oԎV�`��?_7�n�z��r~m�0��}�w��S�&A2D_�*F.([�hgW�f񯷾h;��Y[�Õ�vĬڊu�m�F�q�{!%W�SF	$������k�}H�Ipz��އ����-_H8���������0|U#� >^��o;����=�B|��h{;R�'߸��?�&#Ѽ����w�Ca�1]�N��q^�	�ǃs�)�@U�VI��]=w*�l��)4�G��#ˑ���<���6����)�.�Y����o�ﬓ�z�Y(���m<�ƛ/ �M(+�7�����}����͞4<�yo���zx���Z�g1�֭�@��@F����4*�Gt�m�>뢸�^�B�Xq�_�l��"�?G̔�C״,�����L������Z|�BCP�+{�Ww�g���F~�Ah�����-ȶrW���x#��[#"}��{s��Ý�O40�`?�C�9 ��V��g;���%�y�/La|����"Ѐ��� ���!���<;���G"�dM�=�]/n�R�<0�:��W~���y��f��9���e}�nff�D`>�^��R���1�8儀µ�Re�g��9�>_�2�����i�8S�Wt�,�^��n�θ�֕M�M\�����7�o�H>*e�jiv���Y��\ �%��J$q?y�3W�/�=m|�B��o�V.:�v�=�֌X3ē��ظ��k���T�s�O��`�&ak�B��r��FlＪ�ʄ�|����Ș�?��1޻s[RK��A@HO�ќ@����K p��5�w+W;�A;�w�H�o�!ͬ�g��ޝ��[�ݐv`��0Sh^��?7��{	5@@�D�� ���5�7����u!kgm4��[~4��W�O ^��
�F�����b��V���]�WR��܂�3�4��k��²(��������vkzj#�y7M �q���7�(iկ�/�`i�n�D�D=�J������9=�N�2�0�f>��u%���Ӌ�����Y)���'���/��xo		���x����!�؆g >e�&Gب�e������\+F[[�/o��W������~W?��<5(&%f��ymey��ݴ;۪o���6�>x/����;ʀ� K��\xuNH.���^�����U����������)����K��f�z$��>]�ɅŠ�^�۩~��k�=�EH�*�˥��iZ��D��4D��7�}��)���9�+�m5}��&���%�#�M[��;~��K;���/���Y�\=d�^j�x�Uǋ�����ː}�u�gdEÛ�5K�y6mL�����L��
�[����@u����Vr�oyw�紦��<�{~�����Aܡhp��Ә^����e���OXvG��ƕ�û���=��-Ex ;����	f!�)����iHXǘy��E@�9	<���z��Q��ȣ�'��n�!\�� qm��ʓmG�{��_���ݗ��8C5'u�l >�{h�����;�)��3���m��uc{~1j���� �%��U�ev��JN�7�QP/�Kfi1��x���N�~����w�bky�D7��׽|G��iƝ�@+�nT~Ͽ����d�T��<��L����b	#���Ձ�qAA$*y8����M�-���ʓ����w/�a8d01��v0n�D�A!]���q��{ �} v�[��o���60^�˽#���ؼ��'94����W�\ٺtdk��Q��p���P��r�)¼g�����hNB5K�i���_RV���QJ�=7i�a�#��	~��P�sii��ժE9�R��&�2p'����Z�5�r��Cf���R�j�ց��W�ꓟƙ��ЖW��4H˨Eo�@��+���{0Z�@�w�w�a`��ocy��V#?�o��啯�`"
���=��.t���t���9?\��wޒ�����q�����O�eF:�׹?�m�B����9U��]	lJn;`�(<�K�*0`�����aD���<��Y��a��Y�G�Շ���'$�>�-�W�ʇv`i�p)��HS�Lg&0[��K$�����ߕ=�u�������v�?s�B�o����]�NP+��>[�7�-�-2���X�B�ۓ&ZԂ������'�+�H���fd��n(p��,�©�#v�r��m�=�|���E3��� �J�����a"ة��f�׾C��5�G!�V�'�5����v%��H�S[Kj����^
��j�xZh����D=����c��'���3u�v7G������("��I��e|��>'6�qΨ0�����#��b��	p�`���;�x�F���p*�16�[TO�M+�N]y�%�9>�8�reI�H�I[�?%�$6��۵�/t�&	�6�mف�)�F��Yc�h�o��_�vn�9(^��v�鱁Z�������k�p�_H6x���/�U]�����pAy�tz�G)�K#�M����6����L���L�1��F����fF�`��O M���<�I$�!��?٨xt���]C�����?�*Ï]��*k�ZeT:v�� mtϊ����~��B��,�ӯ�`����OE9`R���x�_�F��W�Ʈ#�R�D�7�)�<MSn�TUc�zҺ���b�!G�$L#�D�gVzs���,�R�`�5�� �I�������֮mJ��/�*/�Bu�Jt����8؍��)��(�@ZB�[܇a�KqGwΧ��^u[�Jv�Fr|�ҹ
��*�bb.�r�������|b�b�z\�Oǔ�z��qg#�F=��8�)�M#_!1�v��1ʀ!��^Q��!�bNJ�'37ŝ���C�k���������ɟ0fT;-�ֆ��iٮ��s����<�8oG�뷩��Ve���cRXWߩg����ʔGN��i`�młz#b�0g�@��&��%���_�"�*ک�rjϤ�� ��_�!�{mW�Qu�A|b0)<@�!���L����m6ӎ��N<	���������������mԻիMĻ��Z!굔���I%Bz�o�bm�8Zx{[���4jl�AeczZ؎�[48Zz{����'�Tgjm�z`=�<E܉���m�������HEO�F+���}/�kln���5��EWr2���;���~�/�������D[{���Ķuܜw�3\Ŷ�ݾM��i������~��+���;^�������80]��"��x��F���*����	�y�Dd ���v�x_����V���N���ۋq��"������Oo���F�����/�_9������?��R����t[])a�ã��4c̑�(�-������JN�-�����[��F��-n��<	�����L���S=��<ކ����AxO��8'ŋ=�<�*T6S�������,������v�;�zw|+�D>�no]d��t'��u����k����8��{T����|5#'z�&}'6T7{������/tK��Z���&*�C���ɟ��m7j"<M���w�|��c���h{ku)�o���j�Je�.g����2��H�O}��ՎJ�0�Z(z|-｡�
w=�Λ�v�4�v�=ML�vǯ�X�;�M����N��N�ï�B>I߿�t_(	�ߌ4wBv�"�g�z��"&���ѓ��8h�8�t�^�[Mi�z�ʅ���[c�t�v�w3B�?P���{=�XɎ=��+�C�����b��'''��bVj���>�ُ�^�pW�p��z�^-��_WG��N�'�
���9A�A1�GL/�uG���O�_�Ű01�� �D8m��s~���x����呎�g�W��ՎJN�J0M��MLя�U�J�0L1���e���P+������Ν�p�q���
�AФ��c=k����^{a�)��Gi��R��&TaB������e�� ���JKR�P���f�ٙ������H�z�"WP�DY��s������8�"	R��x��A~��H1�JX�'��7T*��c��
��0�,i,.j8���$�%ߢ�j��d��B�Z$Gw�%}�C �R>�����l���b�e(��è�D����a��P �)ӷ�2"*(Q&�"�ɔ�A���S1��hse#%o�2Ek����^��.y�H)��وD_+��d�(�>�{'6.�.�@1*�@�F��f�Fi�����h��ے'[
�+F��QhQT��
#i9�ꚠ9�iҔz܉�C8��T)[��En�biIz47BR"���TW��VYQ:��q�G'�F0C�	NWi��(	�- �Ԩ5㝕*I�8mUs��	O�j_~��IiX[�jZ�1#T���v(h���h��qB�b�
e�!�y��h�5/{�D���|i��;��5��N9y�$�w+�Z�-�<�k��Es��O^��K&8^q%h(�]�1^�♪;mW��K�����8u�$�+<���V�r���P�x�NxD�2QErVu���ULY�	#��5u찋'��J�GF�t���@(ܻ q�r{��T�þ�狒�������/��h�6$���N�s7�ݧ��l�\f�ς�!����1���y�(g9!/������@b����H�v�g��sͼ�A=�ϵ�o��~�ڕ�k��U��$�ň����GV�zm��D��-~���ֹcS�,��s�ּ	�7��74֘5G{�x���͒
1N*�'ߚ�>�O�s	�3��@ӕ >n%
�7n�΁g;��W>�$b�	I��L����P�]�^�e]�9�d&��h�qj[6m��S%ިGY�A�\���HΘN��5Y�Q5f�*�)�X<�6e�8u	�(g��0^�����Z�l"�iT�\���E	�.�����(j+�,��e�����l]��)���L�#l٫��8p1 FO�U���Ocr����`Ie����;��@����(��Ž���Gh�q��U�d�n�*oJ\��6X�:�;��5y�PU�D�U'�)��4Ej!?�&����PV��Ħ(=Q�T�1l�ύD�ړN��f��c�ÕGg���/�nw)�(Ev �a����N�Fit�C��S$�'��D�L�[�P�D�&��p-�-��%T�<�JW�*�NJ�pma�I�J�#�%3)����9A�R�!C�P��[�*�Z,I{`r�צ �ؘUCO�D)RNMP����O+�љ�u�*���e�,e�����*���CS�j  ���Q��l�-d�S���Z�M����%�p���1�~�K��yxAjP�R�����s�����s=�:y��U|����-p=އ5�Nބ�j�FE���@�#5����^C0�#u�@^s�!f���~��Y��q������US����~D�w9mi3�
��x�w���\`�9D%uY\�mn6yz`�T0�|O�J9rz�Yǳ�l���L$\TLt\GC�Ip��D��F�S�����ڈ2>t�O-�+[]���}�6#u�X��棖I]ϗC��PĆ4�iAe,{���NO�!��A|˧�M](� ��2��,�'^�J�ݒ�([���iG�c5߈���]w޽�
�]$f]�`����n���p!���a�6��@�n,s#��J"�/��ZL/�O���2�H�v�#k�ABu/ ���&4_w�:�oDr1V	��vݘ��=�Dj�#8��ȏj֝i���
��Сj��ޤs�1˚toSpr��R*=�Ț����EJ2K�x�VeKw�\%0>�w��f�EnUA�r�%��X�'i@m�����n�H��ڊ�B�U�����C+M����1٩fO-���TfH8X�X���o��~5�R��ڨ�3�=���ڱ��J�\�~�qb�B�jL�������I�du8U5���	���fM5�D�w-���q��5�5[[�0H��I$:N�T��t4�ar]S]I�!e��q�X�����4_�T!|o�b�d�t���H1���{�Ԯ�/0�\^~r��~�}�YO�8ں'R�^I󽨅����~W��u2h�0d@�0{�&��Aʘ+j�PE!�5�qkY��b$y�4�|�h�ZQ+<"����,{O�8G�'�������ܪUK}�� ��
E�na[��Y�-�.P��ðQS�P��d�YVB��H�C�C3~�;Y���PŠ)�[^������<'�2���f�"Y)8h�~ğz���e�
����:��r1��y��{�Z�bR
6&���a�{�h'�s���s�
����ԉwo�
� ��T�p�`�HF**~�료��"�O�t�����*n6�M���y'ߥoh��>�2�ȟ�m^燹��+�S��X�:�f$:6ʁ�	̚�1^.���/��Ͱz���J��2��ɬ*�=<�T�X#��8N<L���4��j�i��'��-.��Rrl)�B���,�*���9t�Y��!8f�����]��+B)˂��ag6�?y��%u�%G��~f/�aS;NO���=C���FB�,����e8�~�����^F��&\�;�@�s� L0R+c̈e�Q��mJ�ta�I���r���0漎f�r���zN�Q�*�q��)��
1����e�6��~��U'\	��K�*�Pl�@T�Ѐ� ���R� �f�f���i|���иBV�+,��2�*�e7��gʬ�����z�
�xcO�I��6(���-*�\��r���CE�B1ǔO��Ě��dz_R�_�R:�m	� Mav�y�t"ab�[}��%ې���QJ*YK>9�A���:�`���*�8:�����rt������$\)1lό���wU�nҪ�YVz�jJ�:^�����������3[������ؒ���E��EPV�����\����௼Li�l�HY4&w!6=d��Ê.QkF��E��S6�9tN�x�9$N�fq�XG�x����5R�-��:t� ���K^Xr�xa��`T�F�r�[�� �y�p
E�Q�h�@��qt�H��u
s��������㡷�V,M�P��J+v-H%�iG�P���mV.T���UBn.P�R�>e�n掔�Ab�N�[[��lD���|�H�Rcz���T�u���d� Q�����m|��`����E�4!���i��y?�������p�5��n������5�ư�`{���L6Bi��*Qt�(�6��>�����E]=%(d����#F�
 ���F%��VK��&M�U>�Ej�pE���/-_��ĔT���螈��|H�Oމ1:1V �Չw7��6��ER���iLN�m��(�Z���~i�ʿ���(ܶLי��QV��1���q�Û��^�Hվyb�^� "��|$*^�F���ށ����g�￨���<~��6��9�Lh���;��FK�����K��\T&R�<����@CJ�LT��ȸ�0;��+x���r�[�I��-$g��b�T�w��Ern�ôz]][�.����)�O�W��b����D���f)���(1�����|8q%T�b�h�:{��Æ��TD���Xr�L$�W�ВE������]ⲍ�l7�n��`����S���7������1/�&�����/�-ˉm#��!���K��&��n�Ƽc*�����[de��9c/��}B&�T���#�1������4u$��%&�$W�F��p�.���������X�!O%g%�'�r���Ϩ�;[��ͅ/ �6Kwd��`r�A�b��.q���~��z1U��L��-���8E�� �7~@h�0~2!�&�I�S���I��F�)1A����e���UH���II��L���߱	�*(�[P�˙V^��@h1����~Wf��d�?7�N���P��Ͻ{��lO�ʲ�1����"8���,�K3�*��Ś���0���SL���mO.�� ,��櫍?I�V���J*g=F�3��KUcX<�<fr1�aB�/�!p;9�]N�JA�]�_iq�}:ROʔ������R1���6^v���b��
�zBL�8
�^��j�B�\۾D�����^mb�y�h�v�����)��N�L��� u�X��LfP�(�n�U��D��5�v���s�40��􃑮������#=_�{�F�Q�퐴�͙����Ld'���̅N����	���7c jMh0�*�����|O�v,�Y���>$Z�ފ˟,�{�N�`��1�9�)_X33ի��!�`p�D��%�y���\;�[U=l�\�����(�Y�}E�1�u�L�Q9ᯋ�>��[q9��_LL�ڑm䮗BЁM�p��"�'#���~8��תG��u )�\==�`���#`y�?m�.2�tA����
ք;U��y���N2D K�'�E!�78�+�0gk��񛿌Ig$Z"���=���Q:mdx3)��� j�y8���
g蒺�E*sD��i*�`���.����_��L��+��s}t��cFsc��y-A��s9�jc8����r4�m��8å�m'"�����/�%�=a���q����q�ۂ����2W>qU�}�)ۓ�h���5o8����e�NW���kk�EI]q�����M��vq_Q��?�\��#Ӱ�eM���v��&j���șaQ��9@��H���|~�x���;���3^iϊۙ:ig���� ��yo�,��L�Bq~ev ���5�tH"K����5�)".QI�ɐv��s�F�Σ��2�*ϥ��lxX�������`A����\�B���LB���zv9ޓX����q���.a���v�M�+��Tv���� W�m���j}�۝���J�!�5��*}6Qg`���&n���lwk�u'���Ԟwm쪧���Dҳn�����R����֧��H�t���)�N��|9)���Z�ۥw$���Wj|���'�
~"
)���jr�r��N���of�<�o��������4�����򥥳�h*]f����k�C�VB���|(�r�^���'d�<�԰j�����ɮ S�ԝ��N3�y
H�zD𝧎'�Vk�n�ñ��+���Ok'��yd��%��!����ZqGo���d�ly�'��v h}z�|��IsSK�m#	ٕܟ����B�PY����y�}�j����ɲR:����e��Tީ�i{y!��7�!k<I�
ho_�W0���n�7�xd��'b�6|E��L:m�aǒ���,+U��G�0����	n�׮	�+��(�O��wy�41CRPX��3�U��ĉV4N��UġF�/[�1�O�p��Q��'�v�GF��J=�@&�Gq�#���J��T�C�_�痛�8��fv2=����j�2Vv	�}t37�c�y��Wd�/�C7"z��81�q�>����	y����A%DyFMK��i"��Jyw�� ���d6�M�Ӟ~�广R6���H9�H-UX��t�U��]�����iy��9��S�+&�K�/����FLz�K��1`$hJƆ���@/��f�-�H���TdI-��ۋ����U��`^v�}{!p��^�4G���Y͵�^�y�u�������,���-�������=�#����FZ��8��\MĽ�%���Q'��E���Đf<�"�>J(a?���'݋�Zb�
��:��1�7;E+�$��Bć���̘+�F�<".¼�k����/�9�T��nl,�G3X^��Tf|�2��_P&tZҴ2��Ԏ���&�R�1����%�dj9�YL�h�5H�p9�>#�,(��y�,)z-���%lOʪu�#+�w�I"�1�������\t��W,�������`4�8�����$������=��g�\�%�'S�aW���x��'��4�5:W�)4���0��d��&e��	����jdJԁ�nu�?�&NfU�E�#�������C,�ִ�Qƅp���n�r`��7>:���g���^���������	�a9��װ˱����<�iSi�X�����{O�&�>�&����a7�-#q���>���8M��׳ȋgGL�����$�[[yP0��ơ�j�z2�ߦ�'����-ُ���[#��"�ȑ�u�:b��$A	^��vy+t*^Ҫ���0ץ��h����Ӡ��5����Bw��Kv�0q��%@���J�pݍ|��X��ڼ��«�vdh7}��Z&H��U.8�n:\.�Dm�=E�d�e���T� z�)X��	*�:�������5{�� �"������:!V*�-G�Iݭ�ޑR[���c�Xq�&W�7�:mY_�=>���s���
Qi�qPc)+�	[�q;�j�V]�d*z�	W��K��)��A0�R�)4B�v�5����)̐����S���J`c}��U���r�M�,��G���5���@��ws�S\wi�}Ʀ�����`䭕MZ�Y�l�y�>���;��o�PD�9�������k�E��G�&j)SKȟ�p��$@b�YR�bhK�8�y�D���䇩kLP��b&� Q"ՅR�0�L���[򹹟��g�����0�@%)�#+�/*�q:�p��Pa0`
�h��	�L2�a�R��:�������Z�	����
�̇�VU�VV��Rk�]��1��؎-G�F���j'qRShX�=�G�(5�ToըSq ۜ #�*D9�6��YJ��ݟ�=K�>�'�|n^H�9܏cΒ�g�ᾲx����X�a��y������2}{��&s�M���.�aNf�z��!e�\#�	�T-Q���z����+�UJ���:k���UU�V�ϻKڝ?V���;}��>��S?�v{�J\`ti�l�B�F��ݯ���7H�����нx��x	R(���r�2����k����D���h85fK��m:���Ķ:�uF�-�F�E|��bfJ���.n	Ů�S�ֿ,茺1N���ar�)[;Bŵ�ŕ�8��^������9�f
��4���]�1W�V8��6�`����,� ����l�`�&jq]�� �|qt�)b6Z�ib�|�#���k��`��!���ŕ�K�"hcD�㫿b���$F9V��"zs)*�QYNm@%
��H�@\FU9=���]~؂����D�s�TQK"���L�n�:�X	��u�&qR��0u`���;]���ox�\/Fwq�{�d�o�8p{-s֯K;J=>���*'�nꌉR���5���ȇW{r�#A�Lu�����KU��f  �7~N�턚5����fx�'I�M�-�K%�O�v��̔j���j,�ǂJ$��NN������g���B\l�Ե���7��ZŴ���ȹ#_f�=��F*Z=��Io�À��Q� ��P�cp�ë6M$A�Q�d��L5�a �ڇ�4�=[$n�޼�e+�i�2��_�l5Z
���4�^1�T�:������|��)㤔� �+�h�J5���Nw�@M[�`X,��ũ	�Xa]�LҤL_�*F�p�0�O$\���Ŋ^�����i���������������U�d3�ѠUm	(�&3�7Aŉ��aaiȨ�e�)�љ��
U';
�;|)�ϫ,iRg6���:Ԣ)b�߷��_���X(�X|�I�"�euB��,�Vh�܆��{>��g�o8�o3TJ&s�̷�<�1t��.ߢի�I��\�'m�cK�a��Uk�%��w�t�鄴��u��Ɋyʰ�R4{jge����kD�Sxpp��4��jzh�0n�C[J�a>C�"������I�lV]N6eoN��J01��P'iJ�ra]��وlf>��į���s�t��{s��]I�x��
!y��E'z���i���ۯ,�dI���e$�KRjb��C�%2H���P��]�e�PC��3H�ɱH�6U��Y��d��]��/D���`���fhI�TY�HM����3RV�0	q�34- ~UE}��jdxH�Vy�Xݼ֢�þ��$i��ͅ���Y
�R��|[���:O����yݥ�o�-I%G��l���������\���_�X�ج���?��k����R��W������-
�ç]�\�V|�V���x*\�Z�tMX(��OU��{�T���L�Z�V>K��<�\?P����Lu6\Ug[��%�<X/BN� �aAa�SoP�Nu��*����z���G_�K~A.UU~�o-4�d�����q9�����@��LN��u$���r8�,�N<���	勩.3�<oo��i�ǥ�v�L�1c4am����9����ρ��'<�d�R�u���M7�z"_{Йsgf���IX5�<�$�Z9�	U;xVqF��6��,	�9$?�$�%�����G|8�jdhH��4�?�}2A)�u0b����Cs&3ʄq=�6�K�
֨al']��>�t%�1���U.�]d�Q��\�{��v�R"��H6W��_N%�Tߎ(M�h!*\����X������4���n,�3ιp��
�'dN����3F0�����h[:v���>�n ۊ��Zs���61�Б�N*Z��k�ڢ��,\OЍMu�����P����v�N����4�F���o�JW�n�#3����C��<�qH�jnO��lKch�H���~l>��dX�~�sH1Nc�E��Y ���ԁ��ǝ�����`�tN��l.g �n��S���1�n��W��Kh��1m�j3�&�J�"N
0}I��ù�B��^]�݆���cL�|�8f�P[G�#FDC�M�[�?����,f��Zt�ĭV�C[;<��8����2WГ�W�ܷz��_M�f�S�c!w5� ]���-7�?a-�_��Z������Q��Ӡ�r�@,�d��Ǯ`°�@q��J�}z����C5UŪ���T�@Y,j�0B3�s�Q���B�����z�C¾���.{�+=6>���rzY�C�WzR�yQr
G���@�ĥ)F̋B}�X�1�Y;���|n��׶�]� �r6�[>�<�L�hE���g,�g��b �[����&���a�`��N�$Y�[Va��b�h�Se��B>�"����͞��J��7$�۽v��u���I����X��s�@�����!�j���GP�b)�e��a�wnJ����v����[AVF0�ޖ�@���f|/ ���CM\(��cl^�㫪�f���2�ʜyꪎ-W�y�Wl���tz�=°5QM�"*���#s������^��_�T����`șd3�8Y����r�"��0��A�� E�n�������MO�>I {yf�Vb�ʨ�	����_"�B���v��@�ˎ'ڬ9��׆��f�ɭm�cv,;��J�P����g4��c���!)�I�Q�&y,�jd�6��~�����;̢`@e*F���5)����sp������"m2����7P��
hO<��Ci^�r(��b@����]4?���kL�35{k���zV�����
����J}�M뮲�cǉE��6�����'����\|�k���l(u �.n�ɤ�Ղ�Q�������J4�S�̮ab���C^x�?�c��6k���$��IL�fS+��I�ҧ:>�T��N�R1K��QQ�z�n<N�|�NC0}^��l�ec�LZ���4�!`����������)"���i����`>
���Έ>��y����u4���9������8���	�Gi�;h�?f���[O�cf�<k4noGj��)Y�Q[( ��*:EOa_=�7�6ZkW�4 �BX"ڍA@�u�;��2�C�lFo�C��`b��u�c�ۖ��D��\����h{�x��P�Έ�N�-N��_�4d7D���̦d��<�^��ZO�%K�:�����Q1h���b��Os���E�7�G�g8L�ϥ�Y\tn4B	D�`h�	�\ax+Vm�HG�<=l����׶��_��i��e��%�� UUբ�b�67��7�4❡T�(�w喚��e8%M���L5�ċ+�"�{V@�r�¹'w3��\�|�i�k�=~��+.�j�]����o�p�z���T�Wm��3������&���,������Y�'�#��A m
�i}YN+�S`�
g��<����tQ��Y���^5ӄ�\Z�2�y���K��J�?Sth�ձ�@��~��j��*��EP�21�>�I�-��~A�����ׇ~�&�W�z�XeN�Rbs*ve�Gթ�ܿ�d8ک/x�_�Gi<Y7 F���j���6��ʴlL_[5�� uW�ӗ.��%:	��'��k+_N[�O���Hi|F�����h�:-�1]O�Ҙ���d���5lhG�a�UI�l �bzb�P�Đr �P�2�5-uu�<�����/^�˰��8
�N,p�x)`�g����c���6��Ѱ�\�1���nB�Q`���WE�7�m¤�5+&"��í`�럹讎R�Kl
����*���+�$�a����n��C��V��;<��w�j�v7�^>J�IjP�hUR��XB���R�Ԃ!�t~͠�Oo,I�_D��ὡ�����x#������9�V��R1�b�M�< -���Y����[�.����"�-��g8:�1�T�HaT	x�{�V:���q���-ɴ�k5Zo�1�����}��}�a�����;��������|8��d��k�֠��Z�g�I���~|���9�}��Ơ���i��|F��DLs5L�@���?<~B@~�����BBA��S�d�[l?%Ka�V�`�k�<�G��(�����4�<�(Fd��������tm�G����=7>�;�(:���%�tu0_&D�Ao�MIq�Ϩ�ݧ[��h�=�����$�ɵ�R�>w�c��m}mHW�nq�Ք������RN\6kp�e!N��8�0��3J��Ň+�ߣ|����^����Z�����(����&�Z=�����𿻎�������8*�(����[u�[�Ǐ~��i8�l�2׸䟒��ƍF&��{�-s�as����D�k&P.�Q)RΒ�mG�bйe0�� rە~�a�+�{��A9�y5MǗ�޲f���*U7L���N���k�0n�f��W��1�H�('EKd6i�n�u] J.���S���ڪ@���۶#�!�D&T.�?R*�^��vG�1.��S�Ш�a�*ӹ��T(������^(���܎�ਡ������)3�E������q�����-[�����Ǌ�$�G�Q�8-�U��C}S ��VE^qB��:��C�p�����|	��XHV����]>�����믄���[��������-�`�X��ƸM�<%���Qa��LҖ���ta-G6X+}1�s^��k�"�""��|U��!�H(^���a@���s�/�0�h���|�Ρg`^������ć�X�OL�t55.��5'
k���9!+"/[�*$ns�C�����O.�TG�z^	��y}��*'��e�4��n�2`�Xk2b'<:�c�*so8�٥w0�݂�L����D&�����-yP�������)M!�]��_�<d3܍�MgcK&k����tY��ݗ����hPGR�˟VM���Er���W����ثO�d"G �����Ј�˦-\�"l���k�O���_��������7_~���Cƍ�4}��ys-��|�╫��Z�r���5�֮ۺaӘ�?���?���O?�r̸Is,^�2l��M󖯙0c��m��<�������lK�ޅA��6�q�t�5���ש������ܽg;��߁,�ojq?/Bn2�m@5R�@�c��h�z���֦��)0Dwv�1�%�RYV�������s�n�� jC�W�[���ΚDFLf�^ՉV^	�A�K��"sW_��|�e��H���L�y�����]��}'���.�G,�Z�V�"	����D~K7re�W0�D<�+�k�[-��_�L���$e��C�o�~��ᵋ��lȯe=Ϭ=�$e���u�Q�j�������.��@���s"T;$�P�h�"T�%�e*tL��^Vh�R���A�2�;��=��E)Ol�8�:�V%��4n-]P/���j�L%РH�?�4�V��ë�vϒ��g_}?wǷ�~7��9G�޿f��Gх\�]i���u���3"�]�3��6�����b��̭W�n93x�#&�ǌ�u��MЭ[4k�ڕPn\�~ۮ��ѯ>���'}��^v;"�"�����������Iawv��7��
"�v"�0��¨�0���*:��/h�8jM)��Q�����ر��ٗ_���{�'L6x����?��/��w����}��`��O��`���+#�Yl���dR�t:����2���O�ibС�t����%4D�La#2�T
ŜH���T�whصћl��Vj-FA����|tP)�W��5�|/�!�*���%�nn�JT B��)Q�1���T��TvO��QpK�*�D-{㵗߹�W��x2�@i�#N��7֕=�
�B��K�	PI�I�׬�k5��~�����>�����uo�p���Z�"'��)����&&�3Z�NEm�Da8�������2J�@!�c��g߈�|~���݋o]=9r��e԰�wY&��	�远�l��3��\�r��u�f͞�������_|3h�ȱ�Μ�`���\�0l钰U�W�[�v����m3bܧ��?���G���7��Z�j�ⰍK�n>a����xF߾��o���V��Y�:���b��ux�������}'Ω��SgN_<��X�}M-v��b��Q���"��<�����\W]S�d��g��0����PUSU������P���ڌom���,G$u�R�H"�����Tx�׋��Z�Z�T.X0>>3��v��=$�A"�[j�\-���n�l�̊U�[����t-�}��Uӌ9��ϓ��m��ܯU�X߱��F%~=���R��_
MP��wNx�`�U�RW]0!��F#-u�$���-4�t�6�{�{���eKWY���̚�:y��U��D^��o�[1�1 .��B�)�i:CH���#Ժ@�b-*QK��%+�ZfB\�Jc�:z3����68b��6��_{Pʕ:�n�Jn�H�N�˫��Tv�&j�~L�Q� �V&�S�ݒ�fʽ�gM��b�W��fP�vX*���K�f1t�P��`���NBHC�7f��
+|�Ԟ��o;�Q�,l���F4}��ɣ��ܸ���}�vl���?�䣁9b�q���f��k���*��jXB5��l���)<�XewB�6�~)�!D��"���r�i9�dZ�RE�T1�$>�A�a����������6~���}��_|�A�o����7}���/?���_?��W#�3�ӡ^�p����7q�l:�MmdQ)L*�I���b�"����G�ɺ�P
"�#4OPVR��);M����K�Z��8.;٨��*gѓش$.5I@����u� �;�ׂ�E"���������ށ���&%�I΁�����t��F	�!�|�J�E�Զ�B�#�Sj� �T�*4��0Lq�0f6�A�2%�A����U�꒤�I:j�n��IX�>)�QA#���VO�j[Y"%�b)�J3(l���(Q<N��w?�ZT���'��u���^U���=`�}�#�[�s��s��-X�|��%P��3��/���{}��7��7~��Y�f�\2kֲ9sW,X�r�U+��	[�~]ئC�~���������g�\�|�U��ذl��!�fl�w��s/�p{��h�ѯ����vj��Q@a 7	�L{N\R��A��QkC{��mN�Q b<���Ǵ�V�-޲u��-�G����t!��G�c��Ɔ*�p��m-���m���s�5bܘQƍ]�`���l�B:���چӂ�5c�_g��f��/_�����>.B���{QO^q�ȌIm ��)�n�*lWI����nI�ٖ���ò]������/�y���i΢#w+��PE(�)��J�������V�p��+P�J䊊���O�����imؼ���R�p��ջ��=�s���3a�֩]ح���W_�yU~3���a����b�����z�=B.B�Vj2r�V�VgPV���s����kͿF�R�Qʒn�򠜇x]^�JnQ���ǫ�����]X��,n�����;�^,�0|X�4P��")�[UM��h�+��R�����P�/�0t���x���:��a��+/���6v����=n�qö�Y�w�:(
?���>�``�~Ç�/��F~7h���OߊP�⊴oE(T8<M���D�Ba\.7-#��B��5V��d���(d���Ɗ��~�Հ�FL�a��>_�y~��_���o>4��C�޷ߨ~ߍ�͸�����wnE�&�rY�\F���X �ˡ�x4?$B�TD~DL�K�
�-2)G�pe>"	��.w�<��D̎k�t�����}���z�)W(MK%�72Q�I���*�֚[����Td��-J-ʓ��JGUj�x�<�(K NH}��]���]��Ky����W;<e�@��N��3ȩA�ʘ�rZe��Nn�Hyj��!�Ȕ\�v!�bZ��^feV)�]õ!�GO.F�[v(�-u·����H��aٖ4��BjZ~�ƪ+1�#R#��ݿv����c,��宽��ck���l�×�o�;}�څ��B��͙��a�?���'��<��s�L[<v��1�fO�<ڌ���X�h����ׄm>t�~��?|�����8lq��E�6�]�n������ؼ�]m�{*>��A�xEh�]�0�z �뮓W��8u��s!��pjtRaZF��Y����-k�m�4r�Б#�t�pXKk��hP������������>�N�<qޜٻvl3j��y�"�=��]"B"|�:3��~ن}5��\�J:aT=yՅ[&�a���I�nǨ\��1�˫x����R���ٙTs�Rv>�q��ۙWkAP��l�/0ap�hh J@�
��Ŏ�I��\Z]^������$�B���h�ҵ��$W5���<z�ؙ����{x�M���ʨ����E{�d���j��;o�2�-K�!�R�S�s�EZ���ZbB�m.��������H�����h�C��������x�n)_�vw����t���ˁc҉]f1��S������\�Rc���3�o㓲q{��t�U�����t��

�8��!�D��0��4�BG�d��+���}���Ua3�B��wθ��&�ذ|��Ӈ��ӏ���G�����СC��=x��~?�r�1]��/��@C"d�5d����z�m�M�����.B�<az=����XCk�f�B"��8E��GN����{�����ða}�M0b���c�}?����CE8j��+���3���Z.������i��(|U B� =t*Q)�!ߵR!K�����.�o��f�ń=���Z��[+]���@��_��W�|^OU��
��Xs���k�b�B�S+P�F�H�3��v��.�夻�$����,KK?�@�j�L ��2ۋ���@;5׻}l����R�a�;��#�J�\(P ,	O��B�!�Z5P�afQ���������r����M	������&��)�;n?|�PU0����9�#�?K{��+��]�2�����������2囯?[{����;f,^6w����]�r��y����FL9aޘ����ȴ�&}7`BX؎���B:�Ï���{_~�ŀ9�ׁE�t.µ;�R�L�"�ʗ�0h^�V5#F#b·v�о��U1�9r���+�z���i$�+�#�oݶ~����Ǐ5zؒ%�s҃WloiƏ��z�j��C{ل$���q�2�_?��>_~��G�Ǎ
[�t����Yi`��u��aTLZFa݊�G*�J������8|�z��[|&�c�(6����?�Q�-�,Å�c؜�1�jx����B���Y�]�t�Na2l6�C�F�+���oE
�/��+�����jen��=��=G?Ky�V6j��G�l^�eÊ��WoOm>���=�0�g{\!���V���h�@�l��k�!��L�P"G�;4��.�ֆh�R�D!��v'�gf���Ԛ�Pv��/�Pft׊4k��-��n��C������Wy}��V��HH�F��a��,<�nǭ�lys�|,�h¡ǣ=�Y�u�<X����z9z+~���C"��p`����.p)j�P�st�M[�i��e�F�3hޔQaKfN�4���������w}��jp�Б��2����L�L�Ȉ��j��C�d��+�{�Z	��ؑwE���F�"��W}���_�f�ġ������?�������������O�懑��}�у?6l��%_���YX�Us�\^=�G���F� ��DT��.��H�T0K��)W��r�L�E��B��@��5�o{R�?x'�c�(�4�3�fI�}�ϕ��B��p1�=��N+��H�I��^�2I�V1ف��*�G�ti�N-�0�)�2U!�ڠ�S�*Mz��Ro��͕fk��Tku�S�1O"5B�/`�E,���@%���%\r�ZT�130�����#���We%/�BKc-��֝� 	,RcIn^�v�֟)��������_n�.����x૱�cj�G��2]-T��]��^���uO��9o�i��O=i��	3�2��oG|3hB�A���:l쒱S֬�t�������>m¤��V��?p��������?x����ޗ�?�3pݮc$��u|�O�5�&��`�+��vQDo�|�*G�<x�ĝ�׃�ڛZp�f�On U<~r��٣P��02�Uĵ��*�^k[������u���lP�����ӦL�t� #�vn�z�BA~h������&O��i�(���Ny���W�jωJ���2RU���&s�Ų�i�;.<;�(}��W��=ؖĂ)�nx�L��$�o��|�ͤ��$/8~��+gjP1���xQ��y��{=B�A T�(���e����������h&����OÓb�>�NNʎ���z����g�݊|��L8x�������S@gx�*��ij�P���68�C���a� ~٦.��P/�v�A�(a�J�X�X����+���c9���ۻ� Ԩ��Ю2{�r��3�˄��S�-.Mk�Ҋ��@o�H8�ʚ�l�F�0*}F=��[��B�� �����_.;����������S�'c��FK�J��Y�C�`�%�Qkߡ�@{\� K;]地�ؼ��'�\0įI�L=h��Q������?����������G�}�]�~8d��a�F�:�ҍ�L>���1��b�DnɌ��+D�-�-mXs+~a��W��K���)B:���i�����O�����~�&�<�����������7�����/��>_�7d�7���ÈF�b舑V�?;"����TsE�A�D(gH Q�d�.�r*92%Ԃ"�$�@���qF���L`h�e��FB!9������PҐTV�T^����2=-��(�ؑ�V�ɬ��:�ReD$1� d�x��¬��¼���a3��I�3��V=j�z�\�)�������&�TĊ�L�B�y�Q�H��e2T&�Kl���d$e<~�t��"Z�,7��b�A��tM{o�R�P��\��?I~RHZ@=�4uř'��8�������I�4"���{���.L���܏�g�\}0p��?~��'���>�f�{�������G����~�{����;Vm=w���'/��6���>�|�a���o��O��~ش�S���p0m��]G��t���:���l�M�q���`�!�m�;6��ԙ���ܹ�;��l��4��UV>yz���=�F�9k��Ξ;^R�g���^0_WB{�B����&�fؐ���y��ְ��7oZw�����\��9�k�Z|�-�V��PPX��Y1s��Ƣ�0���ЄIm^����U�O�[�2����V��"ٺK%�#i�%.�Þ���������TU�> k��&;C�R�l��6�ͥ6�a�����!��b�_�O�*T�?iE̠_lX2e�Ⱦ�;���S�lM�,|��W���}�a��K�]zE���5f����O�Xp���_`�\�<�(�n". X0$B�шZ`E�P�V'W���n
���NZ�Me[q�^����4��r�Z��P57��-(0��&�#T�U��c��)Ȧ���8�-��N���R�8�/�ZmxB��p-���z�D����_Ђ!�pa�t3�g`D�����c֟��������L?u�ș�Ϝ2b԰������������џ���jР��>z̀a#.^���1��F��؄��j:�-���V|gQB�Dz�Á�t��RK��P)�4zh3f��_U�Q���8p�1#F���ϗ�������O����_��������o�Ё��bȘ���7?2���+�Ϭ��)�?��

�h<)N�����cl�
*P���AB9�I5)ʒY����J������6���Au,���S�Z�Za2B��+۽^�#yB�D�"
�\iVj�*�M�w�Q�B��71i�b��abs;Ij+gkj��Z!Z+�5H�t��i�ZU���Tl�A�1,�Z��Jf���j���%�t6�Ic�����5�|~��J�k�E�BQ+��Po�ظ��}�JG\\Ck6M~�qҒCW��
#ǟ%_x�� �*
|^�v�|�ڹ��u�c��(arg��ߏ���Ͽ���a����Ő����>�� C&�ݶa�͓�__y��z�ɯ������φ���~�����o?���~�g�>�߈)ߎ���ĕ��������R�V*j���'}FPt�U�Y�Ƿ�!����h˳��[7���)(H�+HIz��<+�̓G7�l]7c��+B9���δ�DD�ӡ��G�@���[�"ln��Σ8&Dʟ2i����S&�����{�Y)*%"�s�<��+qŵ������^�Iʯ��z;�٢j��l���{HZS���0aU����̉5�c|[9F��`��چ�0L��?k�[��ER=�}6j��x���V�?�I�;q���f�j�J�R�6�Z����sRbSc#��Jr��\�|������������ZRrv�����=;u#�&��_�̒�pչbcT#��4��<���E��$p�m�x������&�ɤ��C�H��+��U�Ľ"����a��t��6�p8en���۬b�Q�Upm��hcӤ�_��n� 	��w(r���E�K6Xkm�ЎI�v� ��!va��
�:7��"T��o�4a��)��͜9{����O��u�/�"|���}���|������aĘ����<��%��B 5��
GE["7��k�b��Z�	y'&(B|g�Z
��J�!��M+*����A���>rt�>}��������������?���ߎ�o���Ç<|�7�&����1s��֕��_#B���A2����D�]���M��5�헣9�,�6��Φ*s���(�ʊ�ҬJ���)�լ�*fZ15���^�H+e���S*�)���
��rnB/�LW.�)�(�E������"zd5���,��qn��'y��%�Q��'E��2*����/�=(b>,f=*�<.�W��P��W=�'?)�>+�>�#�N�����UvT1%���8�~��lmId���M<'�w`URkU��TV�md��Fi��XkP����a|#Dx:�͢G��Z2b����g�7�;b֧&1hƧ�>`���+�/9�lӅu{��������~��������������7���}�;����������:z��3����_��F�,<��N^�|�"���q!�k�2
*�޾�h��E&/\0u�©}����?�4eԷ�}�z��%s�o\� H�u\�K���<.��%)�\�"��@�5foߺq��U��MkV�-�3kژQC&O;a�ر�F�	��{�ٵ��È�Bo��T��T��p�|O "��%"��Go���vb4�V�¶G��v~���N?^t�I]v12q�=�	�5�]�_(҈�X�Pq�֣��F�7�����"�u�P�T�(�H�*�<#%ɨS�ٌ���#=z�<������S\�����~����g���y����V�a�`i\)C��f��)�/���Mj�w��������J#h�	�k�������9��z��#w��V\�Ħ��2�E�GYz�c����j��f#�ТW;M6&]�d����D�Y}1f��W�*�w}a��F/P��]����P���/�0t�nh�J�����ӗo�;g��3�̙6c���C�|��{���_���oA�_�����~�M����8w����K�|��+�s�GCg+�<9�+�Ϲ���!���p`0l.!����¨�1)\�'`Do2�>����;f���_~����������������_ǌ0jԠ��`u�w��>c�|6j����,)����C����8A2
�.T0DJ�D�a?%B����
9�g���v���k�k��Zv�ٚs/��O�?u��h�䡻����=�dѮk�ǟ|�u-�b��W�g쿓��n��{��g|�����ov�H�y���q{n��ގ�7aߝ���cw݌�u�ա�o�D�����q��g�A2�<� �?���$�Px��E��d��O9p/����g9�7$$�,#ɜd��D�A�cی��ӂ1��<V��fq�Eb��	CڱSӽ��[�%�
�n��,;tq���+�Z��Ć#������$pg������o�����>���{���~�uC'�:.l�Ǜv_߼��E��ۯ.�}��̽�g��=w���;W��N�/"q�2[og�l<�]��"� B(J��C-56�ͷ`uTq���̙6vԨ�/�6o���{7>yz��,������47/��8��Ts����̤��x����^Ǿ��L~���Y�("�^FF<����Օ�yYe�����K����x�����K-�>u��1+��?z�JtBN_��ҝj��DԫY;w�*��G��j�C"5���3b%V,�c�{�~��N
�M:v�Q�c�3=�#��26�"�	��UPxr����]hrt�^ L�7Nj�T�a�w�2%�ɡs8�=*.-�|q���T�T�jjQ�,�>O��(֛�&����\b�[l�����S$f��d�����n좧� Ɂ��G�͟�'D]�����]̷�F�"lqirs��s���&��F<^�ǭ�T�Ȇ��!���P9�S&��t��7a�,ׁm~Qq!��ok��T�3"�{jT���.B臑�>ᠰ3�o�5k��i��N?y�`�7}���?�����������j⤱�(:�?DF��/=(�A�|-��c�5,��ő�9b�_�C�<��B��*�K�A�!W,M������ B�y�Ǐ��7_��������������~7rȷÇ�6d tʾ4���?=����"��׈�a6X���B.�ΦQ2OW�E)z���J��BW��Qj�8�^պ�[�	U���
~���K�-�lo�㹱Fc;0�G��DnL�Ą6�Z�|&4a"3�؂�&��#p���ɼ�2�I�!^L��~�! �x1Y S�a'&v�s*��S\��sF��������k����R[��A�5����0��Zڹ^��ƪU�:�*�WL�y��˔\��U=��[J��.�\x?(R����?��z3�x�ʣ��o�}>fין��E;�=���h�����n��W�ϓ˟'�>O.~���U�QV_��~Y(�?F[�_� �L��|yP�N��#3�B�a�(mJrFB̋};�Ϛ1zɒi7��z�$�����87-%���F�s3AcQ/��$���T�9u�����e���]{6=~r;;79+3�����ݠQII	q/"#�R޼�~���U���}��o����O7�ܙkwD�g�T��v�:��$���������6��a��!����(��؆5��o���Y|;ن�i[&m8�s5��>���;���;b��D���t(��5rߥC��ކ�ܙ�| j� Z��ipl�6���h����	u�%Z�@e�gF�P�)���
�mV��.���f��d#~�RP`���:�Y��]�u���Pe�Ձ����,AJ,A�[UW�Y]��pI�N��#�e>.B�Z"tX�4�tު�e\[j�n��;��`E>,ێ]+F�E1�^�\!��!~yB����3'l����Ə�>~�������|��?������>_~�׏ߟ8q��A��~?DXSO�t|!��DHgI�\a�[����n��{���ʤqxt..�Қ�c���à!�'M�0a��o�~�������D��?}�_��d@�O���������W?<����'҄]"�`�lj���%D�.B
���+��w��"r�T.���R|g>��FH���F�zz���w��z컰��.�|��H����
{��n*P�'3�+O=��B)�5��zk��{���Y\Ȳ�X��K�e>��EGlL���W1��)e�6��q8J>_��85�����@j�ȭ\�Z=�\�+C��ė��
�H�D[��@��|t����xh�Ď�`[k$ִ:adn��Ē���!Ҩr��]�at;���s�q�����t�eұ��_�7����Na�ELL�j^|);��Ė�N<L�3!�Eg޶+K��M*W�	#3�Cg�Xw�ѱ�oM^�wԒ��[ߧ�%�Yu�Y5���^g��V�א8b��j�Pk��E�6B�*w:���n��/7a��<�C1�Ԕ�_���z���};Wo޸(!�Y|lxTă����Y�x����\?u��M�'��϶S'��ڱ}ޜٗ.�Y�d����&Ns���g͚=cĈ�O_�|�3gW�Xq���۷M?zŲE`�計7����;���¹�����&d�WP����[0�mj�ѧTD�s5q4&����eW"����/��چUZ1�[|�^�J�`$u��u��n��m�6z��;.��r�J�ki��<r�օ�D�Wb�;�:�0���Q��B5�*�T�R����u��un�+<� �F���x�f�jL�/y�Ae�Q��]U�F#:��5t�#��~�.~B�0T�~��y޾{����7kD�٣R*�BQms��=�`9�V�N���\��F�.z6^�/PaMXE+��ö>̿�BlmA�~D�8e]�����fa7B�D�w�!S�5~���F?�?��߷|������4�A�����>�z]VI�
�`A��\��b�L��C�mM���L����3��![$!�蓧���o4e�h��}��~�O��������g��k����˿�鳿~�ѧ_��}�8�����U�~5G�S��Z�@|g�zx�?j?pJq�RY�I2��lҸǟUp�v.�hډ+�?})U�i���G�-P��[&n��8��,�;v��L����V�w/���m��M���r�U&�L+����'�Eb��e�X!��L�E�|�J�ר�r�V&W��:��}*#�4���A�6�ƫ44�Pf�k���'w3���U E�#�a�%O��K���P���ˑ B��,����x�(�P�r��r��j���l{{��]+��G����
~L�e1�e/�Rz<<���������Ø2id��Wv�z�FK��݉�:p�e��+�+xIŴ��Ɣ��������-��� �#�1�[�V�B�t&�Ί�(�W���n��X�ʙSYWT�����;�O_�|Ĥ��5���o][0k���}�#"�?~������9u����wo��ׯߩ�'v��y���>}��s���;��g_�?{���S'���8~�㇏@�+�-�!�E�yYZV��ի��ήY����q�%EѶ���ζ:��S���ig+L)Ռ
�W�a�bۘ�Wc9�+���Q"r�\]�M[{X��.������/��i}B2M�w�okJ�'t��:`�u��z�ݕ|�y�F\a|S��D6��6�U�'o��G$��!�&�>=����-�Q��h4F�ڈ�:��m'��O!����`�[g�S*tY���}y��F��6��!s��.��m:+�NV	������r�o�v;m���a����P%p�TV�R-�j�Q�`��5"m�vD��ܡCG�4hƍ�~��/C"�u�\Mu���,+) <t��b^%���C/��\���цD�`�[�@~�m��V!B"�D(�v=��@H�t6���x|
�6y�ԁ�?z��a7cXkYq��|�?�����~����_~��{�����_��O_���YFe�"l�
q�@�;~T �?�T���?�
DD�L$�bD
�D�Cn�[�l�p+��e�(F�R۞+s'�,�Nl����1��ޛ�m��a+ϼ���h�byl��j�M36��WZ)�AeFV��j]meiL�A�XL��B
�\!Q��rD"{��U"�F�@J+_i�]\����p�>���N)��1mY�Ԁɭ�ڃ[1ą�U�Z�C��&Ű
�+�k�����U*�גʖ�}5�p���\�lmLS3�ࣩ��r{���Bh*�yTMz�2��]*�oм�Sm���w��4���eޟ�fʮk_��9��ݣ��/+��jً���_�Z�<��M	=���UA)���k(,2[�H���V�y���!4Lb�Z�����`h��p��듏ߛ{�ʊ��v�ٛ��(d6g��//,�JK�~����ބb����N:�~����nۺ7<�źS����8����t��Ĕ����u���%a	��{w�y�����v��}�ҥ����������Q��ܸ�����v/_�c�]��E�Vz�{��T��݌Av�Ȃ��yzo��e���x����̳h�J�W�Ř&l��ө5�r��V�*:f�V,n�Va�NE�I+,M��݌�m]tI�P:sz��,�H��#��Hlݼ�a��HV,���};�F|��ؼ�/�N܉B�ʴ���`����h��Q����y�Dء�w�+�����	*@� UѼ`��e���t�I�v��N�����nW ���g�7{\m��1,Xw��k�;�jM��Z����+���x�)3�Ywv'����kT��f�����}��#�aܰ�F9���2y��\��m�i+V.2d؈�c�SK�k�t1���yZ��S��Pv!~��F�t���R�:RÂ���̙�<�ն6��+�V,�>�χ������ٟ���߾���~���|����}�����7�O*�%q���ahOQ|s(XP��?)BD3�e(]a��;'�;�(�Z�������.�Ղ嚰)÷��ͺ�r���;6�Գ�ze�#��bM��˽��rN��-pb��i+Ck���=��z�F-P�G�(@���)T��JOi�j��v�4>�� Ul�ڽWW��DdZ��ܓ�5G��9�x���;/�_~�s=�P����Ebǆ��|ń���س̫	��
iS7#i�<;&�����5�Wwc��T��Q;�W��QʳeQ������	�5f�HL��veɚf����X�!�����D�1�mM�被�'�3���2���Y�Ϯ�4pK�U4AC !�'�~�Hm��o��&���4��z.B��)C�
��"��zAE=��\YTT��]��W���������:9/�07�8.&�у�S'�<�x����wm޾��˘�'N=�
[��ū7S��=q�<����[6�),(�X_G.**���NII��Kx����K����.,kd�kH��F~YX�(,�)�q�2T�l���Ф�ƌ�yl��ӗrj,�8�!>���8��h:���V�У1�o<��<t;���Tz1���AA=1�M���c�~�C��`���r2�1ό�J��`�og_���/9�$W�Ƹv,��܈ΒZ���&���Q����j ��1�� o-��$B�S���M��k�$U���{�-^u�W���^���;�Z�C㴩\V��j@t&ߪ�a��[�W���;o��X���<��X0�TǕ!R�Q��*-�׈0��h�������=u��	#G����'�0���}f�y��4�ǥ3�䅋����c�TѩBS��6�P'j$������ۼM�B�D�	_�t�����0�i����),7q����[����WV��1lѨ�}�~�oÿ�렯>����}�ŗ�|�a�!�W��x��WY=D��.~� (��L���e�UA��dp:\#\��%G�
+Y�������2iX�N�!-�b��yā'
鷨�]ߛQ�Á+�Ȓ|�bjږ�3��ݗ�Z��ml��.�
Dhgh�\�	?�!�h�|���Jp��n��J��D9J3Gm�.B�.p92�֫�"�9�9UT�l�x�\y��BP�3E��7^x
MÎes���`��?J��x���pb���7^x�sbk����35�������P�>�)�*_��[.pD��)���y���<�=��Z��x���+QyڶJ+��jɔx���t�-��9��h���	բ|����,f���J���-���j�H� ޲Y������s,�f*=�����f���b)�'N�+Rb�D�'�x���U��5��hT��-� ��S)4qq�uB6�+5����-��'q�e�:?��Z���dT�Q

�H$NM��Ăg�P9d*:gt� ���W\^]YO)�i,���ф$�����J,P�3dn�z�j?O�[�|�'����T[Zx-����I���V���N�v��e�0��O�5	��di����mmx�{|���5r�t���X�Х�t�ڽ<n��`X����p�Ü�'��Ĕ4h�ݠx6�o�:E蓡����*T������4��#��p��ŏ��EO�DX�+a�6^����]nG�S�s)<n����;:�Um���&�=��f�W�:GVJ�]����V�m�^f	�n��^M�@��%�U���C���r=��X��Ԥ��ϙ�x�ԅs&Ϛ1z����OKOy���\Q^XWS1c�ԯ���������UP�|C(e:UL�������Z0?��!�w��K��9R���	�~����ߞ9y81�eq^Z«��O���/��C���1��7���7p��ߍ\w�����\��%�g�g��!��`P��r�-ǯ��W8
=[�Bjđ�R7C"l�xvݍ�p5�D�1�X&�{>�n�ո����gnU��خԪ]���M�v���[��}��������c-�����EH�ip�E񺐧�s4z�Z0UZ�"�0Tz���P��j3K�_��E��t�����y[O�s�eQ��<Xt�j���dՈ�׈f�:_.wᗃ�b��^�����7�~LԂQmXװ�Z$E�囚ņ����k}l�:�T�EW�w�{�����g��9�p���oH���i�oYz����3)Yʖ�7c��OJ���%.a���@���6_O���P]_*v���"{��R&0���2��������2+[� 5@ʿ"����3k)љ�
�Oa�kM2k{�Pw �xӳ���B�L�J��܉~�]U���"F����Q$e�0S��Y �Z���̪g��H)�gU7p@�����j2��-������RJC��Q1e��P/�4 Z��D�[ꄺj������kk�Z�� ������d6LjǠ�&)LK�(�Q,M �#q`r;V@��]E�T80��]�R6�D.��grcf��b�G�u	5v�H5X�'E54(��2m9v%��#Y�7ٌ�|Qp�UT���%>�a�*�
.
�}H��ށh,����B~h�����&�VL�½w��V�JfRqPG���b�	��H�*�^�á�	X�H�[T�|�I�ܗB׌�~����VL��TV�nb���,�ތ_�R���������r�m7�1|̌�gO�b��9��Μ6jͪ��/�8zh׉�o\�4a��/?��o�?~Q�W	=3M"��Ņ��E����a�b� B�!�w��I�`q�)���84\�T���/9v�������W�ƍ�2q��)c�L;s�0���
?��!�:��a�?�vı;/���$�:�QP�ֲ�un�2�K$@��Jf��$z��*1��F�:ծ6��!(�u�a,���u֫ݩ��v����n%2���iG�Ok,�a�?=���Ҍշcc�>�b�Ƀ%�G+)��\X�z�����+�$�w������1�d��:~uP���31�&��X%R��D�l��}k�̤i�7V�V�e������:/[�gꚀ�Q�A�&U�<rwǍ��?��Xr�IEC1a�kq�Ǐ"��O�9��|�����{��f��<;�G�"��ڜ���G�v�$��q�E΅�i��S-F�J2X�T�c����㫦��ތM��_O;�,US=S|!��T=��'Y[o&>*�&��i\g��)O��x�����5a��͗�o:��^�;r�N��z�ގ+�7�����=�%�4��%�Q��ߩ�WI/�Vގ��Z��\ڀ�aw_��u"XxK��e��ep�T�
>I3E�6J�$��N���)jX�j���©��(t>�%b��|���A�L�K3p�f2Ǟ�7=��/3%U~]u#�w#�u�E8&��Q�V�J�U@���;x>:�����U���

WX�%h���
�ڂ)�D�k}
]@��uM��Ф�{z'����B
�.��E�uN���W���B�^�J����'V
�fօ��D���X6I�p�1��@gBf�BGA�6K����V(�����P�w�םđ�n��ez؉%�����b��ˬ
�J��I'���sؔ�ҢJ]��Ce���
EfFnzNŦ�W�됸d�u6LҌ��Ɓ���Ar�To��;D��u�M�]�O���� �:�{ֱȓ���g�?n��c���j����G�[�p�ְ5k�,[:�Y��O3b������;O+K(�&E̡˸,�-㲥L�Τ�D؆5"$�N�
���"�2��� B
O����xD8���?����w_|��o>��A���1vдQ�'�7vh���c�"\{���g�VPE �&~�Q��A�D�YH�L��"P��Z���}�ƅ�Y�6���J{��	M�����;8�w�yd6InnDuf,�c\�8m�駣���[Vl�RXΓ���$mL�h�R��C7^#΃�3/?{���z���/�U�+]kY��|s����,5��j�Z8��-m��E�cm*S	#%Bc!�x0h[�(G"�2�.\{���r6UӔ��^�'O�7c�/�L�j�ثZ�����n��d����]�"g<I1u���j�;"��E	 P���2$��A\��I�uHYSƷ��p�u��P�=Y��^��ĪmSW��y���]v_����7>��q��c�c��5ئ����S/�>/�_�|I�M���Ƃ}����vց;�ߔ�J�������TG�������K,�l�����XZ�-�R�0���R���w�=�Ȥ���N�{]ê�:�Φ:�is�1,��]u�T6�]����*���!���j�PB9H�
�4�AU��Ǧ�8Tc#Ӽ��W�<sw�ћ��Yv�������x��\�qa�t�ˑ+���s�YJ�D؆�	O�t���ȉ���-C@��ɍ̀LP�M�ڃ�O��Z7��:u:7�u�.�Ω�����9ʌn!�ު��S�·��j���˷���
�-,��؍�a�VM[�s߅��I`A���L`��"B"]
��qaO������iA D(Է�\sj��[QY��/��JˋRbc���ܻ{��?��bق���$�F�f$�|q�ʕ��?��:,�-�������3��̙�3{f��xB�[�F��HB�B���	���iww��n�P�.�&{�s����>Y�穧(�i�֧���>��"��Wx7c���;�w;�(��\���n�w�I��&�p�|�D,���"[�lt�?q�+�3���y�Ν����ڝ>����y�Çw:m������2��ܴ���z����f�G��X����i���K��[�"��P|�粼 �-�'3ʪ��q䥙e04� C�88�5k�m,6�]��������l�f�՚m�� [��Dhkm	D���Ӗ�����*jo#���,�QT����(���l��̕�yrG1�TS$�,N<3�1��3|�R�G�&�b#U��'x�)�||@6٩z�9�顷�w��b�B�D��:Yc��@4D�@��w4P.@�yhD	� ��Q������@�h�̀tlH���&ׂ,���R�
�LD�U}#"��m��B��_w4�'�Q��W<{�R��T�/�L���7f�����C#�hsP�:�&���̝�mD�]|��ڳ��o�kG@"ld�!�7��NT�AZA�-cK�t��&�d��w]���ٍ8��N�����0��g�$W=Ϯ�H���VD݉�{�W[?p�3ԧ��jDnH� ij�.
,���_+�_w'�?=v$�ܻ��[�H��\����·�^�,9�֬�����h�$}���f�� ���^�@/����-���cw�&��K�q�l)mf!���/�(���;3������4}��`I�0�n�w�?����������#4"�I!pIDVڛ�̷9�e%e��d�@#U��?}�����GhIf��-l#]�	��y�[�C�ߎ�&I��ZHe���i�l���F)g b9�?��(��ɥcJ�^%S+F�2xbU�Dx�(Bd4!rD���*�VSD�T'3����ۮ%M�����
�Iu,�
�s.o ��~�R�d(�/���~�%~jA !G����{TTn�3�GJ.���8++�����3ϓ�?�-+|����TS�������7]���z���cMC�d�r�{7`�m�sϢ��r�{"�#�hL�e���&�MJ�f���=����ꖋ����C���:u`��o�����TG�f����ژ[�"L�@��<�e	B�G�q��p��g~.?-�E�#с�G�4�>�'�)T��ϔ<
��a����V���h������������_���?}����d���|�������j�=+;���,l� ����r��\!<X!���,8���gO?��*d�+�ٹÒ�Aᙀt�~׃S���)��S]�}}+��Q=k�[<����7��%$?��}�=�ڳ�S���^�k��\{�ۄ��c��cK1���'<����b�5Ϩ��'i�Ǟm�x+4���{���HR�(Qc�ƨ��kQ���zѻ+�e^�=��C^�[N�a(�S%�,�;D���־G��@�]���\�����At9�V�d�tVA�QhX���~��Q����"Y�'1�$�,�$K>C�PUJ�������unA��/`�P�0��w�倄MG�������j��%�"�.'�~�$�=�TOsڂʇ:���J�3�l�JU+!�zv�
(��5i��i�N5�Boٳm�PH#��흀��P;E~�uZ�h\U�k���u��|3�����/�[�uLM)Ahw�~5]�1̾��{������C��\_�{�dՠ��\U�ҍ��w��v�4�u��w���a���H�����:lw��ܧ�cŔn%���J���´�S�ó9��8<�OYI]�J�j,��(� �u�rtA � L"���F`A�|XP&��ez�T�����ʋ@3<%��_!_9D(��Z��S��PΗk�fT��L��d�I�a��0�,ȗ�A��..w�ɂ ��~�@�O��W٪�7_$?+�k��H��=�hT�`wNV���gMu�o�hm���E��gSuufF�S���� �8 ���i��s��)��=_����˵�<��-����!B	W$"TN~�J�v܏�Vn�����@���p9�|�����ǯ~���W��(B[+{�͉IY�p/�b���$�&���T
�?��X�(����E�o�D8D��Y�~�����k6m"����}��߂�����ݿ�������ÿ�������o�׬ "�rp^�������ݎ/��$	�^�Xi�p�4�!��/�BI�,N?�d0�.f4�*�'�=�|˚(��p��S��y�n#�5|�Sp�[y�W�:�J�7��7��,�q�gf�jB��:�G6xd�����P����> <�U���A-��n�ܙ���nJ?Uޏ9}�Q7����ˌ�%3�fBJ{�������U�ɐ��F��UA'�D�4�4]9E�O��t�8C1�T��L���$Շ!�S�AY3�8M��]�t�� �P��]�l�O�@6�.���z�udm'o�����ʛ�@�I�|�T�x��$�')�������q��I�IL������P�p�*X1�%	�	<`����.�Hߠ��XAX#���2B�C)�V�DX=1vHW.���rA(0BM�w��
��m�Pi��#!tP��3�Z��ԐA��j�(��?��p�<�SOP�0FiSPJ+�uYO[?��j�uǮ�g%R��2���ꕌ�2v��V���tYRiS@TrHdlhDdXD�m��Aw����3//�B�uu6u������<B_���%���K�#â)4q��֣P��=!���ƎC��.�1�(�$UγE���q����	�	�	��89P ��ԢM.\�Dj�i�m�:��c{&<F^�WfZ�B��H�L��#T �W(��9��i�E2��G��,��O�g���>J�'��QMp��JhH�a��={�XwCagKE^njA~Nrrb^N�R./.(./|K#�)h�@ggee훼Jwl�71,�Ϣ�3X)<IM:�Oq�F�D͒�XR	[&�H��^zeD�O:ߍ�R�������:m=�c��v����w��?���~���[��m--ll�ߦ�6����,��&�,�.�Ѕd�g~.�,!�@�C8v����
���>z�{��cV��6VfkV~��W���o~��������B\h�o��𝵅�����m�}������n Bdf�� �ʃ�"������s#�w�<���^t3���H�O��۸�y��/e�������JK�����!�*�Q��\t�p�v^_��*�2��n|l�"��y.�6�S�+;�Ӧ��jI����o>ʨ��R񢠥[��LP<"�~����z4��`A�Ĉl
�0�v�F��^%��eŷѺd���q8Jᥴ��rKad+���i�z����:�;�m����gߜy�����6}s9���\��-W�Y���v��� ����Md�RɸP6D(���;�>
/�k���)��zy㑥�O�*c��~��Ē�^Z;����>Ϯ};�������-a͘}�"υe5�f_Vt߉�k`*�3PPi����$������}�v��"Z�;_$�P�K�(c7{w���xU0U���]�"�X��m�
˪L�����GXdTC��u�Q�<��A'�c{5T��$���j��vʳ������:���[��۵������ܱ��i��}�\����j�����GY�oBjF^�o�ǉ�{mל<{xρ]�v6+֙%gY�>��������CZ�QPO���
��%�@D�(�*!�2�D=�т&~\D^�F/���.��\E� dX=8����'"T!���O��2�aL"�1.��O��O-�8o���|��r",���	�faI��o�}#=�������ܬ졁��ں�ܷo3�Yd|sUemYYA~IfN9!J0�Π��8�I<�M�E3l��y_�f��L���$B��J4�t'�p��.{ٵ����gN�89�-��˯�s��o7���lgmkemm�9>�����eϨg�U�9<w��TQ"
��Y���_,x*c	��*j�1T��l������57����=i�e�������MV|��~������?��?��?�ן��+��; BKs+ ���.V�����R��E��)��g���\�+!�@$�ܠd��`@���'���Q(����ɧW�[�,���V+�"�%͢�;�3zT�b[��>+�y�3Qc%�y�s/o'���L��8��6�!�μ�K�����w+�����?H���o�U�;�҉��fz��^~��Eb� �t�l�y�ufJP�^HNo�HfP���bY>A�-�[e����P���͟|���_<8d����q�d��>��D�����A���MC�܂��d#��Ժ�$J�!�@�� ��(�!��Èvz#I�/��< ��;��O=H��j&���ݸ��{^��I��ţ�Aַm�&�RP��1�bd�_~m�#rUg#��G6~}&�V
u���+�QMx�5	�m��v<*��� �����)u#M��XTzj��[w��]����u�Փ���wР�}�x�G��NjPB�z�|rcޘB������#-�����s��o�����]�������ڻ�q��ݾ;��:����Gl�����$�����Y��ءL�p��PF�HG��A(����44������rjP�W����^��q����X�1�$$7���g$�)�j�\�����,s��K,!O5�$B�f���ੌ���q�E �d	��"d	��!\�\��P�8	'�i���/fq�����8���?�Qr?� �����I��0��ǖ3q"�I%�(d6��ari:�g��d��KbS(\��#��FD�	Ȃ�4�S2��2*�?1�O��7�zDx�۩#'θ<wd���������������p����6���w���la�=.������D�K���\��@D�̽�6"��k�s��,��D8B�"�@�}8bE�о���G.���5߸n�V[��f+~��O����������������?�~��ߛm���ߵ�����5 ´��n�h���0M���r��DEH���4]�	�ӏJ��-*h�w\X;-����+�XdP5�!�s�oQ��q��-�rP�_�i�@�jB�������w"�EА�;�S4���CQ�Ay�����:v�#��=>��:��C�w�^�g�c�ڙ�ܱ{O�h�~/[b����"�3"��۳���9M�h�^:q���x�"7�e�)X�%�����aj>�T!�}W�
=�;�G�]���Aѭ��/v{��/��B<"�C;]�����)(�����'A>.�M(%F�tB(����I��
��9z�������a��B��n�dm��]��/,�+㿋뗞��6w���S)�.%UG�p
�F"�3ug_g���鬦�~������>����,�ؐb���8.�vtR�P����R��-��=��A�w)���Z�t*�AD����o>~Vه	[���5ę�JQ��fT^���^�$���B���n���������<��ؽ��<pb��C��ݽ�y���.���9w�|�]W/���A��v޿w��ٙ��Wc�-n���{�����g�Y����k���:	��~n3^5"Y���ΡuZ1�־� ��ltV���'.BDZK��)����Л�gh����j����p#��a� ���H��{�p�,��+� @\���x G���1P���I��^�+8��z~&�E�-��~bA�2�-���k���@��ݔqtRś��{�DzM&P�A?a�j5nh���f���Ja2y*�`�#��J���"4�WE�P���#�q��!���_q?}�̹���?|���mNv���%"�?�Ǖ�Wn����7���`�/&����U���HQ8:*SAc
�t6
��,����J[�D�/��!��4�LA���L�ˣǋ�X�n�,�];�����o��~����/�ůW}� �U+�}��|����7]\}3�F��RC�c-��GțD(`rDt���U��z�z����tԵO1ׯ�V7`q�a@I�N��m7|v�p�����|[kq���'i;.&V�}R[����d"��8���}����i��>o!*	������ln�*{h�#�~�n"�D�xFf������KOs{��	�t�$��Qx]xV��� )�<��2,)3$!3<5!,=�a� �X�IGE�y��7*J��
�YP��T>o]#J_��ogce�y('��CoPܫ�ϲ���H���OZ�c�I�`�y��^�T.��H���"�S�']��͗K^u��m��|�Qh� ?���)����o�w���*>�vۓ�c��{��"z�.��w�:�d�T�f:����֝7�}��#s�o�oW+�b����3.zG\�x����Z4�<>�t�m��{���t�qw���-��+P�i�����Zk~v\��=;��{oF R�3(��0Ԡ��9�����C ��;�an@���3Ճ�½�[�^��r����\��s`מC��qq:r������7G�<��D�k��ȟ7:��z�[�]�Z���j����}c��qߵ��lD��Q��#	������A�yH46#�Mʴ�K�6�z��`�~����e�䫍,����7�m�P?����3��c3ꆈ����:
E��$��!��]>	&�-v����x2�@"3XlO�HD2�P�/I��d��h2#V�e�β��s�ޓ$F�v�*e�c(��}*Br�'�WD7�4�����?���^��Ȉ	*�J�IO����'����/��9s�t������_��z���[^�h�8ш��E�X�_.B��_��4%��/�����/���GG��9y�ȑ�{vn�l�h�j�w_}����W?|��|�{���m���[��T����#S�_�d�`yL���3`r?��s���GRi�Q&��.�{ݎ���\y�����=��������|��|���X����|�݊�}��r��>�cw��f5��ir4C�g�����|)�'dqEHd˰,��C�'+P�~�$�6�2����.�n�d4��ӫ��(�DS�NR�5`G�X	N8�N�-��Lt��x�A8����L*j�q�Z�xX�(S:O�vbD�ॽdEAֆ�7����@�|�<���!o?t��ݻO^lٵo����歶[�����u�`��#�.��L`J�����G�|�E�q�~J6:-�����C޶�V���PA��Yt�`b��O�t�^8�S;���!��w�{!�J`��D��2��1�w��,נ��&l%�[�I����B8�$
��F�t.Z����3��5�ܫ���;}'��iQ�ᗩG�wyE&��*�y8QBm�WX܋�k�Q�DC
f�F�U�#������ֆq�N*/ˬ�M�(�/Q�Z��:4�*%�;�Ek��7�O.�;V��s30#����W@�������v�;1@�����ԇN�|H6Ϟ�0p�ѫ�\��D����}w�8������z��uc#��Xom�{�����΀5�����k��쏿)�ñ�3��{�c�w��w�B�0
(�z��_X`Nq?�<'�L��[��Uc�-��j&2�ͧ�������Q�����29�b��1ZJT�zr��5k^�����D.�#$и��#=}�h4��d�(����֮x-'�Du/1��)$�2��wHdҪ�R�:����q�j1~��GE���(f�y����Ttw{}EWs#���s7P�ԧAS�w�_���w�76�6��d�8z
�gbE�$%DV/�"�M0�,�$B��#B%21�~^����q��=g��b8���m,l�6lZ\���oX���MkVY��ï��Ǻ�f�.gՌ����o��>�-c0��pv��������rc�%���I�"�eJv���wQ���e�����~���N;��[�������w+��Úo�\��+����
��n>��N3v��D��Ԩ|9���Eȗ�	�sx��0O*S��H�g���c#<K?+0γ��t���@d0��>M8:�M���T��"�#�0e�4��³D����P:��W��(�~o +$���L��%�F)�	�d
�RpQ�և�U5u\��0!=�mIى3gיm077?ppߚU+ �V��a���������΁�����n<�ėIG'�lx=G���ҩ���಑�D���T���9e�v�y��w��W)��1��;ē7���f�A�BJp+"S8I��j�N&�&I�9�Jo�9_�M���p�z~)E%�����z��罣:��ӞA�_%s�?�8 ��q��=�����ĳHۋ�	�>)��ӪQ��O}ݞ�Y8�]п�A���F��b�j3
��]9M2����y�=�Ye�W���(���ׁ/
#<z����{F>�}Rޏq�$h@�M>L*>����G�[t~�lp36��˔\��A��!<�͡{�Ex���=�����$�ۏp:��Ե��*�T��]�WnXg��a��9���Z��V�|���;�����������>ɻt�IU���c)�bR���	�v
$B�z��"�]�X��?�ڈ�[�|
�ٺi��x�yPTak���/3����sP.m�~I�퓈�O�A���AD~za훂�a,Md���Z[*��[�Id\{gG@hxTR&�)f�^��~ېֈ���X7X�E�����*������a�.��?5�G>z�' �Dl:(�M�U3'<#��A!���5I� f''�߼GF���8���2�3R"���߷���څ"ĉg(���L"42�&��׶\�¿"B���@,����a�ێ�m�y��i�������u�k-l6Y�Yl�4[k������~�j��Ï�]x�R>�c�P��>4�'�$L��?��Q~.B�Ʌ@��~�����$*��q���o׮�r�Z��V�����}��7��믿��[py����+�����������Ռ�g(��Rx�%����8���Qp�L�kq��'��A-C���"%I��rq\��0�b0�K�OK�:vVy�H/��,��%�Є"OÕ���(<���P"�$�.b	��I��P�Hb�l��� 
/�k�I�X�I
Gǖ%�Y�@�ޏ�	
)��I�|s��;wn�_��|㺫��89X�:Z;:ڏ��EUu�C،���
k[A��*�5��5-�խ��m��(V�@6��;d��q�]:A� ���cP9Yܯ�#OA(-<G%y��{�U��5�"�N.T�-G:>�c�z��ԓ�f��f��Y���Tٳ�܃>���!��7:�M􏎿��-�y�]�Dӌף��3��� �vy&�x�����-�i��4�fL������A���_��UW���<|x�qJ30���V��ڻ.=p/�I�>LK��Ώ���<��J��r�%T��!�

m����N�����&�w����F>kv���wP��7BU��OE��S�lu�E�cQ����a��WYm�Yk�n����V�ZZ����_o�߿[��&1@�)���l��6��N�H�!�\B;�����A�d����H"D����� <��G�}��A3s�;,��&!�ԯ�μ�y��G[��H�;���4.f��PE�?4:�U4H~ �u�WV�f�������e�.^����M`����|b�:��j��Z�:�v��w�JYe�"�G� .�r��"Ԋ�j�h�ɪ��O�Pҩ{�ݹv�ʙ��O�|�e��m�C�3מaH̫ׯ�����ǟ?v��3�Rhg���$��J��%�|DeB�)�I�J�DM��R4�'�bm\nYm;b���v�߮\����n����[�o0����u���u[o����1,��3���O$P82&})b?���g~.?������Wb�D�$B*C��e�,C�`���ʡ+�V[���߯����?��7�Y��;�߮v��ڭ����?�n�?��K�î#򎻿J����AP�q@D3��ˆG��� 1�-&�dD����y: U<F�i��-&��0d� �f�!��;*×*�Q4*�E��<��ǵ,�f( �+����) $���TP�*:SMgj=�7�a�c}(:x$����L�x�!�3�n߹�f����o֯����m gG+�+W���ˑ�/_���mE]z~ii}k� <{��R@z~yj~ei��Es5#l%2ܞ��'��B$ջa�Z1��o��;����grUPag3�����"�H([��0��h��>���෡��~*�Z�̩GA=����}�#��%%W�_>s���q�?����]ϗ���8{Ƿ��;XqԷ��y�Pva�������G9�O����x�Ń��g��LL�(͹v���[7����T���wVVfyr �.�*�a䳛����h�k\=e�A�kH�c�jЀ�@h����!U�dy72z@�:
���\���].�;�=z����]>{�����n=xp��S����q�,���{	�}��}��{����;Z�8X�����W����/�8%�Hg ��o
���z��ð�<u*�o���gWp�G5�4���^��D(T��j#W3���=��샃"�-�vB�����˧����=:�E	|�X��;[]2�@�_��!57�E&$$$��F�z��ߤFǼ��I)*̠Ұ=��>�}"b�*��*�@�{�h�v�cJk x'V�V��A?!2�c�?��/�܂�c��|�U5q�;������٣��S���r���x6q�;��Ŋs.x=��t��͋���>v��('�{��M�H�&�2~�ߢ�>��ܑ������S��W��s�=���>�{����O��7��A������ǉ��^�H=\��hp���	�,���W�8*&n�������¼�˲�"$��
Y���F��/�~�Qla��G!NGݬw\�}��
�������ԗ�g��xn�����F:_��h�9_|�݄"fɰl�-��E�E'�9e��,)��S�'�j�(\���s�L�
@�(H!�+����\��Q�b��B�D�1��X\�q!�B!�K�*�9*�Ĕ �]�XJK��hY|=G0fBO�)�)�z�Lg��T�ԕV�?�z��q�o-֯����k��W}�����}�G��o+k�14G�g2�]Ԫ<��&3��z2_	���A�dJ��� U.��:��+^��]�o���Ƴ=7_�*h�!�1��f�)�;�3� ��8�BI�Ƴ��:��@j�+F�٪�w�����}�h��~/��J\o\z��C�g5�V�u�����}G]�k�kG�$:?x�<@�����͹�������?�u���KMKI�{z7;9l� om(�p�����`�Я�����&%��>�K�/�}���%��HUC�~�XB��R@P��������c���\�)�}(�~����2��]��e�F����ܷcxcwo�w��Σ'lvp�w�����#�3Nݼ����������#������_�_m�/���7E�d4����@V����`���3�bs�S9�UL�B�␉�.�%�qx,�J+R�9Z�d���Rn���e�w���q�[d�Gf�7���G�n+6{��6,����o��������cbÂ�&&��򺝒~����A�aCy-0�6��F�WE��aE;}�����c�F�r�g"��.�T~��D��HG,B�ZDx�EA;���356���c�/����{�����,��Ԃo�����IOu�t��7�%Ԁ+��v�?�M�F�DO�(bC����>�j���q![���n��.��r�j��U~a�/_�yzgx��?}Y�<��'���u]pL{`�@h-'�Yp�'7��AѐDF�@��i�l5��`0d�E����B!Ӗ@���?!U D؂���@�х�~�eW�bN��>���$��W������/�e�{'�{��=�����Wa��},�G����	���E,Hg�R�j*G 4�P��k\5�!!SE"�Mi�{#R�5��1�t�kZ�PJ�J ���|�$P�j�W	\Hd�`����y_�h�9ЭB7!W�"���{[Pl������[�m��vl�;������r���?|}�����4*�-�狒�'0�L��V�A��RY�Q�O��	S:Fj�\5U:NO��:���L/GP�u15x�<Zb��� ���x�vP�$��5�C�ؤ��7���{ads��0,�O`hUuŝ�7��TW�e˖���<�ZV3\?�2�����۶>z~vN^N֝'Ϻ�D_f|��ztEop\2ᅓ�}ߤ�����.�r9�g��.aqIY����e4L/���F9�w��(&��&�
��̮Q��>�8,BP]/�Cˢ����C�� >�J�C���\���������$16�̹�>A!O��]����{�;Ǖ��*��\Fi���~�\�9>����k�]���d�f�Pa;���W7��'T��&�3^���%'�G$��s& �S���
�+�r�R��c� ^�iƷ���o��$����%sN����J��U'ɳ~�NI�ܸ٘z����_Skwdt�����k�l�57_������nn��y�]��?)���h!��:��֨F�ٗ%�%�oGn��us�
��&���VN�?�/�3�-�3*�b�R���4�|�p�y����W�I/c=b^�qr�U9c{?��3z�xQV[U\V���z��%�OD8DH���K��o��$B$n(j�xj�dw5��R��^����߭�����o�Ot��/���띿�v�oV��������kG�?�y��!���4^<A�1�z[ˠ�>��s��o�p�&�(y��.7�^{�aϥ[������wk�������f�?�������zӡ3s��{������Ng����&*Q�-�(B��ɂ@��ሦ��?��8!��;��jh*����3xR���#�\���т ���4�0|�:���"d�M"���	 "��j@?��Lap���b�z�������yy�߽c�#|kp��-@��f�׬����*84C!�����-VX"�<��� pb�cȴS<��d���fJဈ����IM�,�Ԉ���)�v�k���L�xJx�	۴"�G����afT�vT4���������N��IT���	����w�֑��r1x�/\��	��������S�'��U5����f�'߸s�Il�{R����̦O�����̤�3�vN�坍�7/�|��֭k��8ӫ��[�aI���u=�����Ԅ�-�W�%���T:�%��'����囫q'�:�}�|�s�uϣ����_R��57��Е���&�p����U�k�D��TT1�!�`)Aq�E��� H��*n����O�
�r�y�Dj~u@d�5wߚS=�ֿ{�2����4D�A(�L~��?���1��9���_�b�A�E��T	�P�R�}�Fϛ�F�F�:�����������Î=
��KH����a�]��y�1����3�IJI�w�������ds�����/x<���Ջ�7��*��P9Q[O~�ٙXK��A��)՘���~��$�`+�����'~j���d>�K��|�[�S�2j�T��	�����`p����*�����c����&n?r�������v�=�	U�=�G�F��I5G���-�h�� B-K���'i�P#�}	m&wH���Ϯǆ�V��br���-��.aa��M+/���W��-&��K��
1�V�(^<E�R8:&K�� f@�����w�E���B��hK "��Ȉ�D��^�r�7��	V�_9�\�(,��؛/�ne]�M?�}7��5����{�E!��1%����&����"a�M"\l%�T��ʒ�
 ��0�*�G��z�H���B	O��J	�%2�
GO��p�����Px!_�9�X�8����<�^)�#�Ehj�?�૘5`����x`�:*���108dϞ=�֮���������N֖׬_�îΑ1�z���`��S��q�L�h�R58����A� G�B%8H( p�-OF�� �n>p4�?����C����^�#��WT�7��f�TF�T��4y�#h�.��k

�q��+<VmMEUU��0�e`��ghZ1���7�oj���b�C�=�����?M.K��,(���{�v��'�Z4����V��./̾���L����I�z��}���S[w�o&
^&�Nh!�h�`��_��\�Sؚ[ٙUݞUӚU����U��{7 �LA�U��9M3ϐ�xb�H�rYL6���8�J�����3p�S �j�&��4�%���a��Dj���KW��	�j����kf4�,U3MUM��8*�" "�E~&B� Cdj�Ψ2��F��w��z��UA:�Ie���U��.:��12��h�q~��稍�d6x$M�b)�Q=���ك��q�o\=��~3���QYT�C�;�.���?�R�S��L%|;^C1%UN����|�i88�-�����T�ȇ�G�5�ٽ"���=�,�_1�4 �������G�m��8��d�H\ޏ5�����vڹk˖-�w�=~�B���#�!�(V:CP�,�G��'��5K,Y��� "d�f� �nF�Phw��iByY���ڽ�rD����	��_����������_��r;����׆��*�!���
*M�Q�H���"�\���G��,PZLI�È��O�/{'g6�_�չ�|�ސ�B���ޏ*{�\�,��ad���K��!Y��4eU�K"�\�K.DD��r$z�T#��A��U�H�(��Qk�Κ��g��12_bp Y�-C�� �Ј��*2Kaj�]t�PDS("�Caʫ�{�[�=<<�8ڂ,���~�V�%nX�þ�;�j�H.%ИL��S@�#� K��-<�i�x��s>�P����ѹ"S7Z!���es�\Sa�Ӣ�@����LN��;������ v:	��������}�ܢr »wn�Pު���������7n>���(B�Q��Lr}�PSII^zrPHpji���»�Ròʓ2��{Ǆ�x��ָFL�f�ƽI��r�-�f8��+<)=6"(>�i����\�=}�K}�5��Tp˘�M{OZViiq}e}[YC[YcKYcSxrrAm=M9:"�	�>�u�  B�D$��B�@$��Z�!�#0��(r�9�b�b�+�xy[�(K?���4�<���� �J#�-�t���Ɛ�#�n�b�]3/��� ��i�����8�^�p�HykS\~����^6�nhD�20(�����3CTR�P�pTɕx|�X�ii�.+~32�H#�@��:���:4ě���S]C��H�r�L/����U�Q�	�L%Q���y&��L�_�tq�����Ï"T�S��O^�HǣSs�(4�@��v��f�x{�P�oG���񦸶����ŗWV�EW��]�x�4����GDȔ��3��۷�KP���c��/<K�E]�I����}Obʙ��k�.��"��s�}�BҀ�FLӚ��YM���В���D�Y���_/?!�(M��^�<��}���E_�M��r�����%��i��ϓ���z��+~}2.��9_��<�(��țI]Tɒq\|�7��il���r�8j ����"B�TǓ�y�Be2�P���Y�&k���hl�ě�c��!� T��iE_P)O��	,�@�ha����d�P�U,��Mf32X�#��79)�~/���B.�;��v�f؅;�: "4[���8/9)���1�mv^aQ��0�/Ҁ\(S"���$rP���X*� ����8<�/`�
��a�m*\6��e
80`��B�G���C�&���׃!��l ��'K��F�C��7=XZc{OQQQzjbNV:����tTTT�ԶUUu�u�����>=�U�|__{]UfvV]!��3,���e���);#��<��8kR'���M5��Y)��o�Vc��}�ƒ����������D��PV�<+��TLS��̺�а��Ш��̄t@: 29������`���=w�NAT�U��J$ ""�p%(.��+t&F�A`�)���?�6�%��%C�*G9j 0��xд|Ҳ�M�&�B�,Q<V5��h��Nfp�Hހ<�	�2%1�0�ӥ�Pi�!�Pv�����ܶ�̚�H.�r�l���\~UѓPo턆�&K� Rb�SCg�er�Ì������WC_!�`j�;����g+��
x�D�T5.Q�I�zX�J�"����~���tp)""��D(T�D�QX�����O�����=���u�t�b�Zde?[��{��5��O�?z����0]p?0������3Y��@VF� �]"��4
D�N�]|�|=��[u(�b�!��X�W\�]�}�YO�z������_�!�"|�*hAU���7Oc*��"�+�c2G?7�~.��u�h�!�d��v<~�i\a+M��NI���t���\w���G<b2��N7��"J�E����ŝ��N�4m�{����w�\�_!H�@���D���%��?81��q�d�$�"
����ǃЂ9��#)p����6��3â�pf���q4K"$s�$������<9��#)mM8��+
~��ɓ��<��ٶ�v���9p������U@��Ea!�u�55U��x�-("S�:�Q$��2�@"�<G$�@���<������$b�@��	8��rXL.�(��E* v!���l|Dh��
]���ZcY8���ơ��P;ŗ)��R��V�QPH$�fB��W�hE	ʮG!>�*�q�����ip��C�z_��Q�h�H778=�U��F�t�M{A�9^7�/��04L/?H��L��e2�b2H��6(!�����N_�z�����coo@dRbam-!V��aD2Y5�"H'hRL+	%Ӕ� F���"��j�JCQ��1�RO��hr=!H�E�L�	����~�*��e���}p�c������WO1���UǞ�D����f��E�|�u�#�un�o�ߛ�2�W�8䮡�ھ�����y�<�DFv���)���$g��R%��!(�l�p�±����I!b.���4$,��%('����-��#(���I�΅B��x�
ܽ�G~��\�܂�"D\�q��#��@��Q#Sc<�(pX:��[���66:5=%3!6���9}l����8�����7�N�y��ٝ�Ooy>��]��o�r:h��D��M�j�l� �|�/�C0`��G���9�]���Xq+��5���VВ���nb�� 7�#�|2��y$4Ɉ�Y����L�?v�Y�H�w�,¿�|*B|yY�2�����ջN�2�͌ј�Ȫ�G��m���^�����;����]��[�8���{t-A]�����\�fb:�b�W��Cb`#:G�Q������5�a"o�̗?��5�����7b�{��Zh������2�*�xP:��P���!�J���e6�HJ[Gb���L��EH�Ã�q4>��*_�%Ҟy�|������-����~����������/���?���/��/w���^���iYYY8�D�$b�LH�<� ���'�4ոz7I|5�=Jajit1�����%�C&��f��T��P�b�H
�'3�F�f�i��cH,�P��7w�g(��y�H�F�@�"�d"�F!3iL6S�f+�|�#A9EVAjQ�
!_,3$�t�(�S@���AE����D(��B�\�^')��R�g�X$ H�B)V"Q��ӣSs�L�8���������;|b�Q��GO����Y���m��"�h��ЕX����Rxܘ@��`@��%Q,#�e�I��;��4Q=J��R$z��5��/� pk��'5�c����T�#c�>�(�����r>��7-������롐Z劽�r�R� �"	�<T\W�,��7��3��	�$�1лy2i���ws��Ҭ����1��`�;�$<Bf�+ha�����{	�^��#��悋H�bk����4��M�Y K����2bQ�2Lհ�V,����
�\B��هAT-�E5�����
��*�sjZ��3W�rX��LaJqudFn^ym��✪�A?<���#�������7���+:�������4��AD�Ɍ�Q�Al�˒�f��RG�Qm�����[�X�CP�{���qw�k���2��)�J�T;��4�/��yD���Rx��|�͔��4fv~f���{h�ޛ���|��U~Q��B �a:,��N��q�v�hglǍ�fGo�?��E7?�X2p�?s�Mg��������%�0���q�ͧ�6�E(�(Aj�
4X�ϓy��2t�lI�������E����SP� m˝�s1�7�ڏ�|��4�(����'��7��1d����Lm#e�L��q�7�mWc���u�=VpN�s%T&��M!�z{��3�n<tw>|p��������n�a��l�}�s_���24Og�@ٍ'�<���2	�'�
��R�=p���(���-����:�@�4Ho�^��0:v��駡���n���j�ZY�*v���| K/[a�����L��"T�xj�4�RZ�]lT������$,��ł��b��6����X`\�����-�O�34��� hx�:.��cQ:p$��z_�a����T�F�S(2�DYV(H0TZySkr�������7�o@z��*ȯk�"00|%�������*� �tq..�X+���d+��Q{f����A�����~�&��+��U����hA�
�;���?]��w�^,���WW���S�,���.��n�J
�+ )YD!U2&{S��R������P��_c� "M��4�Q�=N�;�Ã�4������Ę �P�������l&&7?�}���u�+�F竾x��"���b�HV�hA�� |�P���	�%"�(��,O���hA�ƕ�$ʉ�KI� �ĝ���I���j4]A�1�Nv�C���\i}Ϡdr��-��)�R-C=���C��"���n�JQ��/��dCJ���܎{	��ݍ���FҚc�N{ֳfV��P�TK������Qz5��2�c�`h���5�nj���g~.?-E�ڢ����}���œ�|C\���N'�p_ﺐ���9���<�� ��Y������*�!�h`��!�Lo����HM�SãݹW��(��Pd"�%(��e)&�B�gD�ĂV�s�Ϝ�K��$��\}�<{�U\XGӬ;r�T�jd���n�ݠ��a�4�=Jb(��L�<��ǎ��jʁ M]x��\�2��j�@Vߍ���]��<�o҉����O�]
Hz�:���Ԥ� �� �Wx<M2˾��IX�P9&�[{�����^��Gmt�@f8�$[�+�[�XK(�;��ā���ʼ'����>~�ɋ���--=�8���
�P^}�otzxbfLBrbbbrbBJ�MJHL�K��M��N��J�IH�J����N�N�����~����*�u�����/�B��_Ą�D��F���DD���g&���O������bcB#"B�_G��&�&g��rc������:|r�c�{�������57��aEO�R�#2��g�RX�)����+3�9�T�2գ�I��Ĉq�T?b4P����`l^�Hb�E(�	%0�vp%���X.���u�����{*f������rЫZP^A���"��.��R������/��;�S�B��x\_[����3b�^x�e'v�V�g'ܻu���½�'�K2ۚ+#c�=�2�����]n�2=bA roO�����W!���iӮj�1��IsE�s.�P&W��jO%��Ԑ|ʨ8����$jTO_	Nh��� H�z�*�����L�K�]�|�jG��~�dD�$+ƀي1Sd��;@��9�5ோ( TJ�O`��8Ż���I���|�^_�W<O�{]�[�	�_�K��_|���|�A�m�7e��f���q�04���E����"�\�b��K��F��p�.�(��z��8z��o��[�����x�;��B�%*�*W���P��x�{�W{om=�8�z�����(�a��S�9�!W���\�3:F��4Ie7���لҦN�\'��;��}��Z�b�ݗ�U� ��wP�d�+���-�����4��������n�8�i�)� x���,��"[Lb	@($�y\��Fd���`�����|6]��p����󣷞�e���'���g��i�f��12U�JOW�h
5Y�B��U�Dڹ+��L�ϝ�H��OjM��L|��` ��P��������䇀�ć}��	����c�="���v�[HT\�0��6³o(��^���b�����������f�֮]�r�
��+֮\a�~��/׮�j�jp|�+׬�a�ʕ߬\����aݗ߯��ۯ��������~�_����U�����׬�~��U_�5�Xg~��u�֯_��l����7Ym��l�}�����Y���a���*+����+-��d��F��ֻ��s����ӟ�ۃ�G`S9͐�.d+�ٲ)�j�"7��~��A$ͧ���	�TF�D����hg��r�H2&����P9C�ͷ�Go%��z�f�\>t>���Z�_�[�ZF���*�aaF>;�3���y=�w]{�G���\��=}����[-V��:��~ù�{N��yә#��;[�n�i��pv9r`���C����G�{ƒe��BjI�,��#�pU�j;9�	x`�b\��<� ����Q�K%�?���	�D��I5R�F.�g�O>hb(R�	G�Ei<l�PRe�Bnnc�γ׺Ȭ>�er&�0=,P`%���P���p��X��L(�'B��c������	�B4_OӼ'�g��!�Ea$3`g�7�IS��~�XQ�l�IH��deJ�MV�R�����j2K�E`���W˧�M"�S?�����.Dqe�lY'I_X�2�m|IcE?��,�|[��0Ё�D�Y՝�U�5]�-i%�u=̓�~�&R��P��W�(�X���4E�Z.B�P������Χ�6bY�L^5˜��d3�)��3���G3SZܱ���������F����s/s���^�<��MCX���T�2CD�g
�l�%����&A�o[""DfC%�x��~��A巐�xF�^=B�f�`8-x����(�����B#Ě��h��F>A�g��h��j��X���2487'���mqmo^6�=��ħ�%�ޢ�ܢ&�%ō���*�G�����Mx~#����K���#�c�>z�"�XrW;KSL�;{�wߛ�4�Zʚ��*kV��[�z��5f��Y��`��|�s3��-,�:���ڬ�h��Z3�7��7�^������o������޴aզ��'W��Vm�\��z��Mf�l\o�i���6m�6��[�ml�u�h� o�����fs����N� ��`v��ڶ�q�wx
W;�2&��.0UL=�2��?��Ua�kl������ÝO^<��o,O7'����3r�L6&���e:d=[D��|�_�G��������U�C"�g�v)	]��&�WT&S��KEd>s
z�}7˛���S�P��_w���۶�:�{��;6�ad������lFp��xx���=�v���fcec����AXZ\-��U�T�i��TR�<�@,H)�"E
�3�tʹ`MB,�{�z��y�V�8�i�fٌI����E�<����r��r���.=
k�ɥ�Pv#�ڋ�3�D�V�k#K�=z��6Tރ�k'b
���2$�X�� V��j�T�����M�J6O���+�B��s�)B2�	��>�+ܛ<l��T:
����"=��%�48�
�V��a���G��0ep�t�̓g����`�Q`Xr�i&)� b1���4:�~r�?����"D}!�j;�(B�Ô�^2�	E�"4���XZ�։��XCD� �ч��1�,Ed��`$@*����MDDHG���+�,cR�ɂ98��;��ݗ$���f)SP��eHj%u��\}��`�RP���n��5#WB�n�r#�f������P8��Ȃ;��PHdq� �)���\�!� �4*<���1��"����k��d�ɚ�j����n���C�Ѵ)�>=�����>@Y��/�/Ħu���B����R\��H{Q}�%��Z�MwCD� �0�@K��/|N��
��?���7���
	�y�!x3AD oG3�r��W�Y�2[��������a6l4ްr��UkWGnX�r�x�~���6�۸�f�W ���l-8h�a-0ߚM �M�@��7ZZ�Yۂjak����,~ickiggmkccgge�`e���~+�d��,� ��'������}��AT-D7B�o��4�?�+��3���f�a���獾k椪I�r\)�����E73�T��-7�j����V�5�mV@k.����Pv7�;:�"V�l�� +z����c*{I��Gv��cw�oQ�����vo5���n�Y����-�/|�����J�����*�|Y;���U�H�)������d-��h��b���tf�S�#�~�c�#����/!�l�(����}A�ȦRH�����fH4ǟ��+����vV0��*#���Q��B�iFC%r
3D�+�Dhj���92�B 9�L�T踦��
=<�E
�e
��N*�C$Ҧ��rx2)Pu��d��H��h\��2��|,G��	�	N ���K<G@0]y�����Y���?��s���ɤ�h�2L��q!ȅp3)�?@�t��(r'�
8@d�ᙽ8����p�-����~�P��T:���Y��4��
UdD��A��.����Kƌ�@���v��y%���w#ʙS�y(��w�i�a��ץ}��շ#��^9� ��G���8����΅l ���$s�?�����,,��b0Plq]y�-�iJ5m�c�Ɩ�UW���<yU�O���<�}U=XJ�����B-���x����;�w�_K{q�.����H�CT�#L�cl�#|�Cb�]J�=A�SR�Gm���;C\^�k�����畛w���S���-:r�ޗk,V�Y�3�Қ���� K+kK����b�Fss�k��k֮�~͊�@|ܸa��Fˍk���;ژ9Xm�ڴ��l5!8na�� ����,- ���`nm�8�����
T�V6������v�r�h����`�_l�o�[�D�C�	�IV�gQW�j�@̛#)���34���i�i�zV�W)*�^)���p�P�/n��5�O�x����yj=_3��rJЋ���e]ɽ,{�`���\dIWDV�0�ه��FU8���#�M����$�ûM"�k��f�- �(Bk �?����j�O@m�ⶁA<���;#�Mf^>�/�{laeDiGt:�����-�+X�J2�L@
����0��wc9�*�n7��� �#�y�Y��]^�tH�5��n��>g!���N�-nk@sQ��v��UF!�($��9yi�+��| �Q"ӽy�����TS�� jp���KXB)G ��i�g� [���r9|��fq�L6��$S��"PiD��b8,�M��. �g�|_D���>�����Ih�?�O�r#��Xڢ14X�K�Y}� �9B��X]#�ne �:&�B@?�ۇg�P�x��	>�9�d�0�QD� Ăd�i���"���%8��{I�~�����Dswx�:?���}�/w�WJm�Q
�<�(�h�|h̀k�c��"�Bͬ����w_����ٰA��`��N����S"_� �xD��!GR��ڟ~��4u�Y�J�)����6
��]�;5P���0�O9U�Z�p�M��9�����3�O6������x<��0��0���되��-zN��"�~z"��y�sNy1>ﻝ�q� ���𞫝=|��+7!"4�uN[�l��u�����j��;oٽ�i�N���7�9o�ݱ�n�����z[+�-�V{��o�F߅�ha�`���M�� ��-�6V���m�A����[kK;X��EB!"B߰$P��DX DH�C�I�ɛ����)h����o��1��òY3M5/RN�,��i�R��T}�Mm}�,�X��Ă�X!P �_�����۝����ϣ�}��;n�8p�+���u`�=,׫�*ij$<3��'4�������n�_�;;�=�w��C{���pl����vG:�o�����{������d���b��-�˂.��i'��73�Dv(-=�eH�/ "�K�r�k���'�߶���������$?)1�8���?m6�\O(ej�-��e�1 B����x���?�}�3���(h�3����2.<
9�(�����S3NU����t�ǔy�D��̐QhRM�f(���!�-�ȍ�(*B��&���"�%xb	 � K�a��E�`��L��X!�����x.kI�x>�(��!@D���L"ļ���,����Ҫ�  ¢�Ehr!�*XE��t>|���ч��2w��.�pA4D�D`E �o��
x!2;6_D�d���<��E�D�H5$�� ���(�X+{�'I� �W���GT�œ�M#u!E�������u`�"�nA
A�tM3M�J�p$�4��/	�~�O�p����� �lP��EXB�K��A:��h�qﵧÒY�{�:��IhP%w�b��Ih�{d��$��}ʙ�ƒ���x/�ӛC��}p�=��`�wg���1n��nķ>�<?��>=�w0�^����O�\���y�6��=/��O�����J�v�.���o�Y�f�Ն���6�1n�.�=��!طc�5�W~���z߮m�l�߳��b����A}���n�fKpd��-��mwr�ܴaH� �Fܸi&� �L\�a�z3��ͭ,��VV0�����H.�K"��Ǟ�&�&���Q�Q�<�Z���g�U���D��K���C���?Q�0��Z#��eR�N'��R.�;�S��0���>_��⩗�s4�p�c�O]�P���h樺�Qx�d��J�brj���뻻1"[�@UWYl��S]ڹ����K����"ܷg��ێ�Ex���C.�v�2���w�%�'�}�+�7�����wc���PD^Mwkݸ����;�n���a���y�t���.ְꕼM2G?��e�z��ЄƄi_bj]�� ���t2��OD(��9��-�7�����7].��5�g�j�����SO��	��g�����f�J����@��+W�B]81D1l=�?�Y@�d=��'�yW^d�	I����+l`:�:��a�����H��	x!_(B��`�r��iA$�,��Ε �{��bp���V(��ã�xr�@�@��4\%,B� ��E�07}@D��X	�_]>���*�E8��E8B��"D "�8(
�E��҃��R�ȕ�B��M��"$�,��D�*�f��� �8�}��s=��F���"����{��lmM��EI'z��.�8��'������=T9A I���h��.BSD"|���4��� �Tt�WTVtQ3{����^g��e�ª����yU�*��>���@tԡ��q�o����J����q��������'�7�I9OHy��z�KjQ��Bi�P����[�ޗ�=���o��拧���Y|�~��e"ܸi���5{�8��v�e'�����V �ޱń�][��6��������ۻ��-��>qh�у;A@\��;�BD��yfk��fkW��E7�.4۸�n2�`a�����Q���G�b��s��'���9��7�#x�[�.<{��-�N���f����y�<��X�P�+�
�T����r�I�zd���Fi�)�L��G�Ģ�`�&��g��9��i�^5K�O��$eu��ၕ�0v$(<�yH�ˤ��^����/<��z���^g�m��l�;[��a�o���=V{��8`���r�,��a�n�/l�|��N��j�
Ny[S�F�-��7�e�8}E������1F� 	Q��xL�H�L�'DV��)��;�?��g���"o�L���෋�4�4�o6��'Ex���~-���y����rZ�˩�7����.4WG�i�1Ă&���^���lh�(!������o������OK��$�����Q�_ƀ���\��+� pD��c먂+R�	K�B���k �7p��r �^�[Ay2 <���g w�1-��p�~v"|?o��g~.�F[���o�rէ,�o�,E�����iL��Q���^gA�@�0H�TE�3+.=|z�������q��{σ��ѻ�m�p+��߆s�֜~�m����2���gu��沷�5�m7|v�����w������[�^��x�ΓM�w#
$2�0�hj��M͡��T���2�.��M�m�-+o�����m����.���I��ʄ�!�8TKV]�K�����J��C�L��
~�y���ԠgIO��E�?�}�{c0f(��7�ns��μ����龷�=·�=un����k@HW]o��ұY�$�N��cf�j���&sXN�Dx��v���vn߼u���6������;�"��}�%"�#{�۷�z��-H� nX��冕�Vf&�۴q�G�0[�r�U�$����j#�t�p"B Bk[k[�MD[�g���U��{�%*g���⣠����N����פ��m����;�*˫�g����.�"�&A�� ��J�T�P�,hIT�:}�F.�;@�@{L�G�:�JԈ� ��ˀC!p!K;��e���%z�z�Kk�d����#������-�y�!��Vp���O�ڴu������������W9ح��_�yӖm�N�m ��VΎ������|�ۏy�փ��yXbuQzOEjk������`:_,��R�'!�4��:X:�r��2��'&�j�T=
�eZ:ꧨ"|���(�\7,^=(����`�f)�������1-������{����2H?@%=�-�o����5�]'nx��T`XR�XM+aDZ�d����;�̓��T9�\:��-y��g���Bs�E�P`Z��s����)"=C���!�����@ ʄ'���,��dL4�J���t�OU��p�\�2�M�8��/�
(<�2�pv��?����"���ɂ ��>2���R�XQ��y��{�%D袉j�*���5�Ο(��ӵ���^1��?��f���u�uN`A[r���ԐdY�n��A�Y�E�t�ǂ[TH,ђE��R���G�DX����D0�H0�44��I4�Z��"�4�N�C�},9N:��ђq��d�Y�ЈdzX4E��6a���p�KFtD�����<�����ӼϦ?;��u6�əT��)�O$<>������	����8������n�����-׫�Y��A<K��㨦�_���f?l0_g�v��z`�];��ٽ�p���@��v:n�np��'�N6G\�;o�����'�[��X��5��z���{�;nZ����U6�m-�a.!�77[���Y��_��ޡ����&[{xd������x��ց:	b��_gU?��y�[�-�j�Rf!�
(j��i�o�r��gi�����r�G�	fi�BńX�[-�O�eF�f��1�tF�~@Rk��ȝ3��py��j�]��L�G�y�)P���p� �w*�*�&�͕�ԣ�<��`z_p�ֳ?�9|�f��5+��Ħ�_oZ����?��f���k��~շ�uk ��?��O�~�k�g_d�a����B�Z��k���:���S��3%�=C{��~���ʳ=�<�<z��7�3��r�nL�1ȵ�2��$Z�&Bx��L�Q�M$�!x�K���M�W���V��ܖ�V\�`T81���=�v�e�V�2Pۍ�'q�C�Ez�R�� 7�Suf�CEp�'�F�v>Ni�j!���}���FS	��3�(Ѷ#�I��x�$���F�x�*�#s�"��\��j_����l�i�z����ɤS,���͂�U���h�\�H���~��g~.�P�4�EH�E�хKV�o�D( "D:ːE�E�@�(�(��%"��,� H2p\F�L7�t&��f�h�������?��_�������_��=}��Ѹ���=�`" A��H��t��w�C`�=H��ہ��\��WB��}M�xj ���I.0��p��o��0|/SMk����A��z�x�$�W�!������'.����v����׏_�}��˧N�9�z����~~�w�޻�z���ݮ]�t�y�ԑ+���|��.�=NgOIKOij뤱�,�F��bH���\���k~Xk�v=l#{;�m[m�n�[�mv���;w8��#w�Yop�^w����[�7ۮ['�Mv�V[���|ͷ֛V:;Zښ��fo�c��f;K�p'R�a�q q!ҡ��r#��j��6�V�mC+`H3k[3+{3+Ǖ��Y9?�eig8c������P9'�ϊ��b�$@(��ɧ9J��>��fy�9`&P�#͞��Kx\9G3�����Gg�x������&kf�ƅ����;:��w�=5�UEe+��Sjr�	��T�8�b�/ɧ�I��C�f<O���j�G�MS]K�|�x^�A��&Z	��ꞻ��.��4�HMK��.��ƨ�  ��IDAT������oٶߡ#�O��{��i��cg6m����zci��kG���<|����젬�m����7��n,-.x�*����WFx��a����1��!Ň�|��"��
�~T���F�H"�����2&L��;����g�9_����ӛ�p��j��~G5@8�<F;�#J�t�(w����c���*U�"	���ɣ0u3���-d��Ƚ^��WְG#*OǴF7�^d�o>�׭�{32����%�r�A�uP�=M]r�"#ЧP?;B��3��t�Y��/�������,C ��Ѹ�|`�̪l
�YGՅe8
x��D���{��g~.�OD�_Q�"S0T��ǅ��e���~*B�P>��!"$�T&4�^��A��q|:���)-���_�ÿ��\o\�~�8$�����[JK0d2S(��8#T��;L|� ��BƁ�I�{~d&,Bx9@���Z i� �b�h���c: E�@C��Q��4�\E*d<�
n&R����ȄR4)й��ӍH$4�(xIoJs���S+s�+���R�/��n��Zl�����&�s��%�tu��4T���tww��pp�I@�,QN�Z�����V��_o���[��-����6n�b�m�H'��۱�b�v�ݾ����|�͆�V���n�ݰ}�5p���z�����mv "�H�զu Ă�Y�@��V���v,~Xo����+(X�H=+�O)%F�ب j�A!6Hd�[|�<W;�VO�TF�b� P)S;W5H=��?�����r�Ex^7�Od|�Z���y�P_�S������(5�Ձ�#T�
�@\�g�]�ԩdQ��G��"�V(Q	�
�D.�� ?�PmHt~�ݗQa���o��7��u����㇎�8t���K��_ۿ���Ӯ^^��\N���m*�x���+��c��B��-�v6T�c��F��j+_��~-Pc峥8IU7 �c�A�ihl�MLI�5�\#�W�_�I{?�'"�'E�i�d$f�� O��c+��� N@�����y�dl���dr�|Μ�1�F�ؽ� �@�Zm'���`� G���)<W������f�{���K/��ߎNzR�s"��������VZUW��>r'�w|#I����y"MB#Z��3�^d�Y2�$T�h'!�@O�P�c >25G�����:�(��Kg��J���F2�M��d�]1�RL�Ǒa�b"���?�O
�A_��my%"B�C��Do?��!�.;�E.Z�4�bAS���"�ߒ$J E���$t8��f �l���W�����Ҋ^<�e_�֗Y�p������^2�`�&�.dH5U����;���s%K��.� M(�'�jp"�ii�	�������B%��d����}\o�,v|���ɐ���ɸb�TI�)d$��!��St�z��}��>V7VP�Kͬ�-l�6��'T����h��K"`�8��Ŏ2Yt�\*5��(SO)GA��=p��wk6}O�KXp�����][wn����DGk3G�����lvn�ٽ�f��[���{�@
DF�D q1��/`���+Bs����߯�Yc��I`,�v!��,H�b���'���&�G���f<����Eh$0x�]�4]3OӼϩ�����B8�\;Eހ5���%][�z�SU]��b�px����yX��)���'��e@���|)2��/�pT ����K"Ԃ�����[c�kZ��w=��2�2��~���3>2)"81�'��y���w�<CBCSvl?��X���z�����)Y-#]4�ox�0�S�&��NIK[�0
Ad�Bty?FK�2��r�d��X9�B,B��7�(,B�	�=�t���$
Gi�y�Nc �э� �s]��!�~X&ƪy�|�e����j�y���*8>6����o��������w��Q���-�a�ƌA�$iFi4�����tydza�%��,��+���RY�p7�uy�9�-�[YKҀP�8��:��~�.C 
g"J��fl<��33�Cr6�,�oB�«�E�w(��F�GV��T�!���]|~7(����3��#x����>�|R~"¼�
4�
� ��2����/B��EH�W��EIp��9l�!�]N�s��k������{��6�W�Ǥ��b�B5a?��q�^dCd���X~��*:{qP�#��v���^�b=Vl�L"+�'G�X�$H���.T/�q!p�i��@JXb	["�I�<�X A�r�*�J��Ն����r�1�������]J�,�y/	O��"�����`�8�BJ�b�V�"T��Z8�t��W�}�~�����w��^�����Ύ�]�7>����vo.�DD,��n��=��m7�Dt ����?g�|�.Bkk��B+�M@����W�D�8(X�e��4�g�g9�)��=#,?� ����B=�I ]>�U�*,B�,"B����*��CU��42G!��OC��"�*h@	�I�y���
h�ɆY�iLD�b�R$Q��"4�B���p�����tq7�VXY���TY��q�j"��߁m��--jn��C��z�	gN_A�q�����>�e���PJ~qS}9~�3��X_����E��il�OjAT�oB�\>��R�C�����%]����;i����r��C�s�aW�S|2�S[�I-�롅F��N��"���5�i��U��#}z�~�������nX�p>q�zIS�wh؛�AM���*9
>6%,>5���??�U$j`sI���l�H9��T]V�����ٓ�\h3����';�������><�닩'�HG�O��A�NQE0�V����Et�Up��yPH}^/�}}}.|ӝ�5t;����y6��Y%�SU����!I	,��0<|z7As]��,¿��ԏ��������"?���"$�����>��uH�ˈ|I�$a�"%V(�gp3k�����2 �'ı��\��'0����������<������=�Fu�V7wմ�u���l�a
� �9�A���˝�X2S��=4�&��p?���&�f.?}�S�W��Y4,l�V�w�q���R7KO�ϐİ��m�S#JUt��.�XRG&dKE�JLr �/���Z�RG���e�p_ �������R��<G��p�;��=K�Kf�(6��$Pi�M�H� _2�2&[!QI1���W�_ifa�i;<��|��������m��, �v�7mX�q���6�n�j���~�ik������ll6�Z�!��|ȷ�o[r�;�':��Z[��:���YZ؛o�߸�qI��D���j���؊i��*��Yw|8%����+�p�*����+׳ct�U9GV�+�y��$�X(���"�s@ ���;��'.T�>xe�l������@�|cYD�	�\�@ 	��K��ƞ#O��s2S�D��H�D(4<�iVL�^�@�9�_K咶���.Y.�,dR`�Z<�@��z��b��_>PZ��֌��Al�t���4��mzNfJJJ���/�-���n?}kH`d�C��x�
��+dFH:�^������휓b�8 D���|��0<�
�q$%<h��[;AV�ad�n�*	�*�:��x�yze�`X^�?�$��"c&����n;�����������|u������}�VT�W]���?Bcp�1�v�-�{p��ma����xo,��V�Y5��r�eN0���0��M�M����S��{h�?�Wvn��)cq���KJ
�jJ�/^�+���~�A�e����a'n��|�Y&��������{^5�����C�O��G��n_.��rg��W�#����� B
gM.���|��U���
D�]\���Pd�O�ˇ% ,Y��"��@ԃE�d��"|���Hq1��A�hCDB�@_o�f3HUe5e�d�0�[j ;2�?8<�! ���R<�?Lf HL<[D�)��\p�U\�U�'u,�;�|��~_��w�'ϾHN��dC��D���nDUT��nay�]�D"!<�q�I�4��`�*����%�PzĂT�(U�t�	<��P%E�"� ���\�tS��釡4��b���p��*����{�N��.���j�՛�6n4"�"���rt� 
.l��Bz��X����o
.��?� `8�B�x��/�Q xF���e"�������9��n�0.t\��j�Ŗ�������4{VMw�T]d)�=*VA�1�sHB�@=�Qx�Շ�VQ<߅��w���#�1��|��A�m���<���'�Tu��R��4{�|Pژ^�p��j����~� j���<��I
���
�+"�%��"\t!�O��C����i�O�ͽ�����p��
.^�L*j���Q;:.����joLNx������e�!�~�$�¬Ը� �G�ݼ����]�>�ck��
\Ȧ�{qu�)db�v����u\��k"\�L !�/�8�͑��|�#1?�}�7�ګ�D�.<O�n�pƠ�!�=?�~/:�û�
�{�Գ������G.����4���Mqɛ�2�R�d��\#w�Y�@��w&���QgMJ���٤�L~w���6�~ڳ�������v�� ]M)i%�t�j�AО{���8/S����1']�� �T@B�|��~�_��v�JD �>�ܩyV+<�г�N*�v��Y�L��$���7�ˇi�����"�,��eY!0iK�o�
p�[����(��|*�e..5��"�)�|ŧ"T�����|x��ak�Lf�E�-͍-�"�BDw�6��復,�ok��i��j����b���"S "2�(*���Fq���,�{���ȍ;�i�x9� =I�����ȝkCE�	g���:Fx3�#��JXah�3�3]
�/�g!���[�����ɇ�Øf�QQ�
�LŐ��JC�e�u �c�ROS���o��@��P$z��8`ɈL��.��5����9���T�p��?�Ɲl獶�Xh_�6�|�p�U�_�i����&Kx�џ������l7�Yo��A2"���WD���q��&x���5?!P#�Bd*5�3.w�r:�o���bc�`���b�f µ�[��)�PlS��G~��rn�f֌�g`��QE���=���:�[@2A4
�'Q��R)����H�l��-я�@�U�	iy��%M�}*�8˔����uZ�x_;&2*;��9�mmQ�7���X|$B؂O���!��R)̧"W-�sI˔%�2���� ,,�I��`��L*�><�	�/,���J��D�s4z��Gk����R���}_�{p��a�/���_B��!qU푥M��}�2K0�	��{�b���Q��_!F�4� S;�1L�r�+��?I����}�7�� ��A����w{��P�>����EBF�F[��g�]ws��q�e뾽�o��'�'e�f粄bO�X~dPpr�_{cbr�%�(_�Ο�*�],$cg>Oz�I��M��,Ǡ�g��g�����ٗB�G�PR��g���l@�.$@����F���Z%P1e��=��ZX9X^?P4<]�m
�����;�.w��"�P?�;��7�qZ��M��˲�\��XLfa��DS��=�$�c���"���6��"̪i��C�DCL� �:@&�)ʿ�v��mׂ���G��߹m��o�?�aշ_�=~82$ %.�đ×ϝ��v���3/���{ <�)a+�y�T���/6�y�t�ߛ���M��p�U.nlh�#ͮ>x(�|�G���>QM�Nt�yVx=c�{�뒡>�$Y:ɐ�D�W��� ���z
�5TG��h�q�~�::E�M���$���� (���"H�$�8Y:�8�B:F�,�H2�� �CKƇ%�y=��^Vz/;����ŋ��ƴq�H	��==82K"��?�5s{����z�uVv�V�����henk���b# �#�ݹu����v�%�-8 �";��r�ąV ��D�`�����L�M[V��Zg���WD���zr���X��CIn���ˬ�wC��Y���nD�ӹ�ܿ_����"&�$	Š����A���5���5�c��>��5��nc��+���A,�>��������������Ԋ��l>O"���-�w���B�iD�B'��*�����㳸��)
�Lb���ޠ�/�x�qbh�N��5r�6�n��ֈ&瀜pL	<�BB���3�B�X�H)�oFSC��Ǧg�u�c����S3����aN#m�K�*�J�dP M�#�4Gn�7�����ٍ
piR��YN�H�(*1���[�O]�z��/��n��ٷ�Wo��]m�i�!O_���a1�
�����"Wfgg�e�yUM�받,V%�\�!��j9�>9����&<21 �����耇��������)C#F6�x�vrY/U��3��L@D�4�4��D�@(9�QC�/{�U���Þ�w�ܶm��9��$AsN�EEŬ�ń	��� �s�PE�s9���]U6���9}����q�s<�z�(
,����\3�P���'���dH�Ǖ܎|�����3j��o����+v^R�͓Uַ����}3���&z�>���|�*]d�5��	��]dr��I����=����A#��t��������Y���!�[�<�a=��_��'����%xR\�Lg��!6�:�|�{'GW7��훡v6X0�P{ުeKl�Z��Xpx��ٳ�����������}Ö�'�÷�'�I��nqAE��R<���p>5���zDbM���#爄WR��k�u��{��d���
ql	{��:~����.f	�By/�#�)��ׇ�~�K���#���g�R��;z&���]�.9xn�����^T�Tv�G�Ch��;+��
�~x����PB(���aYx+�@K�D２��brg�dzu@d�Ǿk���5������mǏW׷��Ɣ�	�d�mݖ/t�@�fjB��0�B�@CscHr��j`8kHu�p��,h��vj��4j�R!��Dm-M����NLtA��p����5������֦v�	�:���[�"�M��V��)G'P�r2�[X*{������lnk]Z{!5�i�ʃ�J���J����n�1����7���V&^��y�fizrMfbճ˕'��OԤ��O;Y�v�>�\Mڥ�܇%�Ks��ٛׯ�x>�ĩ3��n�E���'�aCf0�F{lA/v��t��V�`5���c���Y�%��xx+�W��}�lMeUeyE7WUQ�������yBO��bU*a��C\�f��T
�Ne�Y.�#�e��\$�5�C�X:����~�d�/T�/�`��0jD(�j��2[����U]���; ��'17mÉ�lQ|Ƌ�{���k2��,o�f�����.���̙��|��î�^�n޺{����"W�%aa{�D�MNi�$�Ȍ.Gfh�������E_:r�Tx���:~�t�;�wG�����?����oj��u6�HMLZ���(�^��� ~YO��"���?R�%����F����jlcv��;�8�D�h�+�������p�`h������Zە5-c���L�gM�y���@� �?U�auS�G�`�c"�S.��S���çV�8�qGȖ���>�o�~YߔSY�H�6����AK������|����֏_��'ӈpY�b�����2���n�w_��G�����3|�Nh��>p�������6�I���}�w��Z������l;�7�Y�����;\v�zNG�<W³�q#��V�.=�4�xrF���7���bH��h��`A�K��9\�L$�F��r�#�_Y����w0&*�8���q!:����"���fF�������>x##�����cOl�������3���U����lS���]�neE�΄���NA���E�ֵ��FT�q�h�e���t���N�;0W�!�P-B[c}���k�sl�P��Z[��`���M�����f�V�VV�A�&����z:��u�Aw��^���lG�`�mtU��vf�52�{Њ�%z��x�]"T��K����/[���SǶ�(L�O�r*��媴;����O�֤�K? 4�l�"�R�p/.�9�����'	[V-�z��ŋ�]�(�)�=}��!B5�����/�Y/
���=|p�n��g�>t���賧���߻'�a©'+**�D&B!�+�E�,�`�et�J�X��x")_��UbI���oHD����q"p�o�%"i P/;����8(��lU/��\(�|-���4Fy{Q(����E���XZPR����b�=ؐ%�)ꛀ������AK�ZXY>v�y~>�cs


*�jZ��t�	L.�U��J���YbA7��A�UTW467PT�,	!�dR�DD�	,:��$�8В�e�>��^2�O1��,Eĉ+;^xǡ�DN��w3I�^OE�� p9
"W��Γu�e�B8�`]Q�::�^�a���I������>HMv�H�;E��1�=�Ix�w=�����G.^I|�S���`qJ�Zk::l]]|��9:|��WӦM�����/�աA
���/��u�G�1�oӦ�,��r��MX������[5M���E�$=˫n'W�����95D��uv�C�"�g�k�(���^2Qr�dz�Dj�@�(*��C{�.���'@�4�;�$C�IT�T�n�<���N%iÕ'���A��|!�~�H��y]yV��l|w?bM�Bre�0��	7Ǥ�P��M[�u5��gM-Y����ʝ��Sg��)yRP~��Z��S"t^��=}=sK3��E�.�a��S"����$bӌ���5htheiX�Naaf��ΔfFz��p����HO[��D���'6�����N����p#(�d��f�SYߡ���7r�Q�$:Z���՗#{}�I��W-�[��}V"��9Me/��XE�zq-rӭc[3�ʻ{�*�J��g���Ǫӏ5���>���������JΕbI��C��ĝ�w��ވ�=���a�z�̔��+Bi�@UCs���e�)�˂###�=M�z���C!�~/���&�D�������
 �H���B1]$�#K(��w���R(M$�Kށ-"#����O�^�!#jD��&Q`s���%��1XGh/E�OSŲJ>��գ�g)/�2�_��VI�{�G�}�y�/��r��f=~��ENvf���������~��277��������?|ғ���k#��d�q�2W���y"�XI����&��@Ɠ�T&2	��d3hl:��$�t���w���%Rp���II�S���zY�~���S1y
W�Ԭ>����B6�|�v�o��<
�G�	p|Q�@�)N�{F߼���|�*��D�u���3"Ը��΃?��7����ᳬ돒�&<���t'55��004$|Ϯ�kWii���_�}��g ����Xg~H�O������֬�HM�06޶eӉcXY�n]||����@&V�߽��̹��7�=�"PyY5xvO'g��ܻ9�~����'�����t����wjo��Uq&��z�޳�n���đ�&7����5�MC.��X��I��K�Yv6�u�-�ȇ�G��	�u}�ً.?+M�褌 %<!w�^����O�_��6,B�N���v���0��̕�O���ԩjNE�9��ԩ�c�A��ҡ>�W<�vߧ�V�D�~8�t�b����7A�33�ذ3�)������f��Fz`>C�5�P�5
����զ���D��@����uk�q�l�1�ն�;�v���+�{�z��[���y_@�M��WrɒjV���[��d�R�?"�qkK�c"�+��9������)�w��>\����NM꩚�5i��Ҏ֧iL�lM��L��rgK����˛���=������������DpB�Bi�ɗ ��5���E�PTQu9���E�а��>�||���]�7����L��y~�f�)�H0
D��@{�	��xTxB����^G��n
�z��t�+��K%r�\�iD�QOp���I�a?Q1FR���ÏF�73��t�r�]�f��[WzU2��H�ھm������!��
	��V����������[6�kki"�Pu���{��U������W�p=��ʗB��F ��u�yeuM��].��b�Db���1y؎Kt6G��&6�W
����DXD�rx�_O��^���a�^�\��q����OK�r���<fe�D8<�A�ʿ*x2q���և)�[��.2��Z�2�����q��7B�ڭ;6��Ո��gtT��'U)�/]��u��eK��mm,���:w�`>3C7�%�=�Z����Mk�L;�U��F��[�u�梢"&�#���G�i���<x�{gxDDDuMS��WdN/[�J��n!��^�n<��z�Ŧ���љ�V���#�WՉЖ�Iɥ��YU;O_����T��Q������(��o��X�+�޻��'?��g4�����""��Fٛ;��N^c�F�ѽ�Scs�@�M*d��`��uB5�hb�B�iŷ�����U8}aՖ�����r>>�Hܝ�sW��;zD��I�����B�G�����2	$��ﷁ���@Df��@`���0��Y�������o�&�j�-a{-��HOW{��-3C�^���48��Ye�+�b�g���������0_d``me���)��O8��������ʖ+O�o�(x�Fx��y&�������R_����a�0"
�!���6_TQR�v7� ����Y�?:�9�ơ��8~ebC����c-�Gےw&G�"����w�ُ#q#rήK;�%����Wb�ܹs�`��6vT�����?��ՈP$SV�6$$&���:|�о�����'%޿{aݚ��/UV�ܾs�����<!�'��\����7P�k�L�W/# ��{;�O�R��@����?L����Cd�(M8L��s8*��^#![(æ���]ʷ�������,�rZ�������f�l�u��{w�w�6��[+�rϝ��t���t�r�q^���������z�ڥ�����:��;��t������������+���

GDc�ilC]l�l�b�י�������\��$���T������9l���𠱢A���z�B��Q�����N��p��iE��=�oߠ�o?�#�P~+��Dq����a7�T5��A("2jǞ��6l�)(R������$rى�'��<f�������5aи�ךme��jo�pۆ���nX�����j��
�����?��=���{w���UTaCI$8��y0"��ղ�G�/p9Y4���v�E�4���=&;�@y]�#��?�TS�y��ЍW8Eji���F�X�u�U��R��i�	T�C.�n�.�<���Qc?¿F��o/�~���ZT�N���,�E^Xu,v����2\� ���Q!|Ӡ@��$�o9�W'F�T+�,e��@���5T�ݓWE�G2h~�G��7.+�~��3O�J_W���f`inhmelkcfgk��������f�X��w��/02��v\2�62��0�Ӏ��HOg�\]�� BP 5��߷�xonc���, SskSs[S����6V=�9���ɇM2PT�~�Aڅk�e<i���?L͸� �i^AAmU�+Fdao7W!���ť���_��ۼ�9�����{�o�h˼�.NhO<�{t�� ��~�}�G{hw��"�gg�|x�Ź��mڶ��±��G�R�Ӕ}�l�O�k��ӈ�}��S�/B�����;9=�杻'Ξ���3��t��023�	X���z��Q`˶����D*(�ϓ�r>W	x*_�b�S���/D(��RD=8���?F�h�K�	JD�!�x���҄l�T"���zƨ�o����U�'�E�:/��r��7�b/}��G���������v��s�Y����%��54�-,�=,�g���W/ۿ{˾��7�ټe���w]\��]������O�C�ì�-:���B�Ǡs@��?
�G�
�l>�% 1Ed�[�����{��h�RX�df��$1%D��e��l��M�"�!K�5�)�o[�+�ᒍ��z�
L�co_Ob�~��{�����A���!�f�5�Y��D�^��/�u�/^��v=&66R=�*���/>����|�ء���ٚ�!�_�,b���G��?u$����W�X��`kn�������[aHp����6mڿTT���������A��S��t3��#����%��b鑛zK��슽^�|�W5��51)g�5���l:Y@���P-\y2\�����maqE7��h׃6��sO��Pr���G��d���{��w�*8�F�^8�(o����'�Zo�H�0�rB�#�,�9*��
�T�}����o���'g���7���A�}B���G�^K&|�������V�#�ɂ�.RO�_dc^��?�v�&�!�c#-Cc5F��]j��������� ׌��������R��v�>��b8���~��UU7>z��҅s7�br_�f$߽{�έ��W9�uuL�R6��*��U�Pu�,�xp�ދ��5Aީ7Ͽ�)�ѕ��[�ĤHڃp�����`������i�O�>�zr><;�T��e�Oy���C��t`|R�7���\�- ��v�POBx�!O$牤��#��t��"�N,_���25� >%����Qֳ�₨����U�B��\�@>�G���zy�^x)~��)��aw�0D�!�l����;���� �ckU��P�[{�ߋ�H�c��M$�r,�g��QS
��n������?`�����%�ޱ~��eV��:m��� /�%��`��A+��V.�^�xu���~kW,ٳs������m�Y�~���Uak׭���t��zUXڅ#�),&W������R�Y
5�n�!���z3KBdɉ��G�R��d��=�g��X�8����w�1�,Q$b�X�FN+�B@(�� �fn.��Pf��~8��*L��M#c���5�Ňy��o�}�7��ۻ���)b��6u�2�?�+,���������������S__w��=ܜ\�֭�t�t��;6��^�!B+\"�y������!�!K�=]��Y��}�֍{v�صc��=;�;���p�ʕ;w��7��6�}��t)_�5p�֜HiS%v�\ğ��D���ʽ�=��gz�I�0���J}���t�\�v:����M�_w�1�F�
�(�H����m���Kz١ꔡ�dg����Q�l�nI~ �P�l�k�s�hoQ���ž�sz%C�{��}��j�������]�)�������^��y=
9�������Y�-����I�fؘ즜��f
dACm��B͸�-�� K}�F�����s��"�PϬ�Ƃpb����P�B�_�0��N�����������D(+d�2�`uUc}mm����m=r`ۡ=��mX~��ć���kA? B�t����&(�ޗ���>}�힤����>(N���t��х���vk�8���(�����uIgS����;{dߩc�O�9�w?�P54B��D��  ��\�߉P$S*�Ų^�rRNE+��.�m���9�#2��5���������v+'�)l�������9n�F�|Q�څ�$B�&B�[9�蛼�W��
7��N��r�NX��#7��Q$�~�Ȑ�������M��7D?�E�ChET�<[/��???hD/v_�ac�3�7z���7��1�����]�qM��uK����do����Ӛ���֭Z�l������O�˒n�Ddp�b��Tl���v�H#w�����;�����+��؊��l�z�3e;C��&	ǈ�qo��dw�;���<e;O�!��K�RU���K��%���:%�@�hD�N:�&:���Q�����A<k�Jb�UR+��'�&��?��C���M"NQ[ߘ��������"db���vt�'�{{�����z�{��cޜٗc��ܶyyHPH�߂��������������{���Ƶ˗�{�]ln���������Ӧ͚�-�v���g|�eh���}�w�oݷg7ԛ���u�d��bQ��N:��J���K)�{ER��+7���G|�fy�xFA/Y�?2i��(�g��}w\��}�DJu�5�F��(K�n���xJ�H�>�EKi�]"�W�}P�N*���Ϋ�7	[���aT�T4	O>���zhe�����R%�#�fqK����X�>�ȵ����B��:xI%�{.�O.iMȭ�b�s;N_$P�|�H*��ݲK���o�!D7��w*,���1�A!(��������ZY�ٙ�/2�#���:�����
�t��g����)P5�pJ��;�� 555655}�BS+3+c3}#+{��G�K���J��)�^U]��;u:�⥘��Kׯ_�u����%U�A D� ]:FV���Z�}���֥^?�q�$�,.��Ή�w>��V$/vWAܾ��;^Do�<�����Gwܱy���GO�����D�e��D��'�% O"r$�)j:B��R�T�#��)_�^���6X�˧��Ȱ{�/�"�$����Ȫ׬^D��l� ����<a�څX�(W�����a�r����ﴌ!�g��ɏ.��U������l��u|Q�D��D��?�TJ�@]}h��s--
���Z��gkh��BS]3��f~g��WG?�@/�)B=V,]�~e��5KC��,�5��˷?O��P_���uyh������^v!��"�\!���7�R�3;=�7Jo���E����H�!l���ĕ{�Ց�0<�q'
���͕{/�9x�c}����nn@ĩ�z��O-��R�0����q�n��+��<���\R��;+��;x�2p�S�e�>l>g��3�M��HJ���FǱ�o&�N�:����A���/��ں���-8�z*���$6,Hf1DJ�X!��͂!�A��󠦃J,�zy���Eg���_�MsqX�|Y�_wH����Pg��"�2х��ׄ�غ���]�����H�"�����=��&Rw-���©�#��	v�.-X|�~���w��]v�r�v�	�-�#���^!.��R��#t��n��SOB�_x�w����{���X�����xk���;�E"p9#�U4���&�R�`���8��2����7���9ǭG�d�K��g�*;+	l[���q�hcsC���Ey�@^~���{�	�LO(��4�"��7>��k��P��(����~�������5�P=R!��D��V��FZz�s��31�n�/BC#}���M���⠚���'��;H�I�Q���a*K!UNT�R�;���+�e�^}Zz�y՝��Eթ�5e-�,I?��Az!��;�b��cr�.�_��������j?����߰}u��+#w�?�m���k/	O<���퇷�ܲjY@@�O`Ȯç��j�]�-�*�2%��޹P,aK�|�s�%B�_T �b.T�K��t��\;��2�-�a�%uɗ����RbDBN�x�I6I�GT�8�?��s��<�?�C=5���)"�fGH���l��#*Ƣ��x�iYE\=Y�)�D�oP�Z�bW6��@j����y�m�0"�����g���/�]��g�R�-���ښ͟	qpJ�^V��V�N��\m�������n����������R_o���U�����~>�ٙ�(�|���DH��
������#��\T�G�b�M.�b���N��m�v�';y���l�u��z6N���:~�H
��gϽl)W�l������%�%u*m�_|�&/��6��v9��v˭�m�J^'_RP~b���ϛ{�oPg�����"�P�}y�k���6��!�F�w"|_{�`�?�ߊ��B�in,�,�/-�y���<� �-��X����Dh��"��|����4	��^.���-��?�}�Ѵ�������ՙ����֞�[V/�_�b����z�Bd����W��vBg3����#�E���:y)-e���[9/�<}z�I���ɺnA9�t��,&�!bj��/��q)�䣗;c������Է�c�b���u�"����A6־�9u����^�Llb�n</
���,V"�$n�y[!|�R����g�RZh����q1>dGDiCK��g'�d�%�<�z��p�F���ӷ�Y������5��n:���������6L��J�7����f�%�-M�|mL���$Bk#M��f��f�(�;j:�]��85Ԉ,hnd�ɂ�K"�3~'B,��]N̶�sl�����G���������\0�}b��EL�d\>���o9ʷ�E2B����4tv�>~�quؽ뗀ukV�pc�ыaᇃ7�Yn��{��çb��v�辻�.>z�hW��}����O/m&�N���\!$?Mw(DC,Je\��'W+SaI՛�'Bl�&8���D��1��uNg���7�x�Ihڑ�r�e���e�prǽ^rG��P��-U�����F5"�\�Y��"Ը�,�٣��xݭ�8����RB�kd}����֋đ�ɭϪ�v���r%�|�E�c��c�>�kW�6��c�m=ݖ�-_�r��__�Esg|3���~��c�_�3��"�p��t�������?��ۏA��~�03�P�a�:_��gO�HN{3�K��b�����߬��1��2a���Z�	��Yř|��Y�-:�U�"Bm|�����a�Kܕ��x���+��y����n��|���:�C�w��%tY���m�����m��^Y��:W�e ��D�*T�AY��:� g��� qE%5u�#c�~�X�臮����D�TF+��F�tQ)x:���r�^Y�ڀ�.]����Ό���B(~�ŧ B�!�P_{T�����I�s~�n���04�� <����bO>�y�|���kN�8��wvu�wZ;ȭ�VaC����We�:��-
��]_q��ӣ�o���vIz��1�[D���]O�~^�T��m�8��$��;��Z r@����^���������C�b�޽��O
�G��k��87�ey�b��]=����WMt#��ls�h�f[�B��ݔ���	��?�����;���:i��%Ux��W�a����������F?S�۞^}���021�61Ԃ,"43Z �p�Dhkc:�L��!��ꛚ�/BP dMMר�)�N� XΧF���"41731�06�0���3��rp;u���CNO���k�<\|����eq�k�V�{P�)�վ���v.G�D��C�>D�E#�B� ��8��U5��,,}UX�U�~V���&���~[~2�6�Y����̌����²��͕��h����(��c,���? �! 
���+8���
�ꀨĎ)i�d���U��ћn��JǛ�JH���r�Ŷ����]zL@�cU���B��M�����~@m�!B�n�#ŸƂd��.��#������a��:k}���G�v^�>p�LIk�0ڟ^~�J�2�bsIN�O6	G[x�]'O���,�_��\hg�-H(��uڿ���5�P��/?���?��g��FG�W�;qr\�V���O^vws[����Œ���oW��})�Ў�(>��Z'B�Τ�q�%Wl<��]��o 8��1{N?<v=��;Q��G�e+Ѽ���Җž�:�d��܊���ı�+O;z`����w;G�����כ��FQHL��>�Nj�mQ�v�[u�(&�Қ����1l?�"�P�����)ʫkR27wu��.*��P���k��i����F$׵w ��n�����7:|:��bO7h�.��y/	�;��Y����d�848p�֍aKt�f���g���T��������f�`�9Zs�/�w[�:���Nk�H?�V��\��m�Z�M��%�^݌�����XS��\��n�&wh�kw��FET�7�ؚ[�������}�eS������t�D�D絳D���k���>n�w��:/\��{�nSc@{�����ox�/޻�pġ��,�ƣ����W�����BM���7c^�t�!���H���nm���%,yL�˛��	�Q:s49����XV�QPBOɧ���J$����^��F~��8��L_o�6PH��}��L����R3pTs43�1��R�54MjF�@�fi����C}-8�m�����l,��bb�kijdefΛ����/Bsl���X����J����g,�H5H�J���ܚ�/*R��_6��j�Ȯo�q����W��q1�3{<-�u�zBvu+��݇��+	I�)NzQ�tÞ��sKۊ��M��FVq���Q�̪�4vqkq��Meum����.f]��Ƕh�T<E���W W��V*Yr���\���V
bW��~
���� A=^ۮ�}��;���zQ�m�U��QUR��m���!�:�ꅓ�[�`�-�@�h�"�S�-8̒���^D��)'J���f��s�+�"�t��g�]�o-�5���L"�0b�Fiu,� �b�:.Z��PN�Γo:i����a㊭[V.[�X{�y 60���\��`���|C���� Eׅf��F�Ůvи����>�۴O>�fh0��B���Z�^��9�8n}#�ΐ�Y2l7y���22¨�H���C���/�N
�s�y3����-�څ�;���G��F'ैЃ�2��n^q��P��<|�
���;��+y��g��r� *V �m�#�u��"��ɛ�W��P�e1����wŭ=��;Nd��8ؼF�߆F�D8����.D����v��]�:q �N
���J9��"��[[kW7gww�� :�ہwn۬��98�������6(�}�� 0_p����-����3]-�\��!��YA\��D����CW/��0��^�rE����3���K��k�]m$2��c�O|�j���kqsL���88o<x���Д�����;���h�&VT4��K���XYUZ_Sv��~G[l�#sc/WW5��������sˎ���+��W��䞱��]N�Ý��9p'��� #�k��Zb�h?�֞�[}�b���-�����W��ƽ#�z�KW���k)���P�[-�?m��}SHl����D�swY�	h[5T�q���|c���p}���F�V�F����"����==m@�N�C���9��ڟ����Z��f� �SD����O�[�G���>~�����t��ʹ�O���� �'C����Q'�&U%{�߉��(�����~Wy+���w�z���#W���Iq��.Qs��KH4%�� 1d�ϑwq� ������ B�P�J9b�ƅ�PŔ�!�o��LŔ�t�$<p�F���$�+��B���،f��iI����T�u��&�8E��)�`�F��!��ߊ,Ȑ�R��aD��>y?kGLB-w$�rʉė�a��P��z�|L��d%]�����	M\�T��C���)���9�~���k�߹w�~ֶ��Z�~���w���VFN��� ���-�t�rZ�����"���h������������|k+C'gL�n�~)���8NM�ƐSY
a7�/x垛	��Y�+w��ndw��+�,0���ȫ�jhx�$9")@�(�����Ѹ�����Y�Oܮ� ����V���Q��x\�P��=��b�kR<l���=����8l����[�^��z���`��U�����Ð8�!f�"�P~/�$��55I���9��;މ���"���`�6"13/����/�$�%[X����w����������A�v����6�_�2l�5Q���=�<ׯY�c��5+֭Yr�dD��sH��� ���#���]dk
qpUX��"�7sf�����.\8�{w�����
�#QJ���\����p�ڍge�W���]���0b
�oT04A��2�J�'4�6?�|r�ޭ�7b/G���t��pg��:��⮫o�n㎊�N*O�ArTc�	�D���*�D0���/�����mEF�L�3z+Z��a�]����iv����{��@|R��5�^�[q"��_�3�P��o8����N� B03���UZ[a��شzuL�u4��i�i߃5�������4�u@=}����lJ���Z��掎{����}����@�z�ѹ�����9p�Į�G�_�~�ĥ����Ye�D71��Z����-�
�����>kv�Vw���Rz.�e#m��3��Y�D� ��Of��Y�Tv?��K�ah���L>S[P	0�XW�fU�)b
T�yO���mR9��$`�~�t�.#�&�=�(A�ҽ1i���[�[wF�>o�;w�~A���Ai�M8L2��,a/[ԧ����n�~�dP#Bf?�?��yn8`�u��3��BZq &�qQ9I�*��v���(���Ȋ���n����@8n�փ'V���߸u�ְ�!v���vFfZZ�?ϟ����lȂ���SY�c�������%$BO'k��,¹���:�/NJ�n�`WՑI49��$�������i׉���>�nf�5sI*t�FzlZQ�h�C0Z�«A�y^0�Q�v���_I�a��/=�(���zPg�V^�݂�Rj���O+9#��Pԣ����M*���=x?/�ȍ�S�J� ��)�x���2$�����t`db��&�w������T�?"B�M��)\�F� qT�����8.($����߿�������g@�
��^�,�`/7���m-]�l ��]�<��x���ދ/����������Z�׬]�4hu��m���q�5y��U�ń�v�/`2�D�Fk��j��ʖ�6rZU+}��b>���jꮦ�:%P�42��FqSgIM�L����u�^����������~<7'7g8x�]��a�^�j���j%�v�p��*��s��Q-^D�*ǰ1��>$P!�	��ɭ�J�u�Q+���*h��D�>��D��t�v͡�j;�/B�� ��@�n�8��Z���`A ��5��47�Q#B��F�4YP�MtA�pnge�ߊP�D���l��������(�P���	�5$J�턃1�k�D�_��خ����Y�[O|V���V�n�z�%����~vmw���c�KH�O���C#��9�Λ�qF�A!��O�:�v�DH�kD�0ꭔ��A�4�C�`�TLqC<�QCl��h���K��U�׋��}�$U} /���S��$�$�����8��O��}L� =��J�����wϯ���Z�=-��R<^�2������6�����I9�Byͤ&���?\�)*h�w����"BEu������<dɪ%6n�?��z�Ό�g��w��_����3���o?~��3`����q������ |���Q����B+���b��vVe��� 3{@�$����#S2���)��K�y�6� N2�Eeݼ��W��
�(�d����ty9�K���c��	xX5Y���u�F;�#�g �&Voo��?H@��,l��zސ� Y��|�-·��*@�����odb��?�?��yh,"�Cb��t�B�I*�/���Rq$��]�O?��?>��o��XY.��\�<t����_g,��+����Ҡ%�����h������؝������������zyHкU�ׯ^�m��k�.�ٶ�IZjW[�D���P�jK�DL:�)�e��9=(Bw�I��'�O=\u[;d�����l�˪��ѤE�����<;�F!u67ܸ�&,�P[����������������9{���#g[�����vj'[�C�(�7*oeV����X�Ԉ�#y?������I=��)c^�^�S\�S�jk�מ�6v�9_��-�X1M�n���f�fN�FE�D��
 ���4΃#��5w5v�GS� ��# ՞�+| '�&M�5��o��5�����Dhbi��Ome�mb:���hѢ�G�pgp�6bc�ȼ�zf�i-�e��3 ��5V�m=yH�Ew� ���h��Ok�����G�SU��Mt��"R�7�g���$:�p�Ӌc���
��W�͑A��d2�sR=��_�����dA��b��P��4��8�A&��*�7����y�4n�;@�`� �� ��X��иJ:_E���|��`[.`��Q/M�O�vq�AA�G�w�����d/�m�gq�d� $�F�R`�,� K z�%p߶����i?[�i������m?��c�_>�6����A�Z�|����~��_}<S-Ë�9�ǯfO�z�����~�/?@���>�tگ�����t�p���𲰥����(�!��K�6�V��la�@�"��T��E~�b��+)�j�xa�������,TD���W�xrh��	@c�p�͓a+ˈT�����n�� T�7%�weR��J�AYU���~(���!���Q���x��Li�uW��uv�56L��O?���/~��'+3Ow� ?�9�~��_�}����/ŮA�b�6�L��3[dg��(lYXp��5{v��>ztْ��qW��]�"W-��i��3�;�n������������\v�q��茢&�0���b��U4u55�הW�x�<-�Ю��VV����6v�n�N��^�VQg.�M �x@5�:XJB�hG�3\MϬ�f��n�p=Y����ۏ^���_u^K*�������$7��ד��|���3`���1Y[O&�֑xB�H�O�ڮ������"�
��R��K 6}�XL�|'fF:pΧ���J\�(P�Y��y�D_{|���v�����������}j���7���v�H�*�@-<ٹ���GbD{�<����3{..;tm����̪*Fo�Ք�I�N?���p1���3�A��?��6s�#.$ƥ��>�Vf7g����q��n�$I8��2��,��`�To�*����7���'A�c�G����^�D�������D��&�1���r�pL�2:���q|���Vl���Q�[�[NZ�-qS�2pN�J�S��!\���WQy�4&�4�y�lj`�Ej$�4P��T��b�E��>|ͦS;��n6�:���i�~��_f}{�dD�˧����_0�?��D��`���������,׭>rh��Qa+�ݼ����tՔqd�;r���*�i��N��] l;��N���˯�0
�q�
یW�Kc�����u�^^�PB���I�
�8�f%X�<F(��������b2S �ق�"�P�]�?(B5!�H�|�~��O�=zT[[��O?��O����3~�05qsq�����3[[#L���A���|��?|�����\\B�B֯]�u��훷 �&�S/_�iij��PJjK�E��M'�i�5W2�����/^�a�g�fdo��QX�R`sz&_1V�����^W"�}��v7.n�bow;K['{wG{O����r����g��]��r�Fb-QTAQ��N�a�{����H(g�����y�a�b4��q��f�䕇��{��Ui	i��]K{~3�y<��yz��н׊*۱��ô�񅛣>2t�k`���ҒFE�H�A�@0dA8�B����F~�Ǝ�)�x�f�)$B�@gv��ݢnFS�Ro��6�������p��F��EF5R8��7����O�:o;l���ʽ���o9������V+&�Qx��&
�xe]9��6��abݯ�yxɛN�h~-�fJ�uC���w
&��o�9b+&ي�Z����,���[XGh$
��(���&�I��Q�l�%���zը����PK�`�d B�XJɈB)Q ��Zs���bsU`A!K!a)�L `ʹl9dw����dp1��8ز�PMS8"*WL��0��v!�-h�����&i p�B���Lj#v� ����G��h�Ih��q� ���5�ٲ�k����"cs]�t6vF�/R�N��7CĎ��Ů;7�X�����n�����a��"����v��qۆ�uՅ��D����9��9q4 dť����:jIBf*�,)�ylAm�a�t
�"^���%�q�]^$ŋ�x�/���ݸUﲫ��&1&���rY8`'l.���sx N 6_ ��B�H����<�O�������@���D����25d(���!D(�)&^��~���)B��/~��G#=�Ev�۶��5:l7�o��L�z.�r �"��@w�/?}mme�{�W7GggǕ+��Z�jǎ�6mZ�|��?GDD\�~��ۉ���$�e�r;��ɣwd�߉ؽ�Jn��604����y�������b+k�}�]*Kсc�*���z�$2p�m7/�=��ܸr�������F�����յ�+G"��tP��7��i;.��G{�eD�[�lyN7}��$�'�=��$�WJj߾)��U>x�r*����Y^ebdf�?sw���U�B�X�P���k#��,�[
{�TԸ�q�Fc�<;+���gh\���8%NС&¹F� <���"s{;l<�fxh��9Ydg����B#B)�@�z��5"�+!䷑R*�5p!��TZn���ۅm��mg��!:��$]�1� 6E���
'/ia�Vv�7���(��[����q{��U�}���%G]I��z�vfA	�s/��s���W�_���O]'�'(�q�|���ˇ�A��`+�Ԩu��a(Tt��&ʉ"A(�BE���o7�z���
K�,��lY�F���ݖCbl{ �,�gDH��4h(�N��5ɒ~�T#B%E.���&큼˕�6������W������,2��5q����w}��,`Y����WNVFK��A�Sz:O���t`϶�'��==�GI�읭}�C�]�~������I��,1�-��F`>#�x.�ct�X�<N�#�����JpaG���`�<�f�"
�Jc3�l���7T�P#B�fL�s>�#�w9�D\�����pj
��L�����?�]�D�U�O��X��[�j�.$P��dF7DHK�o^�}{#��<�/_��_~��7_}�Xp��3u���-�n�Y�z% 'P�Ν=j[/Ogow;��怵��������ѨC^^�N�[�m]�zզ��W�Y�����{��}w��MIO��(�wECcU[{�������-��H �s�̟�-[����nnNa_�DK�����J���z=��:�8ZAN�G]]�[kk��.�������Y��|���'�U��{Z��p.%�EY)F���fA9�B(��_}�:!:B�+[<Q����llo()/�y+v�2��;6^����{3�t����z>�)�I�%}�kO�v��-���2M����)�9M����a����,�93��7�7�}�D��/N=R�`�O.�o���"C}m���/�vsq��p"417S��1�7��5��ol6G����q�����4� ��Xy�B��gO
s.߿{�����ed=�.����(W����'����a&o�'�L�O"hj��x���A�+��H'�Yî�N�=q��ç���IE5]�����7��ݻ�jR̓�]�iC����7�p�� b�M2{��<G�J����@�q|N(�&P#�dY���*��*�D��Z��:2��&��:82��5$�q��>l_u9�/�D���r�� ����"�:��|)�����Tm�w�#b[a�C��)�t�Q?@�R%��i2)C*eJ�⾑��{}C�.^�����akcM��W��y9��ͱЛ��TR ���2_�P?�?�P��@��K|<��6�	��q<s��}["��Z�haam���x=�vE]]E]C���5��R9:������Rd�F�0����bs���W�/�@�B��Z~fAL�
�HB	hB5|�l%X6_�8��
E`D���}��|�*aZ�����QH4�C"Q����I�uuu�Ν;}�tm�y`AH�v6�
ׯ]}<����'�L�u̷_h��������#��E��m�M��w��֖n��N�ظmK���ށA]\L��u���.]�n��/�ӟ?�mm��XT>�v�݇�|�`�����t������iY�"c.�I��d1@&a�Vw��-�l����܈O\�j���ӌ9�s���������S��喵��og���Y����"�F����mP;?m&���M�FP�˺�Wt!�D�O�j$�?�nwԞ� S�Jɽ�$:�AgG��J�۫`�z6E~d�������<�&?KS��l-�YiF��9/�9�[�̃D8e�)�S"�l���?<�L�P�]��5�!\�����9�P���31�1��21�zq��9�x�훀CH3�^<�͸���{c/��q��;w�3j:y�~��@��eA��UASqq]�����7� ,�%)O�Ҟ>9}�ҥ��=w���V�i;��+g�F!5V�ynf츚RDU�&���c����%�ݪ7�ID@8�8�O�l���d�L����O>��q�r������و�W��\�z����6>l<|:��}�on?�&�l���/[���	�[D��G��`�N�B�SW0
��s��H�5�^�,�,���w#k0�@���b�Dȑ�:��{w����-��Xuxo���_��ӛ5�����D�c�� �_�u~16��$��z����������׫�k�����Y
����+�eB�ۏ��aw���!�'���4�Up6Y�K���w�B�Ƈڅ"�,R��`@��� �^_��!�i����ە��?����/���:a[�����f��w�����%!@"өt6��RQ^������<�i��� +�ys�Z�A=k	������+(�Ϯ��@�A�u_L�~^��/C%nٴnӦ޾^�v��.N�Ϝ�y`���K��\}|l�,-Z�qS��]g.Ƥ>�ʭ����l%Be$��⚄�z��H����,���g��=L�K<��păBٰH>�;����8����˷��bn<{�8w5��5��է�>j�����v������e�
���=DU��j�U0x�zj��ug/�ͪ�yZC�Dub����x���Ѧ����G^��3Pv��w��)�l�����9:�jii�hA�3`in
��X�9j��h֋����,��V��@H��]��)H��@���Q#BC�+B^��HK�'�;zb�ƭ{�oٷa��m���?}�BS5���K߈D�ӟT��x�����������mbl����Rll���M5�S�r�;C�����E-�5��#H���	'D=��SA ����i	��ڋ���E9�Ԍ��.^��>�j���nN�h������S���
�Qb^�'ρ�/ro=ͼ��q-�	�0�0��-1�����3�����h�-�������t�3T�`A�fЇ*C�@M|��w�P �B�H�B@ 	��5��s�J��\�!C��!�ärY��sZ��3%kCO;`e���W���g�ڿz:Y�xh���L�_��l33К����|���~������������cѭ7:�*��p�.2�F�0�\v7���t�D8���-�bI1�rK1��6�EЧ
t� ��7b:$
�����F��uOuCk@��5Ƃ �a5��/Bl\�����Ty_�5u�)i �N����_!����D� ��4*��Fh�1�m�m�6o�ps7ԃZx������3(P�)�� ]0o�9���wsqrZd��`���������Ǵi�fΜ���d`kw*&fӎ�߷t�l����Wee�MT���a(zi���"Y�s:57�NƱ�W{n=�q=c�����|6)?�����`!��!� ��#�Ǜ�|��[�7��X��-t������l�Z���.^n�s'�����L*&Q���QJ���i)m���1�p���V4��eVv)P��mZ�a%�Q�Jxh��{a�n��vj�ғ��D��{�g��f!QO^��d2��!��,���_�,�"412�05L�� ̅ *u�[hm��
L��=G�4Ͱ�?�pʅ�F�x�j�Z�Ԩ��OA�451��6wvZ��`
�ᢓ�BM�(�s������|������C'5��*�'���;��_>�_P[MOzT��^��ݘ[�Q���q��
Ė��R|vYWniG~iS���gO�	�nob��'���(�g�ߵ��+/$<f�<c�fQ�pԒ��V�r5Sr��T�i�zZ��~T�%�z��#����D'��d�����X�t�B��:x>hǑ6���'���|#%�c?)z��H�/���~VP���[���C�T�%���
�����V�<1�� B�D�J �'B�US"��12�R�D���T*_"9q�,�A��^`A,.�_hom4���f~�/E��pܰ*��}��ߧ��7����k�����>�<�n<��N��v*���
r����R�ZO��M��fv_+���՗[O���-&�F�m �d�@'O���J���D��Il@��0J��]x�И5wd����!f�"�P~/��995��o���w"�S~a'��K"$R0H$6@&1)d��%§�<.���;�j��3~����9�@\�li�΂��}��7_}1s�O �p$ԹnN�~�IOW>"�>}�",�����	Y�����=���ٲmɊ�O��[p`zB+�[64�_ۈ�(ZR\�DTR��ߪ�gn��>t����]w��x����3i����r��A��*l��ߠ�`v)��\͔t����{���K	�;9eDn~+� %�G��a��5Y:F@^P�E��D���I�doE�N��)!�԰���|ս���r!����3��ΛV[�ꯎ�^~V���7�G�\IȄ����<�_����̚�����m.46ԇ �#���<@������)�0�������c��q�j����d|�|V�pqʂS"������Z���ZO��!�`�M��FS"��g��������	��.�B0�R+�ӎܧ�}�u�� ��էsbsh2	�,T�G������0���y����	r��^�w��a��E!�:�{�jw7[�e��,ί붥�k�;�~�r�Ӯ�8�ۚ�g�D]��y�d�����t��t�y]�`�E������
������o>��Gg��w_�ه��̺�WSPW� �N��'"�UiΫ�<������NB�ô�K�o�>90��#��}�=9��Pœ�i,��_�������#"#O��:}�̹�g��b��۶s٪�yE��{B(�r<�B,W1 ����2�7<������D> �b���#�c�{����J�X��RQ��H4�D�s��%�E������Dhogbc��[���sg|�?�g3���f�V�rk�����N:s�;���?|��w���ͱ��sv[�����F���Φ���nB+�I�,�đX��i����h���aQ	�}�ȭ셡{m�w:.ߛR���\)NHR�v���K.=z��V���[�BL���-�.j�oԤC��Y#�w:T�P}G��x]u(�D��>1�A���D����A$������.����3����>5�+�_WgA@�5���Қ�ƶ����%�K�u�<�=���N�^��K<�\���6=bڴ�����������~YȒ����ϰy��|��'�|�k��8 ���"��9�ea��޲{��UK�<=wFD<HM�dO�?x�������D(��.���R�=G�$e�^�����	N��]{U��7�����6�z�>�]P�Rߢ��g3r�˯f��8v����OZ�}Y��x�8�D��N��e�3��aC߲}��ژ����G�섟�9���wg��3�I��v)92�(�a���Y/�E\t�~��ٹ-��N���p��/s�V��RK���^7𞾮�x��u5����b���������F�Ѐ���W���S�%�	�])5_��D��� �F��##c�1�g���e�mn�qT=�CQ���9�;"]7�����3E��<,�� ���D.�f���7��w\��E�k)�^�Rf>Ц�ވ�.�ͤ�.�8t,b��e���$�y�v�ؿ�z��
BUP����#��PY��y!������O�F�>�e�U�ƹm2� B�rT�Yr�V��*���y�֪��}=6��r|\L���	1�ͅ�/�s_>��{�_���ٔ��|���}���r�B�T)�@Z>�N��!q��#���`�����b�������������  xպ�z���>�P�w�y$�������=�X�Æ��S�d^P\��3��~���.��jB6¶Ta"�29Ret̕E.~K���{�M��̞>积gO�N� B;SOG[�m����9(p���}����|�7������B7_w{��I�����j\w3���W��^���V�3P���A-Jt(>�IS9�u5�uV��cӉGE8�
��gݡ�¦6N/�w��-�H	1A ���O�P�n�&B1�#�gb� �������և)��$�)B.���S��t(�`�ڙ�-�7�4�Ӏ�Č��͂"�F�RH2�L%��2\H%P�[���fc�(�P����âEK���!����~��߿��3��/?���vr���r[�*l��?���3~������~Qph�����c�\}|w�?�v˶��0_�S11���nٵ#��-<���$������q ��Ԗ�|��j����������;�Q�L��'�O:mٞ֎k�Lhj��<F@h�s��˶���!rb��*gJ�k;�ħd7��Y�ژ��細��O(����=�e��Q��!����.�ڏ�Vv�{^�QҴ��ٕ���?w����O�Vm�hnh��}}=���-�?6r��o������dhm�9�h��� ��uu��0���	5��� �� �5h�L�� �AM"T�v����)��hh���&��6�1�`��݆}GD#(�U�ћE���\y���H�?u�i�����)]����n�6�HK�󮔵ļ�~Aậ��`l0b ���Cn;ypۚ`w]�Y�Ξo��_J�@�E�j5��6�e=n�2&P9�Mn��	���|��'��ii�.%*��-�Q&Qm�y���^��C���6\+�f7�=K�H<��(�I�Շ���>���p=�����o\�{���]���{�l�P(��e��Ʌ�X�����*�j���i���O�2k'7���������%�����m�Q\��F�9�6��(I|ո��尽�;c��h��ßSw���$�`�"#p)�!�p [.�1�E*�'U���[d���B��ί�L����?~�1��v��6�������u��������w_|�����Z��4"t��\��t#�v������!�V�{L��Nh�R6����JF����S��.k�9�������ˮ�'v�Pfgž�Zj^4L���E�n�I|��Y���D��Ռ!�L\�F�p��Uآ��~�o���Oh���dy_���- �.2��u��� Y���;��v!
� B���,(�\��ш4��#SpT2D��r���n_�b�<m��`�ž�A�A����}}�V�-;|蠏�DS��Ehkc�u�zȅ�ə3~���޽{��-]6Gk��}���ܶ�޻|�:�%A�>>�--���9����g������"��nwRփ�'��uT�e�'����������O�7�;���L����\Lģ���6�ި�:�,w���S�ٕ\e�|$>�rͱQw�H=ؾqj�����Q��5�]~AXy6��u;�K2AV"�[d�d[��홇�[O�8}��֨�5��{O^ħdd�蛙}?c��B��'O��]?�wM�C��!���öS�0���o�E���y�4"�?�����6�(B]�A���~�њ�r�fč��-`ki����e��BK{[+�mBM��B�D�["�Ϙ��a�p`����Ϫ����zd*BO���b�S�����I�]G�$>w�w�)Ix.�<25;��~*1G'�g�%��xm�E	7Δ�&��?�{�9Yi~��y�@�6N�����:��T�@��z.�w5�6��֞L�ëZeh������>��^}Q7�.W���Ӟ����[9ĞԜ�;�/�?�3�����
�6�,���G;�y��-[7lڴA"�աP.AȨ@}���+�|�Sx/������JС��ߐ�~����Z-r��<y�Nґ3q�j�W��e��'�e���jX>��$�����{o<� J_�x���j�QEJ�o�� BS(����"\�dIp��� o?w�_�f� 
���'s~�F�Lc��V�?{swG+/W�)�������V&�,�^���������j��ζʆ�6\;�F�`+J���m%��nY�Aݟ�+�C�u�����~)�^Ԥ@Zn[�h_v1��_�E�$��(�D�A���"�S���y뚚5"�¦�1�L5�gAEL�H�Ti']���0�-,L���o"d�) �L��B"Y
��"�G��H�����9Lr'ϐ�vR�\�Yv�ę5��\���������;(�������޺ycHp����f`���s�����ۦ�Ö-��������������e����_f�����镐��$8$0(���=|Ϯ��CW�[�,����\�<�����$5�d<�/2��O�?;��o�td�����.]H*--�P̓B�ߺ� �e�������7yD����G����Ql��f��;doPo�[4A�A���P��x���/O>�i@�J	��&@G�]<��Xo���ѷW�=�l������S�%?HI�>�++K��~�l��[�m'�)��`+�x���F�n�.$B}���@�ZS�!��`���:�4��j�65h �F��h���U_k������������������������9���-�͍̌�K���4��k�jDh`d�gl�cl�mb:S[o�<]-S��{u0E;�G���#*������:�ԡ׍������i+�iӾ�f�K�ԑ.�V�~R����PXS�k�t�Dl�	�s�_���V�<I�H�r�fb�"$6�1*�7&�/&sitF蹴#i��I�����x��'Ͻ$:���9��$�^)usLڮ���Z>�)�!SHV�c
n�Q�-��N�(��y#i�!뷬ܴe��m�vl�8y*���# W@���SSR�28<O$$
%W�uNB�2>!�eqEAem��LK{gKG+{GО����"7~�a�6NA!�O��������)��ZM�)��xX�ڃ�l���6�fev)��o<6���ᤓ8���*6XF�!�;*��y2�@�(�1�p)���R_7W#�9��4g�W�~�Rgޏ&����,��z8[{��.v^�������h5�π��d�W^d�*l��a�t�^FUkGImMcGG;��B�W�A;OgԱ�è^�*��5:���Ї^��6^||��֪@�{nl��\{��C�%|�-��H�uw���T6��7���wCf�h.׬{�n�k�TT����L��Ao_��7��� �?Y�amc�G�`�F�Y�x
�@����!M�Ɛ�0�M,L����<�^�&bY� ��$�{�=�"l7��v�8mz7W(�"�p�^W�2s��]5-]��\M�,~��G�}��A��CC֮^�}��Ñ�.��_h�)�[�*�J�ukΟ;;�K3[[k''𝻽�3�pO���蘋`��k׹�{~��7s���}�nݻ�n���*�B�K�w�2��yx�^½'Y�+k�;����>/�� ױ��#���x<���;Ҳ�|���~~��Wu5TI�ϫq����'�y��GDL�$!�B�d/{}���Fik#Tg��ЃW�<��0T��]~(6����'�����!+��>�º-+M͵v�X�%d����{��۴�C5����G<Wm�n��<�?�3�&�U����,���!X�gcft^h�����N����p�m-M5"��2�] _G@�<Ɔ�F�fV B�|���܈�W�#�[�³w�&������#�m�#�T޹���*�����y����	O�9͔���˷.\�?��]O���4W��?Ix���fj|kU\����7��q�R������e���{m�nS�\||���2�J��A�@�J�ً*x�8���(��(��\�ʤ�s�����[��{.��r p���e^�>^���\�vugDDdԱ[w��e��t._��LFb�;�w>~���$�̥���@O? ��/X�������Ţ��陥���6n}�vv��ӏj�Q��R�"�eT]}DX��Nd��,��"dHމP$�2Dg��mٺ;ʲ ��дΚ���?|���ϴf������LS��֦:v��6�`DO'k�E���������`������c��=��Z[�9x����p�Ee+������Ja�Ѕ�D�ߪ�G/�;s#u_���̊�v���QkcJx�xϥ2֛f	:�X��dZd\Ns�K4��b�(D��="���,�A��?�.2q�ꦦ��d!��%B��~�Q���!ob*����.bЄ]Ty���<�Ej'(��ή����ւ���N|Km+bP	^��XG�l,o�L�.پk�e��sn.N���h��n\��Ё��N��ށ��!޻��}����smmm���]�\gϝ{0220h��[����?����8}*9-�@&��$�0�ۆ�7M�������^Q��W�5�Hʫ����|����b����|���6r;��JJ����t=5�Ѕ{�]<}#���`���`A�� �{Гfz&�W%{�Ʃd��͂�
�2���6����׈яrj�!!�
<���Q�_�y����d"�
���>�+���Q���!��5Z�p�6�@�/�N�j��ߕ߻F�~Ou��t�C�9�Y�����^�!>��F�npW,L��������:���X}{�Z�of�kf6S[g��6�YL����6�X�n��G��DV���[5v(Z��K�p�;k���v!��;Q��`�$�l�p��<6��Do��!���(�됏w�����*��H�"��(�X�y�KF�Z9�pj��'q��Q��\~(8���"r%��j�> ��~��u"�^y��̝�+�=�-�y����Դ����޽q�̉#{�l[�f�����_�x�칄�T�Tœ�pe*q� K$��X�8"�������/�G_�vrl19z�+Wmvq]�K�w
���[Yx��!E��ؑW�6�'*��G��_y�X����M��X}]�w"$�5"�IES"��4�4(h���[�/tu��?���?~��w���������?��?����~����_�����3�]0g����p�e�?~�1�A��>���?����_�Ʀ�:/��Xs�A^M'����Omg�X�&���ՄswR�F��s�V���5���.΁���겻x�xN�j��W2jr[D�Ǳ��~���x���aJ���m�!BMרƂp�7@�L����qxtr����"�P�P�aUc#�P���_�P=6�*젊[�=-��z�@=�������to H�mty���5�A�F�h����{.&$]|x���؇�GO��gj���f�n:����$G%�쭻��_�zEزeK�gL����ޞ!�����v6֟����fޜ�Fz�H��p���ӦM���xyy�yz�՚y�H�ҥ~�a+��:��'%=��M�RxBA}S#�'�$�l����(^����Mw���[��_��c>ˣ�7�yRBb�#�0�`���o�K�)�b�����&i �q��v���[�LQt��[��n��;����=�A\��� `ot�'r[�w�[���?�
'���.��#�p�祥���M���굛��;ʟ?�W����pE)㍌�	zG�g�Z�����!�����Z�t̟ʅ����u������|�����֦v�>nNK��!&���k,����7ŦO����5~]��p�)�� K���ᵑ������>D~��oPJ3�}q!.KP>e�F�C�C�#^�n�N������>�D�&�vJ�;���1�,."�|w�^r�Ғ�����.&��3�#fǵ��g-����ڳ���j�����7�$e4����v^~����}%�Cu)���⳸��+ٹ��~�n7	�/_�K������b:����y��q1kW�667`K\��L!� ��oH��¿Q$�0:�t��G��ol��z��͌_����0c.0�'�����f�-ߐ�������RY*�t"%��{Ů���n9���J��ҋ����7hb�v����1�� B�<BL����HAe���Qmmk--��%A�>�Vsf���~��G�}�~����~��_���Ϧ}��߾���_�cڷ�����?��?�����$��bη��2m��7����[����K��h�ՍMVS�c����|l�����-f��z����o��c ��5^>FP�i�������6!
�ɂ/B���^�N��%�?���ш��~(,V�T� �@�i4���q:��z_���6��Z��ZF^�]4��PV��5ի!N�(r���Q!.�|��c�u���_0���ͭ�7ľ�����u�x��U!�Af��	js�Hq��0S����矾����m���������n�����/���_~����������"�D-]v�����+��?��8���W�
;:����d*��������PX**w��!�F ���^�F4h��bՍt�"�Vj���9I8o`x0A{d�8@O�E� I<P�N�P�����&F�؇6������u1E�Ѓⅴ��vD����;��יEEq�K�J�'�LN��,3!�����$ܾ�T_"g+����-_�6��k��c���o�g`bdn�?w��ٿji�Sk���4@fT�P-B=���@��R��t̶45 �����/�t���la����t^��0�5����Bk{[+k�wP�ZY[Y�tt���cf�i�An� E,W�E�u��W�tnˢ�ޫ����v���'���g����"&8�B�}�R@M�^>B�׈>��!�R@;����9��I!�����l�<�!�W�S+���q@bYWb)�b�Gĥ?�gA@���b�(a5���2����n����^�\�7���u������gOӟ�$<I���|;#���a>O�R��L��iH�T���΁#��+$W��!�8��L�m��L~�5������]��/Ӧ����.rKNyN"�T1�&�1�-8V}����H�3]�^�j���zQ���S�D�,8�-7*V1�2�D2%B�xX�x��cw��o�E&��G�ˌ�������/ٲq�}�׬���o�c��3��2�u�53ћgm��bo����D�u�E�b�Ko���5ׂ�����l�:w'�ɫ���jaC"�s�p��H�����	�)8��Ј�l�D��wXQ�Q�oˍbK�фt����=����P��OXQS?4�N��|(�T�WDH%P�D�@���N���=�̜p^����Ɠn����S�x���=�]JO-�������%{N�-*]u�\ʃ�c<Wy���M2 #���s�|���n��&�9�~�_h�����C[k�g����/?��������<=\��nܴ����48m���|ncc�����e��EBD�tYض�^>K�oۑ��B��)au}3�΂7�7�16\M��A���q?����S�F�4�]>
P�C��%��8R�#T�(@�Q����QlS�^D�C������j��AD@u��0��
�x���[y-M�тN���J�j(���nF�󒗗n^��})�a\j��Gv�]:QV����+z,����y�V:�f #s#+sS3����������z7F��Y����Y����<�935[Uh�̀��,!&B#���[R�gZ�:�Y;9.�����43�43�67��4��~_�L��"���E�������ڽ/�nNn�mP�}�S��r��l=��.�oՊ��w�c�J�"��8} ��(�ZvE>�/&X�[9FT #$�E>B������	z;��6����jd*���h��E]"h��/������=n�U�A��%�{�Chݑ��mԸĬ�ŵ�._��7
߶#|ˎ�M�;�D�8ʗ�8��j�)�ŃLi/����s���0�[��9{���:@ضXdi�de���\=skǀ���/
itX�N��<��E��(|<]�͑x*�-���M'D}T1(���5�D(�hD��ٽn�ٹmm������_��ݾ*0�2^vV������<��?���z:۹;��Y��f���+�֕�7CHJ|wryhȾ�����=v3-�������� B���8"<[���y�n>�[�!�!�,��<�TH��I2Y� �{���z�ق"&�O�[�,�A��U�EH$0:	O�������>�U'�+إ���J�߮�M�4������(&��ؓ�Yݷɞ�'��;�{������-�s���'���.~;oQ�u�F��u!aK����u&d��֐� ;[�9��?�/������fkc��d���s�[;��f~�ͧ�Κana�����n���v����9ytٲ���;����O��+��=Ј���O��[�wJ�a��M��ǔ�����X����Lp�֖c{�4�0U�A3��`u�В}W
��2�*E%$���Q\v��/�cH�P�px�c�\yy75�UQ��![6�ݹu��=�N��>r7�r}])W�׈�+l���1j�Z��u�]�:�!�-��@w 
��נ����PûL����P_�@[3��z�Tzc��fF�Mt���מ�9��� �Fڀf��<E3�ո��/\diicnnk��������D8�զ}L��*���Ay5מ�<�m_y���S�Q���>x���k������/��\ɼ��x�A�מ/�}�#h����#7��Q�p|��1OJ�W�j���$�8E�nO%���%U��
�QE��c�/h�H	�a���fsԕ��/+H�:���K�iU�g��e�o��_K:�Pz� _�_���K���(ͬ�%��'6���d�%?{��,+-;O20L���m�w"��6:�iQ���F�"V}�9R���d��ff�|������G�)ϒ�1�<�in^^iO��!�b&S�-���6����#�
{ �Ã .T[P��0%J�N�����4Sҳ!�,����X�`5o�/�VE��1G.�x�aei-���ޮ+B�lZ�~��� � o�����#�k+рM���3120u�_��p샼���V\+�9%�N���6���9\
�E�Ѩ*U@�I(	�"���LD��4Za�?�=�n
��	C���Z��u�ߛ8�A���TT�P�5�A�ʿ)��n��"�#\���`��D�k��Tv���>�������c֜Jh�����cI��n��P��G�:�ۯ=o��T��k�L����Xx�F�˽\D��xGa;��;�|���v�a��CW��/���7g6���*x���u�W,Z�������ߧAc��}��"sG��6���-�7�[d��d���|E����O?��s�nOo�^X؊͛������?NNJ}���ŋ\aAQYem��Ɩy����N9Q�m>E���a?S�Ǒ�r���X�*��T��sG�Ě䚵%�ض8 Y<H�y����z׵�ȇ�-*TL���~�Ϋ��}�������U
l������IS����b��c��<L���<�U�͔�'/�H<� �;+��n�Ww�bw���}�}���!�-���``��B}�pJ�S.�����Z���&� ��:ڿ�����Xi/���`���|
�F�}�y �����/�Ydanedfc���B�Y��3��t�l�Df��E���FEյ�b�{���Ξ�^�kha�y�Μ���Wn�K8u?����B�ԏ߿_��_A?�Xf��T��('�����ĺ�U٥|"��T`�Ȱ�y�,��!�1��t� M����p_�J_�vO��8������nf�{�6[�}١k��5�ֲ�6����}���P>NHDx���������,����v壓��'T�Q8P}˩"��7W파MHU��ሥl.���9�n������2���eqUQi-PR�PU�V��U��Ig��P���mm/����A�k{�O2�� r�d�y�{���b�Z�J�D�Y��#��KW���������������t�w�Μ���߿oת���z��	A���aY��ա^.����!�V��		ػm�ų'��/�ǝH�q�����_��ݗD]�W\��Nd��]��������U��,1�ťriT>�-��D��F� b�I(r�����^ �+T`>춫:�9��"��,lk�?Z� �����o�)j��&BI�{"Ը�N����]������r�������_Q�2�%UBt4�l[l&��Xbm��"�����Ȍ�k��^�p����>��/g�,\s�qi�h���jj�B� ��e^>ޮΎ�Zs�ϛ��0h�!AK����ؾd���Ό� 77�-�W,r0ۼu��bG� ���Ξ;����o���ff�ΫW�]�r劵�K=�}�ݼ8TTXr3�^�����x�Ц6D�ʩ<%K�����r�x��M�E�����~�����I���'Y2�� P����|�H
��;0#bR�BU����1Z��f�ɵg�?kf�K���됤͂�]�l����>��FV!�'6�*�vfLF��G�7r��^�K�=�Y|���F:ȘD�Iԏ��C�}�Ӽ&Z���e��p�,h���J~ں��=�ut1�u�@�����ӟz[�3SW�W}�Yj�ͅ���3�#3-K[�EN�Vvf�F&���~QC+�w"���q��W���.jyC˺�[kZ�=����{;���� ���S�/^���e�E�CI�bwݫ,fNr!7����)ٌ׻,?t��~9���GR��*'��b ,ȗ*D29 '�z��~,&��=x!Ыu���I-�/Ǳ��*�u+��:��:��ZҋjA�������P�������[p�9��s^V�����Z'/�j���3x+��{RTs-�ED����A���x������~>�~�!�a�B�n^�1|���@��v�~A�_��)\2KJdɉ��5A0�H�GY��3��=�E�Zeo;�]<�,�eJ��'��E��f�X�7"������������7�>��5�o��6m�΂�6V��v�Κ��t}�y&�-M�Zx��X�a�ř?|����������B#;����;˫A�P3�;8*٭Rl��q�o����#2�$�TQ�+S`ML��,U��ؑ$���*Z!-�{�>�rHso���zd���(\�����~ۗQ�_�M��6�z����"���F�|��O�"|��L��;b.�F��]t���y�L�ת=E\��z�J�N�������Z�{ǅ�7s=���w=��(��W���_L�_��XLjaP��������)Y�$�Z���o���l�t�̟MԠ%>��]�-[|� ���VO���}�2��kL͵⮟]�: 0�c���£Q�֭_cmm���mnn	���\�$dYȊ �`0���32�df唖Uuv���p
O�A�;(�L�a�q��Cl�w�#���{��a��L�hT�*S�R�� �ƅ��~�|�S��{Q� v�+�:�փ���A�$��!$F��:�
��0���f������-�e��^�V�%[����9�hӁ���}�1�#�=x珳M����̟��`��6�Ԫ1�12��ʻ��NQ����݂zs��g��U�`ʅ����<#��fZ6���&�VfFV��ff�Mfj��8W[��z��H��j��nvMK�ô�̼!�"�\�xf��7�_:u8>)�؍�ә�O���Tֆ%r���A�VF?.�s��3�Z�(:��|Jѿ!T�L��� ���T�( :�A�$)ހ5�4�R>N�����N��wMSK�M[(lnIU��cǆ&'/\��uOO�� =S5<N�6EKxQ�Ȑƥ�^z���Oa0��N�~���o1�����`���{�e�.�®��̚5Y�1��Q�(
" Y	�DA%'%�s�96�s��t�3j��v��̚�����o���?뺧���S�]O���sQ���#g��:�;Jl�ÌyX�Je�3�\ٝRӟ�0�H�rPKY�m ��a�q�~� ��؟�9�*��7��Y���z�u��r��]��_����5���PM����7�_�e�w{vl=q��5݋��:7�X��{v�����������:s��	��G�F�H�D�7���J�&a������=6 �r�=B���i6����껆B�h��O!3�	���N��_!I����`�I0ŕ/3�s�g�&�	T>�)�s�]*�O|�������
�J9z����P����-���5]5�0��n��q��F�f5�J@v;鰾��+����T��rZ�
�p�C3��Ú��̾��ɓϓX���7D&7�i��SgT�Ԏ?��M��C^�V��U��R��1��w:~t��u�8���������ᇾ�7����_��O�ذ�[MU7�/��j˖mP��xQ���,#=����Ǝ�aFQ�14I���8bW��IQ|�h�W(��:8�t�D�dPAEXP�EhP0�P8B�'`y�P�pQl�'�%�L	Y8	�U�:���������'��:X��	#� �d�eu��&A+}�p@���,bg@p~���83���X=N�N��a��(:����$�.�`�S�ܴKu����Y��=>�����=��ܳ�+%��~�d�6�����;�}��k熷(R�"
�w"|�k�ZȎ������[v������Oسg�޽�o��ݶ��w�۹s��m�wn�������>�v��;�ۺ��ؒ%<C6�g�����1]�M�uɥ��ť%CxzTAk\�@2�r~Y�A��t��ex!j䡧OZ�c�0�.d�& M�J�/�����)�DƓJ!Ђ�R~��ĳJ�KߺpjA�B�t#��{��s��[I��R���pH�cX�Z����a��[Z���Ӯ�Qi��W ��?&���o�@�M��"*3��K06���"Tպ���qxQ^���5��O览F����-Z��=_�;G^���&����G�fk�@�ӑA`	G$b����;
�)\>�/�{���95͋Z�.@�
�o~�^�N�gN�<��z��n�3�-M��a�wMW���?���?������z��aU���z�;�--(<6P�C̉�$�?�z�Ԗ�N��z�[8J#x�1:��i<�.G��E3�����mX>g�����V���D�40惋:"Kz��ü�?��y�?�Ns�HW��R��
"�8|:��/"��B�E�o�����$�w}�H$2����"�%�H�u/U4��'Yi'�Т%�4h���0�	n�<fLd���̩Jȩ�O�m�U�p	�dB�����&��*��u�=�!h���u�C���������v|󷿬ѽt��D�Ѕ;v{��.XE�5�6�3�a��v���*�z���ۿ��S�B�ff��X�Fetttqx"G��
��l{�"H$BI�@�?�J���i�����-���J�s+a�y�����^�)Ic�>�hH(W09ė#�Q$3�h#��"o�`���-'ݓ,�;,�ת��CP��>��6�j/��Os:�<b6��h��>+��K��m�|S��b�f~Nq)�~O«� �f����]���Xf���w��������
~�o�oE�M�[~�}�{>�Bx�|��.��*����/+g
l@�Q�~���w���I؏ٲ��TXp����}�~�g�n�~�Qs��Y�t!�&��8�ϥ��l���:fanF,���hr�P@%��ހ�ó�=��	��{cUD�U�:��%֏�Iߐ&^����EȑN@r�2D��i�����U4�s)��6�m��P�d�+��pPaA�}�GH���$$���H&`P�D���`��(�M��T(�ɥW>�1O�3��?�y$���$� Ѩ)�틏���Dx���-{%fx�d�֕��T�Z	��N�ݐt�"���-��;�/�O�>�<j��"���9}��!�������TUSոx^]S]MS]]]9�k�~��O�8r�о#�B��e��\ֽ�~�䑣�w�=q�w
i��?m߶�ԉc�����������"��"��RP'ox��Tލ,��`iY�$�a?]�X���5J�	g��)�h
�����6�q]�%��N?pӿ�����'m����8�Ǵ>��H�C��'PDo�%���J����ω�����&Bą$��&r�C��BC�a����q,[�q&!�k,S��K�4!��A(,y����ooo�lo����/*(<u��ɓ'/\�8z����--L�u��7}�ٟ��fۖ/>��/���O��0�57���9�}�W���#1�Y�ݗ�FWML�Tϟ]�n
��c�'O���a�����t�
�����m}���^�?�2@e�cIu8R/�M�\J��|YڝT��\�]7$9���9&��-�*�6ꅆ݃c75��.��/Cw�'x�af`)�h��=�!4��,�,��ٽv�Ã�ût�B:)�1�Q9�|񓠅<���G�5�S������,�:��~���Tuv���LIp���o�JkI�gn�~}��w�5�mڹe�7oQ$�FP��*FG�7~����m؀�ؼ9�w���;v�ة(�v�ٹs���{�]���nڸc�׭�/�lٱy�֍7oT؀*�� ��2����[�}�y�߆�{�ۺw����\���7��o?p�h
p����70"L�.����,��<==�7�/�qM�PJ��~��_�q�����#�7��I׼� �μ���eN��WoE(��Os�'��r=>��AD(��1:�%�A0#y0�y�!uA���<N������E�
�?М��^̳�<ׇ>]����:�Zv֖�wn���&�q!��O�ß�G�GW�7�f��zG�(�$V�u�Ey5���U�ݍEE�N��.��ki�k����о��s킮����i�K;�8��{���enYac_a�h=��P���i{�_"�1z����o
���Y��N����C �	�Y֐��Bd��/��;yN㌪��s��Ν�uV
X;�����Z�_��o���ۿ{��][!���8~p��E��*g�<�o���͟�����~���O?v�|�3��z�{�P����!N)���3�@�-�avǋ6f3�MFG�*hX��L=�:���e�T�aL�8E0]�M:axttȀ���jjl3n�
�މ:��"QL�4�@2��v��1R����+��X����~�U~"��t�̏D�G��)<,���qa\Ed�!$���D@.�bx��Y����E�3�4:�NeѨL*	>������~Nv6�AǏ�����6nZkgg��p��Ջ{w�W����k�@#>�EG봎�ٓgv������u=G[���>���?��|���M���n`r���՝�/S�gj��d�wPhA]�o������~q	�m�X�P���]S�X��,;�5�����;˨����c�����Ⱥ^���y�(zs��i� �;�픭�a@b�$�o�h����lz�3�ip=��̃�ssλ�ܯo?�(o���b�>�{=*���˶�]1s�uu�pbViV~�o����[v��~�5sӘ�x��ǥC�A�lp�n�Z���4�b���v�]�*g�ڍ۾ݰ/� �ۼk����mݽv��o6�Y�i�ڍ��m>�^�;�ް��u;�Z�Kɗkw~��.ȗ����th�֣����|�=|�����A|��u����PܳoÎ�P~�n>�͖C��|����}����+�!�� �G��d��%���/j��94�5f��WvƖuئ4�́l��M}V�)d����3t�!Qb7�;���5/<���!_:ɑL��3�,E<H��!t�2k��ϛ@�4f �5 H^1&_�HśEs!�]N|^�����S����^7��E�Ծ�~I[��U�&F�Fz�t�B,�Xߴ�5�u���G�t�z�tcS���JK��k��l�o�9s�ʙ3jT.�jh\�3ҽzrB�®���i_���Q�Xى��'t�$�M�V/�9�l ��[C/��^㇩���I DSs,���*�m �e�-ER���P��Ξ?�r^��9h/��Z�ZzZ�t`tzAS[S�ʩC�v�ٺqז{�o�"T=u�쉣Ђ{�#�O޻M�����i�W���y5XN�R���������y/B{�d��z��6�l�A��;��-W��y���>=�o�B�p��>���H��7C��$`����q`�ᐃ9�l���3�������#��"d	ފP�"|_>���*?�>�o���qKo!2���d��"Q�B���4��y��a�Y�?F�@�D�BR9~��⦩�~EI����=��9�g��ͷo��_v�{��ᦱ�����_|�����13�55���>�m�׿�ݚ��ۣ����^��c~���e}�;�mذ�/������;q�DbBrdD��=���f�D���9�&hܰ�������Ȅ��Nn�]}��e��tQce\�K��+V�w�h�\�����˵Nz�r[���y�w�'V���UB_, ϟu� �l����U�Tm��2����k��;u�>�!,�<	`뿅Wt?s+/J:n�1�+<�bCkzFa~^1t����a�yQ%�4�qJh#��3 ��9[/������yF�����io9���(¦�6� �������z�o<j������w�*d�~���.}�W��=Z�^ܼ��} ��im�iӡ��N\�q��ΓW����q\{��{N]\��غGv�ܧ�����ӐK{O]�J�=���C������{JW�G�ݧ.�:�sR��aP<_��(EH�q���=v�����.^Ա���Pۜ�]���� ��s�W��E�ADa�t�j�SV�]2� �6 ���fBC�+�)�%�b��!]<M�O��V�a���(�M2��A��v�u`x3#�)w��C:�U�\�v=|N{סc[w��{`����s����N�9}ɥzp���?����/�ꓯo{���1瑘����&e$&)!nϾ��ٵ�䮃g�:���ځ#���ߺ��=G.\1���������d�Ŵ	�����
5o{��eW]#���(��m���8l�\ �B�D�hAxOlr�	U��ϝ<}�r��
r疥�+[��fF״5�N?��][�C�ݏ�=�o'�����a�?.k�Y�_�����׹tY��e��G�i���sv����"Bv�e=��^1���1���1q�n,�'�kن�����0�EΊ�1��:̍��2�פ�W�{l�wm���am�"6�j��m��K{R�/�E��A����cD�6�>
*��!�ۤ�+K+����?��R�Jzӳs��K".$��	H2Hd�ʤ!�Ie���-��OD�e@URj*JE<����Ϣ��o=���x�z����*g�\��ر���;�^�rv����qd�V����6{�s?������ҥ3�v�߶c-T��ک��P�HY������kh�]�v������������FK[����P痮���{r�o?5��-��W5��߅���qiys}l�K_�3ڪ����Y��'9ꜹS�<�ﲍ.(�Qsy�Jn�J�+����7��h����N��cx����5w���@	n��'��bN�w��?ŉ_��gܞ�̯�"������ޤ�Bޱ���j,*��jjɬ*��J�&�D1��ȫ����/N9�=o�V�|����sf=4��?k�r��	}���w�j[ֲ9r��������t<wi{m��ܮ����K�Gu�O�9��sPӳ׼l�q�鬞ñK�/���~����y���&N&Zf�T�!�l.ݺ�u�}�E��I��A��N���x���z7�������������:��G!��ZeS��s��6���Z;��z���{��=O	/i1ϳ���o�QЃ�1�"@�#�g���F����kΏ�n�>M)Q,]b��� B�$�eK�����"�!�{dF3N(^ �� Z�.,�:^6�IBMpI�"���o8yR���W��?vL]��9�����ջ`h������/��_�T׼�g�����v;k�l�0|�5��O�y���y
�����yˮ�[��~�g����?���/������/aؽ~�]�[a��z1TY�̞z��Uk7�G�V^���}�I:>I�|c�c�5B���-�#*FG!D��,)F�P��O�SUU�������Us���7l�,�n�^���vƁ["\�?4"���/�
o/i��er���@�蚾��U��H� -���(<I!B~�o��\?�'DB�KnO��A	��	�����u8�^�X*�!w���c���:�cȧ|��a��F�-���N/M��,�$?!K��"|�V����?���`I���fB6vt��)��"T̫<�E�CF��1"Md(� �XЅ4*�g�R��!� ���r�.��F6q���������ĤgNV淮{<p��UWW?~���ݻ�_����*G=�;>��r��Ի���~��MS������݂�n��_��o��O���_�Y�_���~�ɧٴy���`˥��{�z�W��gf{<��70DcM���}þ_}������c8�謲ak��!��F�{P�|�����(����w<��<Ὁ-�)�a@!����Yz�KXA$w�%jtFTa��2 �j�=W�K�e�W��
K���y���U�h�AdD���ܺ��!�t�L�@f��C�sC�>�j+4�A��D��� mqvb� ,e�w�#���k����K�
���S���^�x;V҂o�I���&�-)��^>�"��Y׼�<�kb�(�flr����Km�&A�)�-��VV��l-q�
7��Z��-wR�C�Q�fr�3̒1'Z���~b� ����1�P�>c��l��
�F��4,[N#i��E*{��^`s�Y��pE��̯N̽���Y7�-��kĐ>K�j�{�V]��I�|ջOP���:>,}}�K'k>�v0�qd�7%юg��a8� M@��!�XF����(E喇'a�K���E'�y�M��@0��;�hs*>(�re/��;��/����q]3������۷��m?t���S:ڪ�����t�\B�D.C�^�~���HKWO�¥�{�X{=�A�S���b�":GN��+�O��:��i�ɯ���C�|D��m{Oo�}LC���?��xr�me ��M�[�
Ǜ@�g�Hb#d0P�o�xǓ�24"K�\O� ;�{gϩ9|LUE���L�����������r���7�;�������Ś/>���]�5U�����w_��E\�F��^�[F^nvN��o��X9޵���cbd�{I������E$��Y#LN/����k����Uk�VW�z�ӎ>i�1x�����.�T��B�bO��K>�s��Y�0��ꆨ�7�1�y��Ĩ�:���3�xn�;�d�*]��MC�),8�� �AQ���� ��gߊ��b���G�C��a�����D��cT���1<S�gK�,�(�;J��\4��#�	d�*BrSߦ�"���͘T�B����$РD��d��,�����T_U[^U[����"!*)%�����]sS����Սtl��#�e�$�]R$}>Eho{���9*�IZʋ���Ϊ��8{�ε�z��4��T`W����]�;����AO���gtv�P����,X��6��r�Q}�k����}9��i &_�`��1)�f���Ȅ ���ÜEz�R�[���O�f/�Gfg6������U�B�oe,�x�?��	HBq�e� ˔QyS\�H�,�h�$^��.�R$�
�;	[7����'&�>	3��?g�e�u+��u�i��s��.�Oz�s�BcŠ�GZPϠ�PI+}��^�	;C�L�	�A�D7c��5o�i�YI�a1f�S�K��DuO$v�.�	l�	�q����R"}�Y�n蕀�	��]頍���(�|��)0���R�x˓��}X$���5Da��4���H�� 6��,�3K��RXt�"����-q��dET4F�ό.,a�_�.���eU$}�f5�f��D�� �gE�4- �C�R3sA�"��/޼g���Q�C� 9eds����"��a���ջXS� EX����=șk�r	r #x���)�]P6�m�7�<މ����U�sz:�D�օ��!���3�p�)�!�YL�˨�����]�n:׬�i�;s��)�#�� ��]0����,1�̑!(2A(�O��0�P %���%�ɰ��_y�<�z�B�����'���{��I(�+�z�7lط}��cg��?z`ۧ��o֬����lX��{�[�����5���5k��W�c��ul,�n�0��Ѻ����y���5u]����5H��`�0Y}t6J8Q҃*l��!�H\��e:ga+"ӧQx!K��]8���]8��LJ��?�9JBVq��~ �Es�aSo3 �q�W8�
Y��*]D2""�T�P�N�0"�(·����&���Օ��G���Q(�Q:��D�و��n>���W ��EC$�(Y<F��(��hr}>������dHd*�����'381
��E��	&���0��ݍ��遏<<�{���+cK��Wu�X�
��9�g׮�ߟ=q������;fvwo;;�|�)� ��Ј>�n��w����]0�a��l����$�IumMWO�L�$�<�/��U��?Jȿ����QX�����K|i�D�	��\.�h�흡���RJ��؂�Q��1�L	��I)R��L��x��"I�mN2&X����_/���'Vpt	F�9��JY8D�����xȗT��#9D��	��,T��a9����se �k��!�$��<!�) �q��	�`�?�s�����$[���*f
��K� T�#s�����U���
�2�h�'��q���s�"���l�,��	�X>�$��ϭ0gW�s���)�H;O�(�
�:�(�`� ��cTF?7��:>;/�b�Ʃ	�6Ad,Y�(\���VG��nu##��8o�{�kS��-�/E�o71�Y=4����D���d��a�ϜeHތ/ة��ؓ(�@�g_��_S�g!4)�>�'"|�VF����-�;�(�z�D)¤�nw��5A���I5���\jG�3U
�FM�~������������ڐD��oJ^�Ӈ"ܴ���Gw�2İ��"���Ξ��=�������Č���2x��,��)���g�?��"D�����������1rP�ϋp1F���s��嫚�v�޻e��{��8�zZ�k�@�lݸw���7�^���r|����=6���ꚭ�KS�[Ɨ��ݰy��|��u_��X���3-u��'O����/,�P�"d�8}L~7�3�P%�L��;���y o����H\}"nظ*�o�ۇ9�+�;%�^�.k|^�BG
[D��?���H���$E�q(��N�H'�J�G�R�|&���5=������(��;:R���G�XD�$��(��0Eq� M\�:\�:
)h�F'e��2�C���R�Fi��{��8�X=g���U��;a�j`�TTV7F�rD��,�G1�ޑ���:4q���=1)�徵������e=5������O>ټ�����ͧ�@:X[Y�]TWݹuӧ��y�S��/����^�V�pw�u��ʱ-�֫k��]�6�il}�*=+=������������ohT �����>/�MHI�B=�Ӵ#�Ƥ�\*�'";m�&�<�
"����!���@��
A� �!^�E3GH,[>J&�i�e� �f�E� �ĳ�� *P���^CD~�E�D�T1g��h������Β�'��Z�E �7�ѥ��N�{TJPRaV]e�Uq�(�u���U�495�,�s���x�81�izLL�Ӕ
��������������Z�.��w�|~�o�o�	���ON�<����Ѐ��@� �GO�8%wr^w
�G|Q�TXQ��}��VT~QhAEHAMdnQ|r\LԣG�{�5��{�>w�����6�?K�q��urj��K�Ή�	?�ILy@l}b�XrvOuq�����Ե��炢�נ��o���\Y�^%Ҧ�(9�2���x�W|`^O, �p�ɰYDq��d���`�-Q�o��ɸ� ��!�
!�b�s��}=v\)����ˮ�)��E=�3F����)�Ϝ�o�]���f瑭P�*�4�T���C�\��(�\546}+½����u�c ۊRa����9UqɅ�Q�>A�YE��)��(�mE�P��a4����P 8ſE�� t!r����T�����	>��ۺ瀳��m���vݶ��Ο=�s˶C��������_~����%x���nx;�y�C|��9�:��F{A^T=tQ���M�����7k�����Ο9{���ӧTҲ��Ȥ1m��@q��$uj�(����D�C��p �f�X�%�,`#A��2�F��H���t�&����-C2u�4"R;	Ǖ˝����B�C".�� q0W��a,�s"D\�l���|�U>!��22p������T>l���~ڄ�����7�]���j�*X=�Ҳ	1��\��p����[IGu�5�f0<����������$�����O���}"��'�F����><��7:���v����ꆾ��K�O�;~F刪�	���N���/������ɟ~������7lصe�5=ݓG�|���~�fͷ_������/?Ӻ���t��〽{w��Śo��bˎ���;�zJC[��m��`İ�B(�����~TI<�g��d��4�#��Y�8�"�r.h�U�<iUwʪ�z*@ EH�7$�s|Yy����4S0������G�pӅ��" �BHf�ҽ��e�T12� ���]4u��}�/����gNTr���cBYEE�@jyU7��a{G����ZZF!�E��M��Ie)u>��O��R��<�~��]����eo�"�B*��⨠Rp �85����%����
�;va/�����0_UQW.���̌/N..Lr�Xۢ����g�}��-��5�/�m��F���.�Y�D��Ă�θ�L���==K���'%g����ۿ�˨�_�y���+�e[YfysQUht�{��ht`�x�U�J`Ͷ4���i!�c�l0;f� ����.r$���W0Ԁ� ��H�f��1>G��V%(D�#�r�IH-��p
^P�kO6��`�;�
R$ۍ|�S�3ڈ�cW�v�f������v⥛����u��YݳWn\6�mhz�����[&7̍�n\73505�nbbddbf`j~���Ǣ��m\}�!D�r+muS���eU-���\�np������wl �/��;~����bC�$��.�$+�נ���.��4	�93D�+d�Q2�L��,�,2^�L�� QL�#�	�)^Γϓ�Bu-���=�mٲ��/��䯟|�����_��g��8t�2���������������k���wk����X���o���Z�e�"���z͚[6��W=�ܡC�N�9�:4�N�A!���ƱB�@EN�͑�3�,�!2L*������UGl�QVX��S�J�} "K�P�?��^������)D���P~ B�r�zK[��D�E�(��|(¶ޞ��t4��c�a88HҤ}�!�α�)�@_=~v멆>YEc��R�;�*�9]R�0�H�*���d=�2�Gݾ~����{��������{v.���W��f��w���;w]=|K�+�k�����Dņ�;Yþ������v����*����u_~	-x��QMUU��wl�]��~����w�C�x��=y�Ⱦ��Ă������޶Q<:�E�y�KVN����mG�=�a��w�Lgah�^	تw/}�<�M(��%b{�5炴��w�)H�k� ���(��lB$�3r��4W0)�M�y2�+�qEO�����ߋў2�ɜ���D�=fYBD�F��X.'�y��s�M�SF"b�XF�%�v�>��h� ���/^�� ��!"4�8���Q|`F�ez���{������a>�w����-恚�C*�/P3�2`�\�3��$���=-=���Ay뀞�_3k����a�^�\��UQ����1��p�?+����ɤ.Ʊ0����]�j��4��Q \"S��_ڻ>02�E(�Ha�#+%�����!Q�U�3vYw�G����3�;
�X=���vy"[���`�8�D�<����.���X�<�� � HJ�I��?�KH��r$A�r�LB*� J"9 ��h��������Bu��!�k��UTn���N�$����0Q�B�5�T�3�jǆ�|�O������ذ~ǦM��nߵ}�ޝ���>|p?����?x^Skݦ�v�Mζ�#��p9�-�F��+��^�:���~���k/�\6�r��D����}'��vt7�a�r�����0���4 ���ye5a3�E  ��IrQ3�̞X�	��V�R�	��P�\����30���sFU���sǎ�8|��S��_��~*�1�f%�1����5߯��"���ȶ]�<�'~��o��_q�M�e��������˷��nܶ�idd��(����x�(�(E��a8��ΐ��hD��pZPyrR�K���H��yg�I2.��"�������-�Y�����E���W�?�b��r��ʇA�GJ�n�@-��m��]�Ы�������{I�CS�[
����o�U�AY?��;;⑩������߬9��[B[�[2�Ee���$�P���_13�75T׻�^�O�0q��#�Y�.�zW.Yݱ��m���w`�ލ�۹e��CG�Ξ����q��$���]�sz����E�k���nv���s;LeSRasogt�K��.�k�li�,�Ĳ��T7w��5���
��)�h�"r:��Z�'Y~����x�OBy?��2���	Wq�%�t�0>K�͒��p��7)gM�X�q�T�	����	�H"�qŢ �oU�(�/������!�ф��=<����+9v�,��:�I����*~ɏ�jӟ$��5U�tU�U榫�i��46�F��gy=Ȫ��8����\�#¸Ї�6�tL���9IB���$,�?���ѳsp��-�+�Z�.ki\+h��u	��.���m�J��S�U�G;�9����QE�}�K{#��&?���q�i�~�t�y{�г{����|����';�{�G�m�r�_F��Hz�4��zܹ�<n, ����)z��m�y-�,�@�S0��	��݌��*e4���XA�̚����<E:	�(��HTD�@�ч"T,�P,�W���O{ĕ�4�w����u���="�T������,%Hy��2kF�[8�FS;cio�k�������ڙcjg��;s����G��8t�ȁ�P0�N�z����O�X�,)�V!�!2/���M�#���zO�W�Q9�wA��y��j�jj�j���:�gj�VRR��Q7��O�A|-��/�-��9�[�-������?���I�,���'���
�!�T��rl��[Z۟TQ=����y��7�?��7_�%�g���Z�ػA��!����ӿ���&�ӿ��ӿ��֍��EYޞ.���O���ϰ���~AS�ʕ����Q4���1xȉfB(B	F4��т)oϟU^��	-���2Ew�$�(B(�E��߫8�W*��*��)(�"D>h���B2���[;��'^��(����U����s"T�BcA�&�Y�t��
OX���U�ULp�#�Wn� AH%��uL��@}5>.���������n]և'�>z����a�F�2�x|mG�t~A��~Fq�]7w��>�O��"�"C���\�;z��/������߻o��m��8欖��=�K��t�����o��������o���'303���������)�"#��=t��Ҋ+���-\<+�Fzi�N�rcf�*����e]�Lu� ������u�e�U,=/;iX�sf��(�Z�<6�46���-�&�!��y�`Aĝ��D�B�<�M�拘|	24�XAy0"�w| B$�0����<^��c�ӭdO����~��Z�������D=ʫ̩k��/��/�W���[Z����������'+�v���2������g��/�?�}��8j������ڥi�id>F�߱�y���������u�*٬9������'��)���c,�G�2"��R�ڗ^�"��
y�Vq�!�tH{�x�\r����ho�������~�����Ϣ��_�EV��]{����o��h�~����gl�r1z��������ɓUYj�vD�������:�:��;/��Z����Y�+��9i��"����U'}�����c�tl��r�F9ӭIIN�!����W�e��A��%n>�~An���_m�R���������ec���7���n��ž��n�Լllf��}����%�e+`�)L*���zpB���K'�\:qF��Y�S�sz�Nk�P9���ެ�k7��Ҳ����1r/g>���RF=��:q�zDS	�b�rk�"�E���
t�����?E������b���{9sVMC�D[KG���u}}mM�c����<��z�׿X�䏿[�߯��o�������G�V;w�����K�ۻe�&mmm͋N�:��WT:8�&��D���Cβ��Ǆ��`͟�
f���`�(����<"0h2�Q8K��९H��x�N���A�3h�+\��(EH�.��a�	o�_��D�ђ���@�"�bhT)¦�vef�U���G~,?���sOJ{+B4���Q*}���1�>��ҷ�%���*H@�:�iG�1E�1)���64�0sࠑߣ���Fj�<�]?�VV�6��_[�<T\��ҍ�MȎLJkE��B�l�K|�S��Q�����{��)���А���8�T9����[��<r���ݻ��۳���G:y�8��c�8t��ȉ�&�n�ܾs����#���NށZ�f�N���q	���e���wx�	��_
�iб~p����-�k�ү���6�;}��+}�ۉ���������g�� B���l�
�&� \�@z�XM.xī �aY\1���r�l�) ɮ��d�8E,{�[)����q�p���!�|qVF��c��MmJ@B�]w�;֏"���_�eg$%gŅ��<��H�L4�	n�/�N�}������/���)���{�ݒ\��"5���A��������p�`t�(o�y�9FB�\��|��Cj&��c����E3��c���yEC�-5��:�v5���;$�5⒟:���L|loae��K=���``K	h߼�o���m<y�dkSkwG��G��c]Mc��~Xv)��'��� �%=�w;mv��ˡ�p�*�O�'9�>5/��jٓ����a��+���O�7�[3B�Kg���4�4bA��WN	l�ߣ�!��|������
�M*F0���71,XA�7`M������Q�"F��/c�Yu���|�Yx庮���u�K�n���q ����j�.��w��΃��n���<�x�vNUKUM����Ybn/�֏c��JϏ�-zu��ы�k;rḊ��+j�����<�u~׉#�6w��"_�t�ՠHM����Gj/a��K�P\%QM��,+��l��d�����!��iK�(4���#'T��?j`|S��5���W�@��ܱ�}��U�K�۶!i�������\�_���_���u�~��r�������e�˺�?p��ŋ:�H�#�dF��R@�C�!�I�˔�E�v������k�lQ���Rx�s'-��I�#@�xC�����61h"O�!�]� 	�3�����h�*��#�)(EX��G������jЂJ66�-,�Zy��Q�ˏ�OD����%�T�Ђtf?��ǐ�e��(c��A+�e��ٮ����u���"��
C��n8G�v3��3����a~'y�a�_�Ϭu`r�{KZ{�<1A(�i�9_6H�v��i��m(� �^��W��S�И^T�"=M��h����?6"�l{ǎm�auxh��}{�ݳ�^�A���>~i��屩�Ʌ������}c�xM:+]i��ŭð�VQ��)��a�e���6�$��eT�$d�MH���z�P�r u���w�t�cucһ(��-wB������ʜrz�w+(I��?w���|3�D�f6Wȅ&DDȣA�$?�� �G"d�&�	]8s�^l?DG�����:T��*I�|����#�QvG`����(�ؗA�!V�|���9�D�DgD���܉|�\�:�Sb�����(� 4!MU߰z�������s��v2 1�F�nC|\�����-��b��t���҅S�m�

Z�J�L�R�Q�bOھH���9D�}�����;�}�3�i�ē@xbECEc~N����Ύ^�>*"�0-1����G������hE5��W��ԦDh��t0wx<�ZP�}� �go�S< �+:�;��N�nޤS����Ђ��%$q(\��wE�<���!�5w͟��Cs��Q<�M��e�hf�����6T�'���9�;��2��<������������������&�לW�35�-���m��6��e�4t�W5=�yPC����� 0:T�U;�~f���5������>�y�VQ];��;/�~���r��VT�KFH#� �i�F�w�5A8Q�'�Z"�#�h�ͭ��>�c�A-���T��4��h�k��^���;yR�˯�)�������o����Z��_A~��?�]����s:����.jjhkj�(Q=waㆭ𞞎��a�&��f���hx�`|/�ʷ0���]1���N3�Y������C��.$��̲���2��3��ַq�Wt�o|��w�!�g�I���J�3jz���e��JBQcD^s� �&���b����k�*!��#"d~ �֥��0�A�G~,?*����0�5H�׏PZ��oH�<(^� �W���>ѫɛn�b3i��>{�#��C��+v7�^��1u�0qб�w/��+W;����-8*�#fL-%S�,a�e��Z^�OfQXh�Ol��hnI���bacs����]���wtt�w��������!!a!��Oâ��cC��'��ֶ��v��t���4�:1�>"o���t���72�7��;�:B���4��/oh9��w^G����5�/�5�~�ofK�mQ�$�,��Q�_9�W�ᴲ&4�z=��u��{/�b���@L��Oq&��G	�%��-��P2ϯ!��T4)����+��{yob�R"��b��r==����ʆ�S2+[{����_�y{�xv�v.��KK�{�|���ӣlT�'�6��5�����{A�*Z:ucLUߜ,Ѝ�<�{;�l�֍�>Tpҋ��Hϧ�Ζm�W�ʄ��ɣ6���R�R�"^\�t�h@î�����Z���/�BC��m�B�z&�x��JX�|��Q7TZ�p��vMd2�)�鵥��֏�,m;�q)�$����2�89J�⍒�^� �ܪQ � �fFxo���e��Gϫ�B�,��k�v���KȜWN�""�s%�cw�3B�	Z��B*�'�P�B�2o
˝��J*b���1��)�c����AM�%�i���.+���"0��Ǝ��!X��/Ⓢ$FEu����Mg:��.�k�сf�h����{���j��U��:��K��^�3��ݳ~��?~�ͺ�����t��b���a�+�ٍZ���~I�^q�)�"��i���Y�� �d��*�	�Y�9^�@L�C���Y2W�k~���Y�-��;s~Ӷ=04T�w�у�N�VQ߶cߟ����5����߬�~�����o���5���ێ;s���]��ۓ�ԕ��{l��#�:�P#d:m��Y�
AQS������"|r�Sh|Hf�o����/�v@s$�%\�r?<�|�I9N�+�Qv[��R�o��N�7�E�0-��}�V�fJƧ����2�?����+�>�����e(Bd\!B��d�a]C��ʛWo��
��G~,��D��9B�B�Vc�0����#J�Cl� �����(�a�+[L��Z��� ���A�l;N@������g�	B4wv�)�_z�pf�%��cͮ�L�~�E����ߓn�oj�TT[��u�>����ͩ�I�ʋKM�x���? ���w�ٳg���III)))���)�)��I���!Ѷ.^���i%�����m��O��o9��9��u�j}����sz&	y�]c��QLrf����ؘ'��ۻS�vp�_b~����Ѷ��a��Cv��g�9�����N��)]��'����+ZD����}�N�t�2bNA2�������_D�օ�#B���p��H(���twa�]����d~�?�e���C!N/�-�y<��5�_/$;�Gx/.�%$���E���A��Y�\��הF��7��O�_������9��a.U+�����e4����v0W�t�i�S��:���#?m�RP���������e�(�ۑP���A1I��aA�m���������9y5��Y6vn$
_$���awK�S_'����|㮅f<.�+�,�N}a���qL�����l�2�����Wd4a�&�Q����lfӠS`�(kZP��Y�?!|%P�x����?�� ��
��8HJ�,c M�����N�.�-*ʴ�s���}��f�k�8���k�c`$���c �&3}�F����V�l4c|�*�� ��"�c�����?��K�S��fס���r�ҵK���i^ֿa��Ԏ�@��W`�ӈf�dT���+�9�8�2�X=�,�'uR��	��D���"Dr���7������s�;.�T/nܺkׁ��|�������~Ӯ�wC��������5k~���}��7�>�j��?_��Ͼ��?Y��?|�y��'��?��7�9��7̭{���[�Q#T:M�a|��9c�����ܡn�Lf��-�'���"���QzM+��U��	�6��״y����w�����R ��7���F�=� �M\�4G.�Z�PX�+����UX9y	3�ld�~�E�\��Q��Q�R��:F�a�,��f�1ld�E�p�,���r��#Aζ�N"p��d�5�b����XS(�lY hD�L�TV���	��1�%�iE���nљ�M�Ė|���o8���Yrj�X�Ǐ�GE���^��^�(���<�������<
~����U��]��S�2��i��<ʬ�'������>˫)jɬl{�Q\����"r��C�_&x��ZXܼmi��t����O����蒴����m܊y��������Eה"Uk�*�`x
�V~�W��%�P&���"d
xL��.��b�?�X��G�&�.�!�)Eh�E��Y�TQ��[�����i��v�����u--�����A���?nw�M�*kX(�x��x�*�,FU1W�hS��W�����8-ǃ[\�9M���Y	�5�F�q���-n�ʬư�rk&�X2C �:Gh(��q5�2:[ȳ� P��ÃLQ���C�$�D��bM3R*S��NpE���T<N#hT<E����ʖ��ˣ�t�X29'[�	PJ��dmu�9���H���M�B���jcs���u�?�:|{4+o�O��{*Y >S�Ȓ/1�`�A̔���s`�>�:BGF�f�`��#���&0"li����%����n2���mFS���>2-���QL\nMCfU�gh4I<E���s�V4/^��RJ;�7�}���C���>k`����l>���E5}�owӺn�2�˔B���Y�pϟ��A#�yda��C�L+����Q�h�,��24�?B����
���\1���?yN��	�CGS�w����Ƕ�>��������嫿|���[��~��w�I^��ްu����9�c7�'�}�(��gɃc�12� $��d�4[
|�JL���Ƶ�2�zV��Ǖ[�>-�`��o���a?>��"䭂������{\m�Jr���)���=�l�zV_/-2p#��7����l���²�Yo�P�ZFr�2��n����fS�������WE���L��3��/�y/B�J�����t�A`҈,:�M��84�AbsH,�"Ͻ�ȖB�q�����P�ЋЅЂ��Ioŗ�a]E��!�bi8�l���M-vy�Em%�A��Z;��K�%'�=����IL|y�ȡo��������t.ii�ݳ���<;����.;�2��>��1��1���i�ނb�Rԍ�B��a�^�O�uVؾ���0laC�`Q}sI}sH쳲�Ʀ��̚b���O�'w6`��BZ���nD���Q�mR�ǲz��tC�2��!���izu�6���X�b��P�b�r��Dx/�����,�I�3��D�x��&zg|�ˢ�	~��酥�9y~!�fw-7���G����q}�e��F��f�Ixً���E6���,�t���;(�֑ۜ�v9%}o�A���{2�D"M��s|꜈=3>19$@�Ȃy:gY��E��u��va9~Y�9@��	(�QH�_�HVS@��s@8�(�-���|�����l�HL6Q B�'����i�
�x��$�_:�@�P9P\���u/k��=�Ϛ��6,�˖�"�!��/D��E���B.2@Zߋ��_�%h:��8��,�4�}�9H�W��Q��.6Kŏ��6���F&���sx{?,���N�t��D�l��i��7�`Z1dH��q��G�dm����v�����F8$�zE�|��b}?8&����s��h"<[�2��"{%�mP�0�
�#�DD8� �h�i�Ԓ`��<�͋�*W�kg#��:�M����!�T�.���w��ٝNn�}b��Ӑ�N�>xjϡ����u����Ƕ�?�}��{��{X��{��]3����1<Ї�Re$�G���S	(�䡄 ��x; vT2�Wf��X���$�B���2�y� �^i�����MDr�,?��wbk�ŠUl_6{g�җ s�o"���Z�e������.��Hໄ|Q9Ȓ�E����q��c���~����;=;�8�P)B��Ga�,��"�G�A8T:�JG�����C`
 D�I���RC��H�Ȟ��M���â)Hr}��;��	�Ԫw\��w���̀�9-z;��9Fnk��ni�).�O~Y^^��������q4��Ƣ�
��9�>
)�h,,��k�j�l*k��`�[7D�0q�Jcrj_2ճv�k�&IH�ɓo� T��0M8NjMg7S�&�����,NWXΗ������D����K��v_1�q���Y��C�[�bM�#�eV��| �Hb�pJ!B�bɨ@�X������dQ�'f���]�'e�F���9Ĺ����y�|`fUb+(� .��?"��ꮚ���&E��Yp/"��EU;�����j�Yѭ�+�I�E�}D}�{�$a��� ��t7CȒO�����_y�Pe�@uQwu�^1y+Ս�e��%eU9�a/�В��	������7���oP�E�d�80�o`�3B���˔)��1ċ��M�r�B9V<�Oa$��l	=Ʀ��4� �  }�R@�1ѫ1�
qi�`��1�ʛ{����'�<D)�Q���O9X���}ߋc]0�m�b|׽6��  ��IDAT�ex�!������b��5���0�I̭���KsS4��PO;
5҇!>�*�_�Ժ���R�H�E�zFG�<o����v���rb�������Ξ���l�X�#��n�LJ�2����T�̈́4�+�H�ݔ�!fA4D�����a��)����A|���)�HR�A6
&�aDH����l���qX�7��U�V�7m�oB!"�փ@��^�p�D��	�KGT���>��{����S�R=|����*{���u����v8��ࡃ��:v��	��'�k]�
OF����t<QJ�Ȉ�),}�鋊���A&���z�X -D��+�W\{��i�@����t�r�X�y��Aѷ�V����7�Ŕw���0R��k�.vsߴ�V=��͂�@���]��,|(ؿ�(������f����IL�E�pH�!��AT�N��i
29
��i�P�D��a ,t�R�C�����hf@<w�-�EmO�y�?�� \�_F�ִbY�F;���;���]��PX�������.wmڛ��$JWk;�J��6v�4��[T�ҍi������z	-(N+�W?��4u*jC�=˂L��٥z�+:�f��͘j%Ɍ�C�X����`|���>�����y�H�axD�X����*I�{C��4�ǲQ�%��M��r'!��1��`_�w�%s�OD��M9�^��+���c��xܿkdln�^���ǖ4=�/s9�cxD����ݣ��3��<���#��+�G�	�Ok�5�W�����M߰���9�-�ӽc�T$��{:��e9ș`Rf�X�Z��~-M�M���F��޼iU�9ֈ�O]���f<V
����ՠ�c��@z�-hG��ќ�1v� ��u4����;&XΣEs�x:uD��_"�F���o<N;�����Am�{�# D��i�f2�Q����q�Y�S��ה~(BePEL����S�Z�d��) ~U�=I��_4�����絶��5�c}]u�)1�qO�ZZ�2��?пe�geр��yNc�Old�`���4�_��\��\��m�򹹂�27o_�l)h��'7�>Lp	�ȨBW�rRʇoދ|�XՅ����t`�-���a2S:w�A�t��)��� 9z	�.*�+�5�^���
'��=*�8���#pz��΅k��u���Je�������=�r�:T��W�;���ʞ�j{��C�m;����݇�C�<xx��C���߾o����w�߷c�^n�wB���Ln����52���g���L�Y����Լ�s�WI8"���oz�ߴA�'9>=�| �Y�)�z�E�좍�k��v{��\��;Fߌ��8�g�Ծs����j75�>�j� ]@���G�_?��z��ϛ@�+r��w��~/��斅����'>��)����Ky2:��P?F��a8Hf����J*�ra\H��(4�).��|�G� 8� �;]�AD8������	�{E�0�JmÅ�t�ѳ�x{�����'�8~�݉�w�)]C趞�����ښ���gT�J�0�#4��+ �����{�'d�W�����	$�
æ�'j@q/�߿l�O��ى˖g�۝�b���-^E�8� �
�Q�c�Y��<��f�i��r�!A0�΍��F%3J��EȱJʽ���Ez���Od�{*�K�1�6p�I�	�k_��܉1����<I�����E/�����L+c#��H�ȃ�Y�*ȣ ����z<h�����O^x��ހv��{q��-� -H���cl���`�������U6��_�$��q��8kA�"���}m���2�#��q&kvH��#]}���(�?�8���i��}��ݰώ��~t/�(��54�:����u��Q9F1�M������O�o{�Y<��8%����øA��gx�ٲ�;�� ڂ$|�CV�0(/�D��"|�I4C~�������"�͢2(TF�ʖ��lĞeNj�ء��0�[��.�I F
��_h�zP9�5p�}�~��e"[�T�]�1%2��~{^JndH���q��^��>��U�񸤶X2)��o-�,,��/��/��E���gxy;�<eW�g��^sI(�k%]��W�ǻ���@��Or~�9�^qy��f�PҊ�J�;"dH�I�����T�BE\�ȶ
A�`�;��0��b�P�:l`�[7�v���&�4�9�����/7o�y��Σgv=����m��(�y���c����]�}�כv|�y�7[�C�ݺ��m[�m��������bݺ��v��68���E�5��ߩ�e�D�4�un��0�Xf/�򧇹�1�d?K���fW��)$1�xJ�=|b�)`M�&A'm��4��E��1e���FI^�J ���1e�4Ys��=��]�-�����9O�Ş�t���YhA$"lm�[Z^|�j�cf���'�'"�/.��D�Q�B*Q�"c�J~`AD�
��,$?�#G\ȝ����Y�$=�'�-���4:����=ͮ	H.mÉ�q�N����Ѻ�Pm]�-m����ֶ�5}=�$M	��|���9�k�$���X�O� �a�xI���M��^�Ø,K�ЂVLI1���n�% �T�
F�,=P��GN��p�e� �%ȭ"�V4�C� X�V4���6L����b����a��A�%P�0.�V���|������y���s����u.�ϭ}��������y�<��>\<�@Zm𸊖88���b� :��FAq�������BCEcX#�v7(��+�
���.p+��8��8n���>�P��۩^�f�>I2$���f����z�^I-�5���[/=H���K�T�$Y-�������+^�������8��q򻸉������45�(=�蛂�s'�?��� S!B��B!T&e�	g�ܒ����l!l���$��ao��9�g��d��'@-abx�@V/M�=�aj����>!hg/��'m|%/59��5)�3�ݱ�el��}���lnܾY�\�c�*sâgf%	C��%�M吖�Җ�b� {qn�o;�s!pMl�d����1bЈ����;��(1TopfSa*"�E��+�q/@��/�b�����߻����ٍC�.�1��^�ˤ��=*_n?���3[�l;zz����E�u��G�o?�n��[C�=��|�a�כvA~�u4���o������n떿���G��l��$��{����U3ƚ�p���Y4}E�G1�F9�(�4Z0�¯��K,z�IL{׫�v(�˖N������,`$o�b��4"�����������e�T�#��np%����L���g�VVW�(��a�Ѧ�΂�2�]��1�,��hD%�g!D�[��t�r�P��F�eM�Y�h�<l�G���xyF�F�hD+��/*{}_�tdDiA�C9�8Z�0������.%5���������KImk����A� �ݎ�����$���q��|�[n��0{nL��Ϙ�O��dìi�t�$Y��g�|
�)#�,o��{ϸ20ԞR~J�)G�s���\�BW ��	?/B�8�#fq&���1ѫ�w<H�?��\��Ǹ�T'c���	^/r���\��nx��O�`m�L��6���P���O�?��b���RC�>u׫�*�#�8��C4FB�Уl���MBw�����/K"��-�Z�-�.JP��f��N�2�8�����I� �ڰ�Q!@M��&�Ň��=r����:�b��3F������R���CTJ������.�� D9��&�,��	���O�8z�y��\:�(}�$\y�h�"DD�6/�"q99�u�%���z@�I�EhAK���m+Z��ɘ3t�|����{�;"U�����y�w����
��rӠ��m�j�����Q�ʳ��ێ�'�im�~���3累\5su{����9�O�R�Ks�Ӳ�:�[�+ ��e��%\gii��C�'~cT���c��<�S�>���V��yq���0���!�r;~��#"�y�"��2������!$�4M�Ȝ~�PԬs��}ᰦ��[��3Wv��>y��y}3=����T�L.�)0���uo��7�;�DU����q����t`4yXra����P3�r�J�J�z�ٜ>�9g�����̞�"�Цǘsc��1�,�7�Ȑ�k�	�@����"�'c�1,�[:��N"�{%+#�y�+%��A�hDD�B$U�r3Cq�$|���O	�~[mw~��|�U~"¢��S���Ѹ����~�r��Ĕ���$��Ę$�f���A�l�6�b.��'�`���R=�����4�@�I�t�D=$^�U?����o+j�ȯk	�}		@H,l�Aq����D�@�j;A�I�7cD�,��R{�3�I�E��滏$����IBK[����'2���,����P	bA�@�PQ���,B	�P��~;w�c���X���gL�(�}ZҎ���I#��N�-���r�Kzg�8���E�6�������`p\�M(h?yǫ�=3H�Q�|(B!�4H� "��-��|⒈�"&�'���L��a��z7s���nB�4�9M�"���0DT���3#S }d%�
�*2	�s�΁�l9v<�	��]\v�N��.yb��� �hЗ��s�j�dT>$V�/�L��l}�&D�2�p�,�'�#{�����3"T�ƅHs	m���3x�V�0"X�b��tS�xp��;����1�w?䬕���{F'&�w��V�Gn+C�7aE/K�#2�2�
#���kz��$�3�8='-($���NH��@[+���%$#7�ERthTHImwz������~��M��Z�_؊�̬E�`��`@i��Vե�)�(�#��!*Pɇ��4��w<81��1 #���j������X��x����񊀷�^Q.^����n~/$=Hx�4�;$	r�#�������m� �{���CF8�:>�=�묱�C����gb������񫶱��h��̜�`����q��{��	�i�lUMOѤ�L�<S�H�"[A���D��%�_�"�@#R$,�4rƲH��s�r�h�ɗ0xbdT�҅���!2A�Q��V�7EHb�BS*}�������#�qP���~���������b�W6̩A�j��U���aZ� !�}8���x ��Й�қ��_����-���em��ڎ�^,�����亾e�IUP�y�#���.
Z���E�DqaH�����P�D��L�,���PѤ� r��Y��
*@�C����J���)�B�y<�3EH�/��+�e���t��h����urM����Bn=M<f�\2*<q�3�]BY������5Dp���q`��g�7Cʺ����zƜ�����dT��F���ܼ�Q]�yϣiCBʂ��$!-Kɫ2��	2��`���8����kU-��~��������w�?�E��I6�l�{݇)= �Y����)��r�>|���j䀸6��́��ɛ����O	+�7сo��O�ND�uA�^'߇U��T�U��^�4{!��L,R����u|"B��w"T�*�� M�2z���Ǖ{,D��G�|�.��9�>�b �|X��m����,=��t�5v���z�.��6ও� ˕I�S�L,��kimڽ��~rA_���cUNj\�����S���m�z˻F�=�,\�8?��/���AP|��wDdj	U
�?�]���"e/�!?+��.�N�6�]4����|Y�]O:|�^����:����`s�������<�jq�܍���/X)�w����T7�����7���CW����vP��뛎]�������i[�;gx�ƽ6�O3+��0���t`iR��K��3&��i,�R�)̗�r�p�"��E���V��ބ����<�B�y��R�STN4��b�,�;��y���P�EDHes!dR�Ժ��z�X|�q��������)t>�!P ���t��5	[:�4�O6��aY�Ǯ؜5sӲ�p7�����L\�:�le�s������%�G{,Tl\C�%����9}�ᤉ��[��l�ul|������l�u�wd���8���aś���ǞD6���"���H��!���I�����G�B(B2o+X�N��Zi�e` o�wN��E���5c�G��EPKZ��R (#�d���1+P�#s�/چg@|��-��u�/N�Ŕw���v��G&_=s����qJ�����iQD�@��S^OP�LR�La��k���c������7&q�z88��30�"���v�7�OF<�b�m�.�^|��D1{���͹����QC��2��la"�����f�
+*�/�ƕ�P9��_�Sb�Q#��H� ��ͼ�>�?ʜ���r���*Q��)T�! �*n�L���ҙ�BcQh�ʡQx��L���K��R��(�#�A�� y��4�E���ϴa��0�e�F��,��*&��=��4���r떹�cDJjȋԘ�¢��k�Lu�8%m#�����>�^ve{LjqFYs�%�y#�����8�-E��\d�{���=�o�R���զ\@LzjY��Ě�zJn;4��/��;���^�-�x��O�k@փG���i��!.�I�~)�Т����1վ�%��m��O��9��}Rb�q�fJ�{ByHvuy�����_�9��ф�M�Q�x�����YrgRy���=J"���
*E���~{�_�J1��ą�Ao�ۉ�wQ�ϋPyR?W]�|�l�R���-��o`8�"�X~T�7E��P@b��A���)�ѝ�$A'9�wT��9���I$}���U���h�ͬ�>9����)�B���-��Kky����o��v
�ӵDi-^�A��A����b����:HR��$�#'C�(,��"��!������Æ*:Q��Iz�+���~�,B9�;	 �p��5�S��������
�|�0{������/���7c�(�3� ��7�F����k^i9��!e�������n����ɛ.7}�?K��.�t�9�asfM����E�c�E�e�9����4�Q��[�:g4n��<��`�^։�x���ׁ;k�{�7�gd��n�����Z��0HG��!�u��w�}L]D9�棂J�R+�	)9d��J���\�R?J�����jw�Q�ys Ƃ4�<|�i�q,���DQ��=P��[K@d"���t�Q|Q��5��Y�c��ň�	a��0��3G�L��b�L>��Ǧ���ܱ�46�pq���j��v���������=Ou#��F�i�e�x˝D�+1�E� ϛ���1	�6bY�QE�Q9t�bNy��e?#B$rR�+����9��k�|	9�H��`T �I�ZЯR+�u��C�U��Fac�tY� ���Y�ή�*@��Ы�95��guޡO�ⳇ_d�=}��V���^���_����K� ׌2��	(
s �G�i*K`�B<CJd���!p�D��ȕ*֚�#Q �dI)�%�SD�oO܅/��稘2@*�"
�p8�V~��l2Q\+D($C��$�ǈ�c�Oˇ�F[:�wD�%1�dK	���|,O܆���W�z���?�NyT��\[N�+�,9�������?�6�I�����E����v[=�|�^T��]/���j��$X�(�wZ��w|^sX��d��i6OԬ��U4��P�yd(�#���Wr�d��;���b�
ņ��1�4A���<1��e*�X�a��"��"�(��?�_u�^�6!�7I.^q�! ����u
.�Li���ǈ<2`��:���;!��q��yvZ���j�~�L��1���WR-y�W0���`� �=*I���Q`���ǉ#�˓�_;�}�W]5�
R��i?�,��h�F��B��<Q�Y'W���7�د�g��K<e��p�y]����A���i��֚�-$P�Z.ϡ�p ��4$�\�� w�UĴQs(S	h>��)PÚp��@I�)��d�{B*,��܇���w����~��w�9��v�l�ϣ8�1�I�$��ُ�������1"��h���?�e�IA/f���=�@�ؤ�Լ܄�������tcs�������a|'�1@�2�h�8I��E�BӐ8�+���pQd6�݈�A���@[+�9���2�B�E���1�ly�(��zmWq��ƫ͢�w�r�-�����D���;��bTR񈒴rt|������w^��g���ڹ�eV0��s㛽7���-��x��֪��N�+��5���9����l(�{5F�ciB؇��%G�.Dt��������\��০�����p�"B�����]�E�$���7��/�Zz��Q�ˏʇ)�Z�;�+ފP���C*�����7E�X��`"�{X�"7�#f	;i|�G��L<2kn����ƞ�{�_1P-��C�:<�U�\o�Y>�5 <���{�E�eb�1��,�>�D�Ax5c��(k�r�/�v	�[��}���'y��}���/m�R�Y�0D,ȆQ��6��"q�Ț�PW	�G +��w
.�&�
w	p�"�G&qi��Sdj&���#������wu���!R���P�0(�P��]��+	P*���V�Zna�נx��U�f �_�X=Ͷ	�.����+!c�����^;f�U<"��O3(�^���U���,5#2#�:�-�:9�2���`�������Np�|��i��i����dx��ejt10�IhrE>���v��n�oh�]���<�|����L�O ���g�T�,藃�n~+�̀�zr���7��.q�>靨I���Һ]�{�>&6Ik�M���^�ih������:�#*P��Q���޻Py�\��\�D��bx���E�E<���#����`�``h4��f�0l>�˥r�������	a)/#�S^�edd�d�?��c�O�@�c��Dc�`yR,G=�4�i�P���2j�(�n9ҋ!��
�@��<k|�>F������Q��{h㱋K�奝rC��}vU���QՀ ��J�m&�?z-$��fP�g��&��F�n{�Ȇ�J�����2��گ������DN?��G���ɣT&]H�A�,!���@>�h*����ޚ�j�� ����FT�e��$�#�A!B^CK�����}��ϔ������R�$d�=2%Cg2�Lt!!�'C� �֣X���f�Jk���h�{�ijqn��`�rR&v���X:̩�H:���U��\
h��;�������ĲK��	m�7��eP��`�j���=$o�*x�@���!� �%�����Ƃ�y���~d��yX�֏�<�]8 b�W%1OP� ǞEs�\-D��!(��E�U�(�W�!Ҡ�&��݄�Y�o��ᖑCt��F�:��t BKz���G'A����7��pPp��ae�����Ns�-3|���QFp~o~�#MnB��t�I2�i�"7?�$[��4�!3�"�����^O����9��,,K�kx#o��]��bp���:��h�KӾi���w�����-���ھ{�<�*����'�Z<��+COiڇ��7�_�eu^r���%43n���Xe5}x�iV#��YXfA�(^��|	�{�5��9A�x��!kd"|+�w���	����O�����ah,���p
�-d�|p����2F�A�4�F�1�H�]�d!v�p�\6����+�۷,͍�oݼ��������YR���5(N[�d�#�Ds$W��!�P	
O�����J�|�{�œ,�$G2���Jg9�e��k4g�������YC��Y������_��V���ݿ흒Z�O��"ԣ:i!Y��U��34r�K�|��8��ӭ����Ѽr�+��ajt%j����&a;��Ebw��}$F?�>@eS�#4ą� �l�b��Y��5BY���O�����(v��["TF�o���V����=��ja���U��O��W"d�¤���YJJ�x��b5�+����U��9��,���K�,�.�溦wG��&�F�6t�Wt�RN9%�����5��V����,�u���ϖ&��o���Q�v�;=.h�f�����)�����D�l>����OX��WQ"r�=E_C mpn����L�י�p���UX���M�Ʌ>GD8[���"DV�)D�BG����q��F�JN��3*�����%P��>�i��Ik�f7�*�uF��]v
Ѱzt�����f�8���I��s���{���߲{��no]�W�nai<��*��&���)�ҬhiN�4ǃF\���N�������DZg�'�G�&>O��N(m�z��>B>d��R�4���F��cs�}ӟ���V���+C��{�?,�No{R8��x�''̼�D�נ[�Z<쐃��7�� *����f�d�;�� �d�;�a�C)F���C�����:��"�VCQ��UF��w0~�R�HH�D ��2�FfP�*�E�$r��Cl�O_6�`|��-�[����?o��10T³E8����ŭ��{�"|?	�\o���Ca���{���q�I�d�-��H'x�	�d�-Y`I_�1�R��\bB2z��_��3�j�m���%�p����^��²��st3�:��Ӱ�}�ꐖ}Rv���_���N�O�_8k���z�����V�@!B.�B
����0��A���C�1R(B����CY���n�Y��!�:(��aA�҂���U���r}G������W��X��"��ʇ"lnm/.-�����"�q���k��䚹{�a8z�-�b�(��{�U�r��s����z��>I�����AHZt�5n�5߭׃��*��"M|��FD�/���"����	h�{��t��j�3;.٤u��qӱ팵lv���lӁ��x(B!�����W?�/�c'��+ mX��[�~�?��a��卆�h��Oe/(bM���"�!"T,g��
����k��U$�
�؊^s�g0&Nm�jXz>ͪ#΃�6S��[���M��VRa?7�苣㠞4�� Y��>�WdVH\�}�0#����Aѵ����7-nu��u4��;�6�d����ցBe��ҭ�dW�&�D�7��ƍ�Q�e�!݇�.�����u�fA�����ҧ��>�͌W��
�s ���[a�4�=���3�Kf��{�?���:�#s �S����-�V N�D���9D���H^�� "|��*.�[M�#�* 0�S�g�߁~�Y��@`#Q�bA�!2$�¤�[�?(3_> �6�%L�aƫF%E��y��5=,�+�d�M��ǸbA� "B>Q��.DT��Py�[<���h�#YeJA'f|��
+���W\jG$1���U�n<�1u�
�m��(`A�"�ĲK־�m�N҂GD����	e��O�|__5 Ȩ�F�V�O�M(�|'Bn'��Ad��ߺp��~;@JB{T�$���z[/���2�9".|+����"�X~�|(¦�֢�R��"�7EH`I�R$��Kd�����W��M�p3$ህ[-�(8�FDI-s��
:�>�tL��E����"<h��j����Ӽ�{��z.��xy};��Fچd5�gN����i��F��w24�=H�?�2�|�A��9�LbA�40}��ٕ�/��?5����?����A�Q�ʔv1��@�K�	�9��̓�S��[��B�,B%��C倘B��<����7;���� ��p%O�����^��, }�
,��'��5�#X��v�R~�;Y��hc̍��<���Ƣ�_bx|��@}�{'��>��FIf}���c���쬬���[\62պy[Ex�{rڣ�	1v&�g��MS�����vv�1I/9�<��Vy���o�%�g!���ɪ�=�{E�}B�/�R;^Ԓet^�_�w��R�~�I�~({�8�$g�22��7��Y=�|視GhxQ�dE��h	#^��ĳ8��(���?��%}�t*V�#>#��Ȑ&��T���P��	��@� ��R�Ģ�FS��1&��3_L]��Ʒ��(t���]�k4\5���̟�dw����YaZ�0otR�(�̨@��K�|1�'�r�B�!���
|�i�m'`��!G�����=�O�<9H*�4�}�A�u�ʳ���jQ�]j�h�eWW1jG��)�%�d��T5r	�H.�0yx��5�
}R�޽��~�ʃ*��
;v��b��^�V�V7L��;��v��D�.�Ї(��`�Q�VfՀ.���J���w� ��"|;���"TX��F �D���������C��JJa8�R�|Ebn�4!�	o��"��L����˨��;���cl-� ���F��[^�:k��Xr"]i'��1k������*(ſ�Mo=g�Yܗ�N�p'�d�_�V1�a�]��L�5�O8k������jX�1#��^��D�`���<B�މ#�o�$�`��+��On���f��nv��V�onԭ�.uL���d����U��ߊ���"�<w�^��$VįA�0��>��0��j�W�C��qk	��n�gB~�`�W���\�L ��z�Ti�O�3	H��fX�8�2!��_�S_��u�S�Ǥ5�|}=���������/����/v�]������o������>����.l�na8l��2K��%haL��_���2���y�ØJ�����4����j����E��� ts٨$����I�`�dtPr�=�U�0 �}�V�tk��=�˚������scRV"&��2�Ο��,���
TZ�H� �S�mBޟ�	Q��*�@?V�Hu *P����P�4�S�.���������x���r�8P➅6y���)8l��X�^d|�hmI�.�B&�q<!��#p��S�o'a �cB8B9K �@�Ȓ+w�ș$OX�Gмe�шe�`ZI��i����mC�(ja���VTa�EY����=�o�Z>I�)h!��uR��@������ś�cr�,\l}����9E��V`��T��H�A2"B��d)�V�!��P)B*K�������7E����`���4����d&D�������*N1��,D��#��,��m��7|�E�C׭O�9lP����Ђj�j��~�b�K���U����;Ok��L�_�٬�E�����E� C׈�1qN夡��-��fn���8W�1r���[~	09r��A��Ʈc򊛇p�r���E�amT�p���Yy4oq���ͼ?Z���v�/���Ҫ�7VM�7�V������0��	�5��O��.B���*m��۞��v�&�5�� ��V�?����cm؇�&i��ۦaj��������rl���!'ff�$�Y+i��`�8��W�.�����~O�\ݳZ�[ڝk�ٙ{��o?}m��;[�_�h��4���=�"�����\~�q;"�e��#M�a�S�!�hx�喿�(<�z3��.��K�#^Ϛ�u@�a�G�2k��ųN��{xǚ��/�?o����m�y��է
;���ݧ���wk��7Ɋ�]ɒ��/>Zv�]���`�*l{@�k�5E��m�ȅ	mDC&��4�	�Txg�te>Y_��+��+!�����<��-J�9s4�lK9���m�O���:��A<�7�󊐏����) !���O"�2��x&(c����V,�e��*�IZ��ϲ��~=�®�+2���k�����|�R�5��Mn��&2X@�R�	 F�Jf�*Q��EX�@��
�)B��
׏Z�1�DW M�J��R�Z�ŝ!��K�JG�oR�y��zǹ+;�]��q�N��[�3��x�64���"���8���LuD&�*��&�C�����g�R8h2	�d �,A�X���)�&���EX3"�*����U����aRz���p|��?#�o! Mr�7��v�%�!t�1�0$�b�đo����)ƂL]~���JD�tٽ���W���Ղ��{��G����I�t�A�}�D��g1���B UdM♲Q7T��Rw��s3�E6|ΐ�I]XX2C 7!r#~s�J�R��j�j�Y������\�Ѫ�ڿ�k}8����Z[�H�"`.�~Mp�MO=Jg���*'�u��� �!�nU"48���T���넗�����ɣ���|�X��xz8�ޥǯò�Q4aY� 2�
,3�6S7c�ϼ��W��z�澛�}^Ǐ]b��W�<�eW,]qe��>v=�R0$XvVAn�=+���������i\.�E'Ә�9<:[�,�h*��i+ξMP��8��g��y�R,w����T��=W>ˌ�a{�f�]�"(�4a"0_	�pcbS���Id�D��e�l�Rk�:���ϐ�!
d�*�嘤�\x4I�T0�,�'k9�Vȵ��xrs�W��
$��"�EH�G��� �#O����,�A��|2j�Z������N��r�V�E��YǞ]w�j�(M�/��/rbr��6b�ƿ%B|h��?��QS�J�Ś<�ҍXJ�ƂlT�+�dht�2i�@�*@R�b2�Yw�̺�>8�ί?|��à�lAEB�y"sЏ��8�*:[�,x�K�%3UQq�X��W�re|y�H�-Vf�ނ,�o���	���(_E���߉���-B�jV�摚�����h��^�eZ���V�J+E�$�#[���dh�24%PWҕv��
0�\%^{f�K ����� ��e�l�#Kb�-�!��?��3d�@��E��舁+3�d��J�HiS�5:TjS��*�JkM�8�ݦ��{ӛ��f[4iG$����:�c�n����=��3���n���)�����?���?��K���&$D���+�k����@�w	4v���S�9���h�ByMfI���D�-UV���<u��\�8I��~-*�vNn j�A�և�Į��ᨰ�,ۉ�qY�r&��JuFŲ=c
41ɹG�\�GaK��X[w�p�n������%�#��ϲ�y���ċ#��|'+[��Q�]O1�?>v��)�+���r斚
:7Sn�=�BL���,�t�;Y��Ub1<��D���$��)/����\KeG�$�BWç�w=��]	�f��&�o�՟*�*������'�dF*��OT=���g�����,���c��}7��Չš��E���d�Yl���[i�G5���N�~9�m��ܛ��*7I�B��@"!_^3 	��8������"��5���'�y�����l���70uZ��T��A]`;�+K$�*�xh:G�ʒ�1��Y"��Ɂ*�@���2:�Ĕ�r�i<aA
�ϝ ��TD(#&�pQ%U��Z�B'T�뒂%*+!'���f�ռe~7|��)�<R�L��
$n�/?��Bo�W~-[j�0%#38"�;w�w�����p�U�V���Q#Wnf)̹*;E�;�>Y�ßQTy`J�%�RX�J'��
�N��PQ@���R[��
�j� E�$K<^T���8Rh�u��.T�J�T�PJLj5Wj�%�a��R��I&m�%m��E�\]{k���~Z���껛o&}�Y���
�gPq�Ɵ�W�)B|u{�ALEbS�7�b>Tj�Xk�L��+3�$:��ۘ@� E���T2����+w�f�9�rF�F�f�<i����}�y��Lأ�i�N���s�٬��Pnr:����C���y�d�~��(2��d�-;|٢<��3O�1tX�	�W{2}���{�>JRd��(E��w���h�iG���p����v�]�a�JD(��P�[�.S8K�rS��1��U)tTr�x�7|����n]	��t��ѧQϲ%�?>�8r�^ߏt��{��G�/<��/�*2��'DT���,B�jJF�+N?�&�+�v�+{n�_��,8|�E�z��8���=�R.>z���xE)���#:�����o��;(&�"��я/_,5x��l<���7�Z]��)@�r�L�#AA��"Y� ��J38����It$�&���%REɹ8�D�&1%�\9!�l��*V�%�^dt)JL��O;�7"�� P󮩩=�S�y���
�����د"�Z�Aህ�$ef~��r%J�_��w���k�	�@�8�����B��7rUx�HQ��\���U���C�' �C�; jr�V����4�=W� �Ep�%Z��%w��6�V�[P���
=���y��:�c�|8�bH��H��H;I�S�ٚXSD��o�o}}9ٖc�D��P����U�DhE��B�x�6�'ӹ�n�A(7�!��R_;:��"��Bވ6m��Sb�L�0�����v�'�9���;њ�W��z�����(?q�҈81��<��v��[����9�<���֦��,QOU��}�wf������⢑KEs]i���G���Ϗ�|�u���ï�m�5b�-f>�ՙ"�d���R�; ]��B\h-E0��Y�ǱN��{�Z�m�`���/bV�|7������c�|_<J��>��̛3A�u��%Bo��
���?G���~��΅��tb BU>��7���q�Ǘ_'�O:Ʊ/�N~��cZ� ���+o�$n�o,��jU�6~% \�F# 3�F��߉Pav� !Bb}>��"$�U�с-<�D���Z=C�e*�t�*W��J��L�XNʳy�l�4��d2D�a*C�����s��4~J.?����$Oe���jJ�t���!_��kA|X1}����3sA���U�*¯�RS��t�B�b 5�Z$����j2������#D�=�굦�}�6 ��0�F:b�p�!13D6��`��"d�u\Dˑ����ZQ�J.S��V:��R�]���PҮpҮ�*�I$�I%�� mO'mK��%����=X�	�a���)j�ީKz�j��i����"�[�F<m?1��P�q����]��Z1�@$r�J�D�zE�V�a�s7����z%e��o�e�'�J{�9� R����ɋ�^���M,�)�<�HY$D�L�ҵ'�,��.�bT6������/�Dv���&�d��VL�eyػTѠ����o���v��r����$�S��������Y����{kԊ��ο�f[�UE���Z����(��y
�����O�ʔd��&l:1m�O�E;�]z��a�"�Q2���]q��bЙ׹�B��ň��Fq�R� ��"$���u�CU���j�f��E�G{Ո�r�ˣA�-D`���H5Ԑ͓Sĺx�Db/K⨄�r���l���͗��N`����u+e���`^�'DXӂ�!FT�"�{�?'�S��Z܂���!U1dxGEP�XJ�)|4�+�aI����Xp!�/�&J��p`�&J�����N&_F���ib��-��d2� G����!��H��O剟	���2�应,���������?��}���^V��p�7�3��5�{AA���`N���=�+���zO���&��PK�g :��#1�+nD�^�=O��E(���&D�I�t�-�� b@���n���׼�vg��+0���	��M�fF��9���ڑ����ֆ�&^n0�_�D��y{G�>�-�5���o«	�T�e�&�r���W������G��|"*{^1�#��h��"K�l���eҥt����8Z,]���=�8�E�!AX�#�|�E�������%3�\}����'��F��3�� P�R)��;Oo��~׹�BX2Wt��Cs��%����$�Ќ�v���p�n����4y<mG[�8�\��p�}؊S�R,�V\���/l]@��k!�zl��s�)�^w�g[_�ףY�|l���x*;�|�����b�'�F$}���1h)={A�+�H6��u��z�3�t P�
�No�
%R"AUj�R���l�D&'-+� +") ;`Gh�q�"��� w�7��<АiLO�7�%�w�D�A�{>#�2%�Xk�+���8S�������#> H�*PG��j�R%�/.ėq�c�hM��_,�Ŏx�Q��B�V��"xj=W�c+���.�( ���Ċ\��ʓR�
!s�,�t��@2h�:ߋ"�,���g�l�$�'�IsE�ׅr!���N�z�kt�:$ ��T�z���Y~5��3U���@��jt����ӳs�� ��_E�����?!�{ޠЛ�����UC�SEUo���ij�Yl��ѳ#�C/ޗU"�V(Use�8�e���-�|h�'雝q���?����2j�M'mM��)���vE�:;�|T0�T��d�O���Q�����I�_�#��P�X����B2�.��RT!�E1�͡Q�T=G(�֚S��!����K|�Yr�/��:��V��%��w�	L�b5K��
x�,f���eg�xrH��Ct���GBb)��`ʜ�_��,��hK���&�܂/��� �7>��LL�x'J#��^���2�#W�/?Ȝp���P�^��Muv^z�#�����k��^>H��i�E�m���]z�����hz�Y[=�������=�����Sw^�&u50����@�� ���<�<��Vo���&�R���Ć�s��DB���H$`G�� K:���<�@�8�C�E���\��C�+����F�)A�t6�%q)?_��Η�����E��S7���څ�A_#"��_5r�� B����fA�a��Dh����v��
!_c�Q�yJW��`I���b%M(�s9���̒d�E�A&��	[��cLZT9��R�/�Bt��BCB��A��e������5ɗ*��t�f��]y%_E���E�%¿������ɻ_�d�%�.��?��Έ�Oh���$ ,�eZ&����y��o7F��K&�J�s ���}�#�Κ7�7�v(x'ID5��0��Xg+��=�F��\�s��;�_��	���&���7���+���K�a�έ{��ȈGE\Tȗ��rD�	� E��
g������wBS[���tym�t�9!����U�s^�m��^�pc%�R'�VImr�U/��-��1!�3|�}G���+��#�hW���]t)���{���q�F�B�U�tJ��`-��I��eG6\
�}�팋Qɟ0
�]a��?��H������3n��t���0I�H���R�{��1���/Ӷ܉yB�>͵����F��g�Mt nDo�`.,�{
����1�C)��v��'�Hd *S��\>l33��nݺ}Æ˗/_�dɢ��,Zt�����4�L�j�/ )B4	v" �������k׮��L�L"���\%WT�Q�~�Z�U�4:[�F���et2�^b�R�Ef�WC���*�F5X�j+Q�:��F�� ��!ܡJ=Di X�#S)U�b9S����劉-H���Y�/�?ƤD�e��8��@L�hB`��LDƒ� �����S�z���˂�5�� �T૚|����A�P�߭G��)�?���5�f�}����/%���@��QT��aU��!b�H,l�b�<�]ֽ�q[r��i�w�4�����7?�|�b׻ֻ޷��y������Y�x5&.�X��2;��BkPȹ
�W�Π��j~qaU��łZ�Q#S�/��[��h�&�0Z�\����y�~�f��+��[T��au�p -Ǟ��S���D5	M"�f�"x�w��?b㱎�%=�[{?G�=b,�?���0]��3V?��E�1�-��(��\�aG���t~2�i/.+�Z�����D,A D&�}�Ԣ��z��luK��T�|����K!��]����c?����)��a!6lȁ�oT�}v�Н������N S����2|���0�g��(^!Fw`�"<�)ٌь%���6*���uUq��
s@�C���K���,�<�����S�Oegd��*"a�FG�<xp���k׮.X�`޼y��e_�̙3G�q�ƍ������O��/;z���Wr���������*T�S����$ZTZ�^��q�J�WiJ`��z���g�4Db2
�:�h��lR��j�Z�1�F�7��"�i�v�G� DU�:����(lQ.[DeV�0�-�b	�������`�%�
���!��	�!�>x©����&D�������k���	�����ߊ�&"���4\�l�����2��*G(b��9zJZVjz6��M�Ƞ��b5�C���C}bs.�.P�)�؆��Z�;�|�~[�	��n��&}�"}�,��0�a�S�эSW����$�b�!Okp����b	 �~�֨љ�:���Q��$r���Tz5�A\�J�`��>C�������������D��`q��>�x��H���0}d�	C<�ŰM�����s�ﮋj�BH�P�]馃t���MW��&׭?]3���k}M��kWn���*�x�l�{kvo޺gOf�SX�ʶ�ޗ��o&O���s(�&����J����2��R�x�X5*�t:�Á����Kg��}uaYr��J��G�{�u����_8� �6�G��~�k׳�S��ǯ?ary)�A�!�N�\8}��l�g8�<�Nj�B7X��3�,U��cu*5;&#�&����K�ȣ���w������X�"��O�5{ڬ勗v����e�ˋJf��Ç-X �[�j��9S&M1l��C`;z�p`�葓&��<q<l6��Y�߷wO8ؼY���)eHEI�T�ݨ��HE@lHPnz2�y6�:7+�Ϡ��R�V/�q#^y�6���S�jS�a�հ�7��1�e�j�j����U��%8l��� ��z_�M>N��<IX�S}��6ѕ�A�B��B ��:���<	[����+V����M�H@(���	��!AM��Y~5��3ğY��*ub�����U�����D���0���%J��Aeʔ����O�o۱���+V�]�n݆.A?1!l��F�������+�/.�!1���P�)]��r�y�1g{,x1jӻWԢUa���U�DJ�v�tyrCl��D��]����\z��&;Ƨ3j�P꫆�C����i4F-|
��ʊ�ee��e�RD��0W�pQ������aQ��4o?��"dh����G�i;l����~m>ݧ�cG�g���[\�F^�n��U�����^�or� ��Za�����%_��/7),�[4j߻˄y3�v�4s�l��l��!���_�Z�{�t6-�e�""��Ρe�BH@/,��x��<�J��;<z�۞_���"���U��s>y�)�GϿ�,�sa)�XZ1v����J�+��߭��wZ���~�)�ۉ��{�5�B�I��ٱ2geEIye�g��J#�C͡e��D<�x��e&��(�p_�}��9_�@ZX\>{��63d��Y�F�S�&�.,�7�8i��	�Ǝ;f��aC<���A` #���O;j��1@�N����֫�/3�N�2al��=Z��x���%� B�R���I���%�3S9�,	�����<8ǤVڵ:N6�ݣ@��f�Z��o2��&�݁z����^���[n�!��'�HA��US�yD X��!����!�N�p�.�B��s!WLt�.�-ȓr(O(�"l�)=���ߋ���B�D]� B�R���U�_�ߔ�?�w|��=!%���S�ڴkסc�N����3hА>}����g@߁�Vox����LO���E(i>����\�	<����n��@1�	K��`�ez2����k��\�0`AT�_-B<Ŷ.���L�2���B�Q�]xf���n_"B�VDldaYX����㶖��+K<2>�KI����E?H��sqÛ[GmbFe�3,34��T�thE�Զi�>�{L��vݛ��y$_�7�=un�׽����n���y��5��4����f~�Ǖߞ�<��u������0r�����4��f��|x��l��]���I����~|y3�/*�ã�7��Ơ �E����)(q��^�}]��V`XBZƛ��aq)�ܿ���囯��:�z�ٝgo�:pa���1K�l<uMYA��g_��^�;s�Ԧ���ٰ~E�QS� 3�]UZ�x�\�+?����K�[�fgz��Q�a�G�޼r������ �)uZB��)���Ϳ���4�_�у��cԀ��j>uܸ�ӧM7v��a���ԯ��A�GP�ȡ�FRS�C�n����۵��K�QC�9^��*T�S�N�)��똰 ��k!��
�ѡ������������������,���&��b��l"����	����ƻ:���F|�ׅn��C�DO��A�]}	�Kwh��R#>�,��Z�*�6}��Q��r�2�7"�Cb4�we��!�OL��� l>M�@�
�
�H	��X�~/Bp�����N�*�T�]�;���K��|������j����<�\P��	
=~�/�z�߸���G
E p�|9�LIL��sa�ҕ}{��9뛕��f#��R��+�BM��Rj�I�9
K`6�̫�o��d��l�R�����v�e.j*����cA/�K �B��\d�̷`\+ό���C�� �t�9���{'w��*��z��b,./��ٰʢ�"w����I���
�^}|��E�F�}s><��MY��P�:7�u�Z�5�����o�ޛ�=��/�ooԺ�u�Y;�Y���������|�i��iab�L�⑧�A��Oj�XLjҖԬU���H$�/;�^:W��ڹc�D�)+pI��������������-�M[\����ܔ���T�JUB�|�����g�3W"x���S>g��z٭{o?��i�V�+��>�|����|[x�V�����-��=����W|��=����s�[�y��)Vj� �Syq٧R�C��Q�̴��K-X�Y����ݽp<���O�*.�1P�?�2�8iq=��Ԧq�	Cujռ��m~�qĀ~[V�?bĸ������B�cG�0f$��2nd��u��{w��q�_ڶh�m����*+�aJBl\T8 ;��({�������\z.9%99*"1&���;4��"�>������_���&�n4�UIQ"��
Gh��)

�g�
$�B/� b�C�U�q)~!��@J��W�U��� ��E�"�ᗦ症�x���3W�x�#����k갦����R����K�5��^p��E�4����|��L�C�\1*@��*8<�u�N�
��	D X/|@���� ?y�|т�;w��t��˃�U	"z-(�2���SԮ9�&�8;�/�^@����V���Ӹ!�#�'R:�*'���:j
�vLU��G�&��G 0�	J$A�lp�������1�!��cx�۠�\Z�N+�!��O�#,r����&Vab�<	8� ���[�Wd���;���Y�����ߡW�����hvZ[碅�g�$?{-?�7��|m�\�u/ۀz~���Ά�.؇s�����^��u"��}
�fߵ�"lڰ�ը-p;����аO%��ܽvه����s��a�[��s�PL��1I&��D�9����s~���XiV�{��mȋ\f�#[w�^��^��ڿ��ٽ��-}��������R��f]|Џ��N]�{q���-��l^�t�k�>��\������X�	+��y�����0��,gc�Ni\��k�������;��\�i�/�ɑN�xT�.�7�3~L�N�t�2��c�̞4q�ȑ�7t��aC@����89�0f����A�7a�Љ��s�Oԧ;����?6�_����n�r�SY�ӪW+�zMVFJ|ldzZ�ͫ�F|l(	��� r�\��U'��27}}���!��g�G�{���A��ndO�L�R�ɋ0y�<��,�,��)ˍ�0��0,�+�IlŨ���
�<x��V���M�f�;��y� ��X~s���|����:B���/�RU%G���-�B�� 6���F�B	1�
�ą��"� 5E�AU�o .�6���O:$ �g��f��H�3�a�/������"�G�"�׃e ةn'�<�4�Y"y\�}x�H�������HBJ��	��̘�KgHdr� _(zKM�9B����|��5MM���/�6�D+FMb9�Q���Ӻ�9�˂SKN���W���ȆL���|�U ����DeG�6<���	j�v��-�gI��s�=7��qѵ�]��n�cB�h����n`��Z�C�V���ӣ'߽{����Q!�o�'G��F��VjɊ{|���׷��<�)5�Y�ӐɌ��}�WLv҈U��	�r���V'� DH�$�������Z��%s�K��%�w�m�����kx�+�{]�X��y4X�s�~�AXcҩ�lX���m�V�a�ܸr!%1<;#����.����ҙ]Kό�1SF659.5<�����C�P�]{p!��=�0���v�:w������Zyh��#��?�u��ճ���.uT��#����s�}�>�|����[��|�&L䁈P�.y���B�pIp����O�(5<�!"� #V��顯�\y����󛙉a.��c���;��U'�ݱu��:wԽ�����9g�ةcFO>b�� ��/E8n�`���e�6?���q��m~��Ѫ_k2��\*��2�:�9���}N�\6sjb�Ƿ�<�ˤ1s�L:����G��Β�ڽ9�������	\~�3�6w���{9{�e-8|;������ԭ�g�\xǵclk�����o;�,�$�2��Dj�]�ڽ.�y3q{A�5a�(B�?!aA.��"�ͅ _�Sc��7�TÖ� b�7��ׂ
��u�~��|�?*�s'��̿!P���K֤�	��5��&������\�@,��ټ�{,X�(�H�l.�P�HD�"�	J�R�P��e�QmF:eӦ݉�Yb�J.�K�r@,�C�U�q����Ȫ��6���r��ÏQ�c��'���+qq�����92�@�	�Z<��Lԑ+��e��=h��Q�]�mv�7��ΩP9���b�O(���E����jW��Y�z���7�]0oFX軬��g��(~y�##%��գrD\�szz8����Qف��ŉ}~/.w]T�����F��'y㼚"�]x�L�h�u�@��u�"B!�jP���s�d�=�� ꋸl��D\�s��I�&��w�����v����w���{��Z�*����p�\d���p��ˠ&*�����[q�O`�è�k�/]�}ن�v��v��İ��V�]��Թ�'ΞQ�4�b���<'�nۮ�����u���U���x�s��{]n/|�ƪ�)�/�;�w[|�+��	 B�Mf5IR�C^<�s������Wn��ߪS�i����BP1��f3�/ڻ����@��Ə�2z��a����A!� tX-B��c��DPر]���h�� ?�Sy1�F�w�v���~�[�n:w����gc�3SR޾|���Ӕ�xxI#�P)YR��adԨ�W�&�}vozw����'w�y��!���73�d��at'�&M�:�
P�/2D������|��3���*��2��D�(�]���pa5�"�Q諂B���P�X�I�%�#Ļa�[O �S:�b�4"�{G���Pf�*����U�������� �9D�h�]�Bi�������"�K9)-�Y�ᑨB��Z���x�T�P��"paVf."VDD&?vV���
$�T(�J+D{��q��ݪ�?.��mŻ�X�Oqũ�|!����{��xa~2��Q��%D�RTz�X�ǒ��%�iQ��Gn<~w�����g7ޗ�t�ۡG>Dh�u�D�B�Pe���<�u�֕+��3��e�""B�%'�Š�SS����ۻg��Y�ǌ3bİ�~��zS�94�*�"X�㴺��H�0��*�k��V�W
HW�HW\��խO����U]xq�,S&M��Y�aCth�b����fNرs���s<��ʊ�	���z.3=9=�٫�GO�z�Ѯ?08Յ��oß�z���Ήs�N�;iƢ9[��\�fɒu�.\�����Ǐ�:z���3x��3������V͞1i�ҙk��<d����3�6_J�>x������fM�vɜi�{��BZ���Q�h���o\�qa���Ǎk�}P����MZ�d��d� ɢ�"���2ߵa��}{�<`��a3Ǎ�<j$�CN?jƤ�𥎭�w��J*�~.+.�w����۷ݰn�ԩ����{�����޽}+)66+-�΄�(0bLDxvN�X.>���ē�o��n�=y���F̽�f��SI�'&,�86��$.�U3j���7�2�����&�V�x$taBG��Y���Q�����"pz�G�TM̭!�/��D�o���u��#B��'����"�G�z&��2LD���c�~�!�C���y���'T����j��	 I�����[����z3��S�Q�B&�K$2�EB�P �O��a��E�ٌ#�qr�2_)��@�rDne�yTiY��g�nz�d���{^��c�n�)'o���Fk_�^T]���ܧ\LR��U�6�������' E�rl�cZ���H��v��鹁��{5��GZ~����+B;�)T@^\��_�7qB�����{��u���������������7o����_�8�svϱ͉9�0�æ��iyQ���E�:p^� �sA�J��̵|M��@����!�\u.��O^x-N�s����WVV�\�3���Μ9u��~�W.ڲ}}hDPJFBjv�ǈ'2>�ޓ�붭oѡ����c��ܻ��+H+�
��N˹p�?,>�����6mظw�Ǹ����D�������Z�¸�D U�8�w�Ё=��_�x��Mۧ��̲N�xAd�dς��:�����O�����%r��I��Pcȹ1ٴ�zܺ�[�S�
�Ǳ����jo��³@)�K�C��2z`�	CqN5d�a�" X� !�	��N7r���#���ұMǶ��?~PYQR\��T^�����{�w�С/^�?>,,�֍kϞ<�IMN|��޺5� �^�~��l�}�~�w3�+��=�s�ډ��ӻ��s(M�`4h��؃TS����KT`�6��q%y슫s�>�3�ؽ���I����$v���F�n��j�L�g���( �"$�d_ƕ��	�*� ��*-h��^Hd����;��]�aæ-[�;������L��x<A6�
MR�A�b9_ ��+B��{�#j��
B�`A��������R$�FL�'XS�����S\\^%��#>�*�T��D�;��P $N���?�����"LϦ08��K��|#I�*�F�S(T���@��Z����RX���d$&˹\5�K�P,R��Ȃ��e�[�4Z{g���YEX�[� �ǝ��&���ISo�x04 B �s�
�¨���uei�Q�ʀ�n���^x�uH;�H�H{RH�����ۡ��2<[�@�(����Ow�޵i�f_ߠ��"� ~:(*/d�Б��O��&�(꾣��(�e�[�a}|�Z��|u�/Y ĩ)B?��"�v!���������U��Q��Z{o�����|�V�	DH�iӦAz�ڕ���Cps���~�cRb�?�.�f1r#��,_��ؑM��[��Ex�͗/�1,��g���E��LN*�	���GO/޸y��+�J-����<�ͥ��-yE�e{ϐe&��w�_�y����������t��m���R&����{���{���,r�GZr(�G%�&$��{���z���2��H�������#iLke!����XP�g�����8| n���'��o�p���'�ܿ�������9��KA�ٙ�ׯ_}����˗��=~�8JXXxhpJRBZJRl4Ĵo�����ؔ�i�q����@.]8�4��y���{�>�̇��Cnfٟ�J��x+�:��/���-�7�|�h|�l~���B��Dd+������U�Tj�P|����K�6j��u��ؾs������8hА�S�_�x���3l�`VY�H�_��ڂ�"$jb�����2_E���,\DTM���E��B|[�a��
�K_(�_-B��!5�~Nf�P�t̸	\� ��:�H�b�\X�Rٯ��~�2�ل"�rE:��2FP4xݍ��.�����\�E�[I��6<oz4��1����z+_}3���C����:O�¤v<�L,Z�^X9|��fs/ՙy�Ɇ�:��H[�H��m����?�>,N�'ДH�n��	"$j"�֌'��er�Fg��mZ�Z�@!���,�	E�RA�!oL|侣[�(��"���~��Կ���}���p�q��!����"���k��g%�Jq�C���Z����$��ȝW0a��1�ǽz�:>)1���E�d�xZ�E�S�&E�����b�M�W 2;�V7SkN�J��a�5/��~�1�Й+>w�l��{�n\f���De�i�N��[��[}�Ȕ�642(�cR\��W/��\^�� (m�Sr+&U�j4�z��К�}��>�U8�F�dj�-EZ��jL�2[h���N_s�R앮�r��*eeǵiRw���N1t8q$(p �,T� �F'�.ԯg��-�����@�VQV^��'O�D�D��'Rit��Ri�:=`1��6���r9f#�јg.��y�M�r�R��;g�o�z�V�^�1 N��r����W�i&,Y[�����&J�,�'M9�����bG��^ �
mN�� \X>�K��xB�Z����mشf�F���I)��cr�4->>���'�V��ֹˬ�3>�"0"���ݨ�Q���'B��G��&����3���"�Z~+�y�UD�?��A\� q��A��߬7|W���đjVSmA�D�I,ބI��`A�ވ��T��R��P��њ��\NtT���l�\,� J�XO;��j��v���ַMV�|�qz1f���H�n��f��H��>�6�tJ�շ�^��0��B���,ˌ���K��U�2�my��܋�W<h�>ꛍY�-L�5�߮����+�A"����XaVh��7Z�Cg���.�֛ͥ��0B1T7J��l6�4:|� �B.��x���d�FCg��=�%5'�"��XﳱM��!"�u�L�h�7E���`��}M����~{���υť B�'��&L
�d񹱉	�/�Th	�I-橿�������r���*��s76^����u��#u|J�Ko<�w�o��y�Wlٰ�P�����D9,n&l�ȵ&�3۱����iT�AOOMy��ف#',ۘ�T,Y{���Pm9Od5�
1��L�1+���b���J�\兎O.7�o���6sb�ϵL^vl�ҝ�9Y�R��H�R3���~G"��w�������E8vԐ��۽c��}�h��ʊ��Sii1�J|�&%--95�!���Z�B1[@~�^k �jT&�./q,<y�V���{��_\>qnݚ��cY�_��:�eÉ	����,ǧ(�����J1��P��/uy�b���e^�
�����c�W�R�@U�L2mϾ.]&Sl� �1_$��d.�+�<޽;w�M�:e���p� �(� B���Z �"B�kT(�]�{��Q�
���#N�#js�i��M�'�)�*��*�_E���V�]r�޾��#ְ�=K�%���/(ֱ���K@�ڂDC���s�������F�D�Kc-]���7X ��Dą ��BT����pa�'�L72"��L:_"3�6��X��.�H�lx�t�o�<�aۇf����4Ɓ�:���3ꭼ��@L�Mj/��z��S1�H�+�hn�y�3\�E��<�\�q1�v�m��W]V\�7����������#m̪�*���'�7=��e&�'��%���\3Z�BmÇ*���gSh,J#�F�h�Lf�Ɋ�������d2D
�����kx����@:o ] �U�������CS�ˆo�� �"B!º���I=v�
bZ�?�PXZ�)*rx�3f���
��J�2�":*��,l�v��_c���3�1�u��T��#���9�6�Ѓ��'K`���:�Ƕ=l׽Q�w����ў,�)�eC �ʔ��������KQ���iBQ�
��U�SX�)�E3��b"M9S�bJm4�1�/O�JrQ-bs���"��g����,�-�n����KvGe�XK�*5��@�4�g�1C�����������e��1#����֡�ύ�ۻ{{eEYIIQII	�B	���LI���Ρ3�C�TW,�-xv�A!�֢�ڲ��6�;�($���"�U�T6=ja+9*Y����r�����K�y2�K�v*�v���V�ݪ��֮�ڕ�j~!AMB��?HU��%
��p���7�ރנe�D>M ���l��e1	�S����;}�Ԍt"A�b%
.Bo[��GH���x�7.�m=d���$D�J|�U�4�F��T�Hc�b����l � ��$��9=p�~�)k��2�Vg~�'���'�����k����E�c��,03�F��@G�Ht4��.2�^�.B|�@C�b����!���2��ЫCB��k�P�1dfQ6oݦP�F+`1���Z� z�B5�Di�	޻�(��Ρ��c�
8V,A��z9��G��>&-zR��������fq��w;�ኻ�D���Y����C�4b�
,Ό]L����o6�Ⱓ!{C5OX��blv#��^�oHk�I��I;��l�i��yۅ��Dq�Cf,@t.<��Y-B�Z/�ZP�Ci-�9
-��jW���E!���xS �J�ښ�Y�٥���ޤ4='ltY_뜡���a�-�ˆj����$�|�w�q�:�%mO�/�J�����"�;��#�M|�[HLB2�NE�a�B�s��Mo�7{M�\����u���$�īdm%&�|��m��_?ci�c�O���Ű���J>3x�\�.(��	�� h��MV��������r�<v��j�W�Dj��c
�-�<�à5#tT4�;G�eX,��f2f˭�b�ҭWo>��W`�X�ݣ��Nh܀ԫK�у� ^�"�\دw׶m�7nT�j�/X0��S\\�RHHHz.B��(B�D�֘������E��q�
g���t�m�Q�0�5f���7xS��T�Z��XP�C�k�V��h�V���mv%���N����+Bpޟ-�Q��)���ҧ/_?|�^��E(�A�l&�Š�X�����8�s�J��Gq#(\�x�O��7"�Z��X�һ���z��!@]<���t����jZ�jOkr�n�6�F���Uظr�wb��*��F�5E���[ye����r�����k���Dh`���M�ZiR35���Ul�
-T���]"�\��*�P=M��	Թ�*�k�JU錙dڭ{��l��b��	�9��z�N��_:H�3Ѐ���!"��tU,VQ�R�yr��|�P �}��K�|��sҒg����E�\w�sNd6�6D��@H�`� 9���2��	��'BZ���l����o���/��n��ï�c߅e`se���֞0�ި:�Cny�f���}�i��^�u��A
A�_&Z���� ���r<��msB��\$���D��Y^��|��G[�_�|wNY��"�[��7�!����P`mP��H�D����9���/���m��.���*)3�=�G�6~򻰨,��cLJ�$$h�\�"�(?c3����J�b��,�6_V`{^��}m���'X1��.�+���ܼ�8Ăk��B����ҳ���ǗB��T��f���19���CT-W�Q�
1�ev�ҬRk�~�6,(C�(I������QH>����\/�f3��*~^>��*m9�s���K�_��"��'{��hC�̌�~��{�>�����#1~�Bx๚�#vF��=rp�^]Z���I��1�.���qe���A�����d���%�_��X�Qc�>�i�yjs�@�'+�$+(W���,*|)Eh�u&��.�;Q�Gi�S�
�|�9Oo�7�� ����n�i+�\o?����/4+��?�%����O���7����v���/E����X<���-�e��_�6r�A牠*�O��B���7OI@�l�R�L����r���P�Y
3[n��=\�Z�l������F�W�������yZ'KW��1��L���rx���"��A�䊾��k���Q��Z���"԰��8���J�����P&�ܔ#1�����"�@�ΐ��\Dϒ�QC�ܔ%�R��\�T�*�L���_!���b���B�'����G�@��py,6���֠р�v71���S"$���k7�A�w K�Gw`�*l���_�[HZ����\��W�������31ay��;t�܀N{?�?��˭�b��F�,���o7[���������{�x��;��<��b�_����{j�f��8���G?��a���3��	��Ԙ���d�\c��E��Qy
[��!��!�nP�Xw>�k��B���0sQ-T.��Ύ��9�X���v��Έ���������Y�?�� )�H
��0���端u
!�H�s*n�ݤ�O���?�K��E�'L=y��D*O����D�%�,�.���1lѱ�W"rCE�wS�cv<L�b�o'
0l����
�����/��;�8��ޣg��9t����M���y�����7C�v�A/���)��)1���ɩ����I��mZ�X��Yr��Ǟt�}p��[m��}���8Q�{�"���\�+f�=�4����xw6߼x��%��d0Ee�'�S'�r��]{t�0�W�����|�ÿ���!��1Ca�1r0xH�^�q6m֐�g�Va~a���Y�2|�*-4k��:�L�@4N�ѓ�j9Fbs(,��d���v�+V�&�Üj�G4��M��\�L8�#p���!P-B��VͿ�D��� B
�+!"拄��\�#$b)"�r��+p�\&��`��LS�J(��qc��z��V%,���a_���鈒���RU�!ˋs���<��IQ9������(���`��\��Zxz�b>K]����������/�՗���L���Ѹ����Ђ��R�&���V\�?%�*¯�"��IM�m��5E�ɾ�	!u���:��8uf���B-�^�$�DP�YI�ؑ)2g����e+�Y��6�\�.+Lx2ئ\��)R�YB
���ͪ�H���!�2#�gP�B�P���γ;;�F�^�T�P%>�EQ�q��x[��jB<(�?����l���}��ֽj��÷�>�ֽ!m	"�j�#�ٺW?ox��N�b���-��z6�K��"lX�u�lx�r�˟66����w�����y��l~�j��	�oE�s�_��c;���c��=��Ɣ��c�C�!�r���Ԍ"ZKa]q�Ҵ-g��{5�b��/es��Hn-�<e륵�o �7���ԜD��|������@�a���H��Z�=���o��@�+�n� b�/"��"p��\�K�:�к'X��Oz9k���Gn<�!(9e���sC��h"U:]�-T3���^Q�� g@��I�'��\����すV|���ˡ3�>>��",���6���CBhL����.^>~��Wn=�n�/]��]HXX���G�S��M��F�<88��ɩ�t�$߸r����en�I�B�/V�i�y�>̱&۱4;v�5e���IZl���7��,�`s&�z>��[�����7���O�yv&��MM?w�t�zu�tl7d@_b�0a�0|��B8T+p�a�Ə=v��G�2dĀ�=:v�ܦn�Z��.��W���q�������H\�i���%�	eTC�I���O���V	>�Â�lB���1 F��b�M�Ic0�VBT�i�N��n�1�dί^U.4���Ux��? ����EQ:#�TK���,1*�ȡI)PT
�]�2�wM~"�� ��f���8�B>x������J�\��O���O��D�M7���P�LF��(�9WU���Dŗߑ=�M�1���J#��wY�8�����TXC(��	LCA<ך��bY���P�g���b�x��{�,��1V��4�r����!���!!BOl��J*>}F�����A�p'%!B6�ޘ�/�M��-�Sx�jܘ��F.޾���QY�S��]LB��J��(4Y��LB���G��L�y�ޛSW���.#6C@��R�5W8@��&�1��Č�WA{ B�����l��P��TB�U*����� �#�dr&��Pd"s|���i�U�uք���5�����6�5���Ǎ��g`��j/{�hc���>^�c����؂7�k�9��[?��R{gi�GҾw�oH{_�v�%�x�����R�s]�������_&t�{x����3m;�)�bBu�T�j��d:�Xk��m��]��J��Jlw�~�V_��2��Z��Ԣs�\�p����Y����O�rl΃��d���VS��8	~{��0����t�J������YF��17�}w\�q������M�2r���ѩ��!5f���X�&K�a�uy,ߕ,�2��C�`X��2Y[��-�c/"���D�̜�dÖ�K]��#�ڝe�׭^����Gaa�G�i�&�Z.eKĴĸN��a�Ps�޼����E�Ue7��j�X�8��{��F�^p�%ؚ�Ћal��9_Ҍ�R, ��h�5��L�r��Z\�n���
�?9�]dFNRj���/���ѱm�>=��2`�����1#k��P �,8f��5h��>����ӿ{��?4kިu��o߻�P�@�f����@��^-BS��	�	�B
��$��:�7If�ɬ2�(&���E�2�����4�F��&����]-B��(B9�~�?�X�"D��� 4.�A�j�B���oa��9���B�w!W�ax,� �N������R����,�!bA���2R�Ý��v�Q��è��7����T�����!���0���cGn'�>���^�L۸����V�`��vu��{F��ߌbZ~l鑛#��<�0����*-Pc@8X-B��7�����,.�,��$�*¯��M�YU����E:��q�Jܠ�?�a�<0v��g�9W���2z��U��)�D��U��M�����7^.?w�;������[!�%��� ��ҡz#�ǃ{��f��}�V�6��V�Y����J%2�
��`A���Ssi�ڧ
h�f(t'�����`ƍF������9i���[����hSpӍ�2�s�<�ZkMH�u�2�c��If�퉤��]�=1�}Q����a��!�#IG?�����v�>��9��.֜�a�"L����د'c�̿6q���ѨH[*�:�Z�\�S,����/;te�G�Ell��h�`:!�71���3O������9�o?95+���v1K�1 ��������^�y-��������
ą_D�o&��H~f���z>��Cn3��y�j����n�:���6��F�<v꫰�4&�U8"3����hπ�[��P�wa��->�l��8	����e'�����U���aH¡�W��f�[|������}���}�q��ݫW��v�VD(.B�Zm�+MZ1�w�܁Ϯ���������;W�M�ŬQhu"�CS�Zv`�V�A�|Fm�4r���$qZ���4��������i�C�fTb[����;��^+����̈�,r����v�ЩC`��A�ǎ?
D�q�H��Ǝ=n��#���H���{t�ݵ]�6�7��T��zݲ���_T�",��Qɹ�1�9�
��d�B�Xa�j��D�3�� H�82�Q��>�C��T'�;jt����!4�����%'PS�
����?!�F�	"B�J����2���Rt��2@�ViT
�R��".#|����!<�e��lNRf抍p*p�Q�"B)� !B�BJר�*SX��À��w�s����,.���h��S:�<�o���'K]�>q���"�4�=s_����m���d)�w^�z+"����ݏ�l�+�B�*\�r-X����9)����S�wF�W~-��*z˿!	"3!�E)U3�L�a����o�2�U]����8t��w7���OX�e����>�"�ϓ�Cf�J�3��H��~�zԯ'}nG�䪨\C �a
 a�������Z�>��v�T�feg�ə�)T*Y,½��­Z%Bh�zc���H6G���(�9U�g/;w����?̽S%�m�I���n�j�)����6�S;�|�)��I6iuL�s���H[3H;2I��I{RI{I��IbH��H�#HG�HGA�!�SI�s�Iigj���|s�10���0q�(�r�ZTh:*��Ku6\�Z�G�D�\v�Z���F�}��`��˯o�JU�����+��	�$��r�����D��RQh���1�JL����^P��WG� �?D�����H?�,H���s^������6�ߐ�nn9��s�P��QT��;�D��9|U_�HW�_�+������2��������^f(>ߋ�|��4�e,������~���8����G�?y���3sf/X�dŝ��@��4h�f-ZQh��PPU�[F��ȳ%���,zq��E،ξͼ�"}ǲ,8|s�Â|L�KW_�����j���4z�k��K��ߌO��TJ�Ĵ����������Ƕj����u��y��aǌ�9D�[��GO5b��#�ԻK���w�k�m����]<���k���JK���d
ĸ�iل�L�@�B�e���ʵ��Z���t�E4�E�-��(�?�w��j�P��u��%*�T��6��j��u�Z �����Og�nBz���Gr܂^��2|� aA!���-�ҕM�I+��F�[y����_��*t!\M���'J�������ŴbW�g�_q0�LW|`����]�ҕ�tt���v�6�0���4M��ʍDQ8��|���2Ԧ�"�Z��R�@o�� �k�9�p���UD%K�9�Y�,�e9�e��"K8Kv#$���5G�Du���f��Ez^�q��2x�bm<Z����Y�.R��,�#��[6����Ybx���!�>��P�2D
|OT��޴Ys{��ӻw�>����{ؐAӧN9rhߛ�/B�?dg�g�g�����%"R��He	��!�,�\)��{��!��,��rS\��q����EýQM��6ۓ��.|�ӾlҊ�������v7��=��{)u�R�ٟ����oe���'��&��œ�Œ�G��E����63H�Y���M6%5Z��ߞ�����N,�c�b�l��^�C�f|y^�Yi�M�ԮeGn�|I�3cq�eZ刍��n,�c˭[�&���0Ud������2R�rV�ð�YZ�5�����f~���2�3��`k�Zq^6�|�85���o|D�ΰKm��=iĶF���0a�[/�=��g�N7|��QS��d���t�6�e�>fٺ#��Pw\^v�a��S���O�q�q�Z��E�Y�ϱ�x�U,]��C؅�w�M�6v��cǏ=f��)�g�߳s߁��/���q�*�ZiѠX��أaRb���@��r����4h�f>� ��P6����4ݧl�g�_�k^�po�f.�s���@M��b��R-5�Q�����-*Ɣ*]jF�%�ˉ�I�s�ƍ�3g���O�[���Y�N�;�Ǎ;z��4`ذ!C��;�O瞿��Ժm�v-:�����:��j޲�ڍˎ�8����s��e�%ŅE BP{ZrFF*���`1\-0p�w��U��j|�^���&��B��4@���E�\�z7�6x���#H~��)��k�w�~��4Zំ�G�P��rT�Q��2&����)B9XF&�I���b��e�8a���߾����.�&�E9�dADW-B�R�4����o:O��iQ���4Ge���0cĖ{����K��˽����\��8G�e��so�s��Su�4��ͬ�O���,M�h7xz\.��QG�V��*P[�N��G�W��R�@oB�V��"b%"7ӹ��i�!{r�Xja$Ֆ"�O���у�l��Zv�ְu'�tw�c7��>I��w��A�e��gӸ`AB� �� DhHt�Єr����(��G�8���Æ���ЯW�mZwhӲ�#����1#G�۳G!��� *7�$j�w�U�d�]{�m?�`�1'���vCH��j�Sg��o����������nK$-|Aaíq�m���1�M@���������z^��Uy���3�_�����_5_r�կ���^xȒ�1,�dej�"x#B�w��M��r�$R�E`w�X�i[�r�ٮ�����<�� r��C'��i��T%G'{.PLF�}$�tJM:��s�\��Z��^�	DX=j�ʂu�K:�y%�GZ�,��qr��A���i��N��x��GQi�ŞWYu���SGL��.*-����㨪^�V��=e�ϼ��R$�vcٱCw�N=�J��i˱c�?���Qzx��D�Ey����@B'O�>q�L��ջ��}߿}���cv�ƦF�<z�I���o��i&E���zx�Aɶ�*�F��0����Oo�}��v��7� �5ǯ@�8q��I+w-?p����G�}���n{1d�V_��jB:����l�3�W��z��]P��];غu뾽�vh��Ǧ?�۶n���νz��߿o���z��չG�]ڃA��oI���C�&�:�\�z��S�;�T�JJ\[QA�B�&�"d3<.B�F@�L<,����ӗh�R��D� �F���� �1X�U"7��*�T
�>��`��=DP�w"���|�qI�T*S��q���
)U%%k�t���r�1�S�V��H��0u�G�������Q�nP���{I#_��̵�hr�����*��.m޾KLc^���b��7��,me���{���)���X��)����DL%�a���`�[����*z�(BO�d�B��#�%���M�p��$6�0�b���_��������7&#y����+��Y�������t���_�&��5d����ϡ��"B�h\i��}&M�9a¸I�FO;lΔqsgN5lp﮿���mP߾������S����j[�Mx���L��*Q�ly!l����v�i��i�;Ҧk�-WHk����.������7\L�u����W��aك���i�ݟ��Z���jكV��h��u�%o�.��u�%o�/�$�Ò�=Vv]|�Ӝ˿�>�y������,�A���xo��B+�"B�ֵ���a�^�������/��?r/S���7aϙ��78��T�w�ќ�T�Ą���������miM(i7�t�������������H̠���L�d$]4�.�H T�Έ�`��D�f_!M8����?N^�s�:�Ʀ�䙋t.��1㇎��:,)��2��������S�dI��}.>��Uc��;t3ʄa�LS���|<Ml����P{���ZavX����?m��E��dR&������r�K�e*T!-!���jԐ[(+���4G+g��:5��*5�~�qߍ7���?s���YR3[_��D��kOO�}}(��ko)|+!���������+)����j��֝;�.�%5�q���۷3r��ac���ߡm���6mԴy��?��s���k԰v�:�:�:`�z?4#6o�C�Fߌ?l������6��b��RZPĠ�F�E�ħf&�P3�,:���7ER�D�'ʁ��g�'�@X�7lR�Cjp)L�$B@e���� ���0�"�����|x����z�X���80��\z�
��cB�~���@"��|���lVZv&�`�j����J�r��B)zM���1C;l�ɇ��T�g��,���7S@�����ۯ$�����O>�7uǬ5h�O��b����m��gyzg��6`��3!�lUI*G=}�V��xo���r_E�U���T9�[�R�\��#V�
�%l�J��&�ȕ��ز3p޲�ɹEi���Q�7�����눑s6g�]��ϓ�Vv�48����Z����u>��� ��� �,��D��ˍ��2j�؉S�L�4{�9GϚ0j¨����گϤ1�&�=rȰ��{���ՂKRRs��B)nA�XC�A�T�IZ��J�v,�`_b��t��ݾ��)GSʏ&��H.>�Z����L��R��B��7�\�U��*��*�EkoDZo��o���ù�7:�^L��x��׃$�rٻ��1ƻa��4m�G�(�6��fB�á���`���c��S�?%��]�0F	���&Oi����$�!_$U��u 51���\2+���g���o�#ͼJZ[�0�'_����}�uN*��hj_��\��:�!�U��(Ig����\҆Ҍ���I#�4����_7��tb�����q�+JFL�2fڜ��T�@MÓ8�'�bˋ�h��0�u���5o��_m�yz�N(�P�h��t���k=�Ƃ����eX�@���L�����ہ/_Qɹ2�49&���
���U�4ߡd&�<��䌈��:�۾D�2���i��IU8�$6�C\�\��A%�b]!!4�e�R��B����f�@1u�ε��Ҳ�Ņ����'S��������I$R�Vmj֢O�~Ç��oȰ�#ܻw�Ν;�hղ�;k��7�׭״A���v��S۟�7��ئ폳�Lʥe��=����<3������"���|�X$�EA$r)Z%B��b\� \H<&���D(7{�Z�ܐ�0��4 ס�@��ә�~�\@���_�@��F W��)�d���5����b!���Mc�3)d��.��yRd!O��+����*��j�eE�.���wb�O��G�V옱�H,G�4�5e�!�� [lK�Y���2g�I����r媬�ބ-�sT���J�F�[�������V����5*S�}�2�Pi��x6���1�׮ѯ�oK���"C8�/$�k9=�o�L%�"�1��(&Q�n����O_v`���|o�K�x��3{���dj+�����w��И8�H�j��m{�EƤ	D(*ӈ�*�P��J��K�
P}�S=^�xR��e8Beb6��БY�p��i�z�o1n`��tjռe�F�۵�׫��~�4n��㧁{AZ6��W2EZ�XK�h�d�T�=QV/��%�p`G�%�?%�+��i��t�,UE��S��2G���X��p�J������i*�
��1���0�GaÁ8"�a|�Sc\uWo��U<�F�W#:�'���	Do�j,,��f������7x@�Z�Q�7���:�L�w����+Ŋ����c��%O;tiܥ6����H%���f��!須t!����I�D���!>� ���B�F��4؏��@�>跤���\��J�6~��s�F'��,� -��C,b��8r�F
Ð��g��iL]Ϙ%0����&�Z�F��b���
�R���$ż�4$�59;�A�f���FE?{����������
��H�|�ɥ�8�k��U�D�zu��A���H�`��,] ;��¿�WyJ_��A�RhåB5�\ޔ�[6칔�-(*�py
�j�J{��i�:�4jجI�;u���^];���s@����Yضm���� t�t��e�����tk�b�z ���9wL�SX��ŨQ�
�.6�"�J��͠rs���I�T*FQ	��A��@`�gTW�C4%*�P��UZ0��Hva2���D�VX
�b��Pn(R�Kp�� E�P�j:��\�6���ߡ2��'�B�?q�	���\��т_�jA�T�A&�Db���u��ҥ~~��N�r����Ǐ:v��㇎?r��ѣ'�=u���S7<�!r�Zw.�1��@��}�B��4f�?'p=<��5����=���������������/]3k���n?<y���]��z���W�o߶n���{�o۹;����%k{�ꗾs���u�1�Ά�����|�o"d���,(�������Q�r����q�TB�A �C8�:,,<)8,���{O"��:�w�襛�o>��������1[^��2��������ݽ�u�&��S[���ܹS�f��?lؐݻw߼u/:>5,&9%���'��D�3�N�=yl�����?5��ih�U"�7�I��p�$�S��H��sZ:b�"za�̚$+I��� N�ș+,h��.���*�r;On�*lUG��S�8BM�X����H�P������Ҵv��#� ��-S"�"DU"V�4f�F��∵Z��p�F�S9:Ө��R�D�QIu6�ޮQ봨T�@{��g�
}||��L+����>�x�غm�/_߰����6�y�4>�4�iyX���:{��=t�^:i_.�n
iGiK:ieB�!�F>����w]w5촴N�$R��[���hAdJ��f�Z��:jě�������\�X�S��
�S&÷r�Vty�>_����yZ;>=N���Tr�
D�2�cB���ݿ�a�S>�|.>|r��ݛ����~v�Ц+�*K�h�N��Zȳ+��v����>�m׫DF-�P4����A���"P�r1���H�2i���4�9k7ｐM��Id�s.Θ1$�E����-��ҩX��K��������u���ׅ�{��R�~-�޾��ԼE���۵j٬w�_n]��(���Й	Qq5E(b	�<��/�Q�T�qj5�*|�:XG�T��d�2|@�Қ���?cJ{��S�rW�\��r�^�i�8�g��D� ��x'�%Oaq+�8�Ju&�T��>5@.�A�f�Z�C��;n�^=����ڳG��~�޵S�n��t�<z���p���#Ǎoөs��;\�\gwÖp!!B��
e��z�Q����+�]<:o��>C�v�ݧ��!�߬9��?|�����s����c���2`��qc�����჆�9r��1�GΙ2�ލ��dZR%���e+֜:u�'@p*�D��W~�?*U�����"s$.)��Հqǝ:{�����_�i����͞�g̀V=:5�ЮQ�-:�m�c�/�Gu�ܳ��6nZ���ň�kgN��;g����O�3|dϦ?�:b���A��n^��\��{�� B�@Jt�����c&�ߢ>����O�����GX-¾=A�#��^<y�YW�d�p�����2C�Ԛ*-H�� v�؞+*hgM\�
.�+��C�v"�*�5�$�(M��(F�
2r#�(,R%�*��x2�A���2��Z��NMc�V��+�z)��(!������!B�M��Rh�*9��� &3��^�p�}�5��T�V�&-�u�q�:�6��$��@����u7'�#��-gkisi}imiYXéo���נߩ��6���%��B�Ӕ�m�v];v��.6)Ƒg3~Ԅ�c##�9NVz�ʒ�P��l7z����n-�ۋm�R��Hg+���zGk��ѩ��̤���Y����x�ۗf,��`՜�[��>�}����Q�1��v3�4
mj�G�o]ٳn��{}O�߾~���D�G*��I&qBō��k�2%�Zo�m�E�=yֲ��|�T\�/�٧�?4�ܹkMv�нKg{w�ЫG��g.��}������u~�7�Z��nլ����m0��o�sȻ�y6��L��]lRfb5�¡��L���A(�R%"jT*�V>D�
�X������$2�MD|T�^�Ζ�EQ[���%Tg���O���3�z{%�/���"�T �T��e�<Ԋ/�[Ӆ5EH4��,�/��ez+\u��B
��.(�����C���{���^��oȀ��0�_��}��}���׿W��?�kw��B.�O���hē2V�0Mi��oǹ����=~Ȍ�c��9vؐ��Ϝ<q�����γ�T����ԁ!#��w��Y�&�3i��ٓ�̘0a�I�'L?n�����.A�e�8�:�9s�׹z��H��ۖ�t�Un��Q=p�����-U����8}B�p$"�T�I˺r�w���'����\e��ܵ=}F���)�e׆m��ܾGǟ�wlԼ����j߫[�^#F�=}b��L�������:����?.^:r�ʩu��뗶�:L�1k��9���O�3�
WZ-B�7�(!B��7N�8fd�n3F��$%�-�:�pڨQ����pЀ�C��6o��5w�ظg�	��1���,ԧ�T��%M�J��sD6��F����&�2�6��xE��|�U��!J�De%�����O(�z�k`�#���%q2h�`�շ7ՈD(Q+�Jn�ɬ�E-�U�Pou�tF�Vc֨�c�ܜ���� ��,6�lRw�تM럦L?d�0����7o㹡K}ZL>�x��:Ӯ�f>�f��� ��?Rg�&Ӟ�02�a������(��N��?6!�!u��z�6�q��!�Ǎ{/���i)�\�\$��tENOi^QY~IYaiiQEiɧ��2wA��^�ST%L�uB�A`6R�5(-���À�Sx���lxy#�e2��L�z����r��d�fg�H�����/�۷{+�P�z��Jk����Pc��+-Lx�\�*T��\�3@��N��`���d
'?��q�fM��]�}����`�� ��@Dضu�aC�4��m&N�ѡs�?��}�VpѶ�زq�z�;�l��x�~_���cn�D��X-B6�!d�d|�Z�x�mX���(�k"TY�a��"�:���l��*V�\�эa<�����Aq[	�Tp�c���Ls�����[��ݼ�M2El/�W���U-O���"��ח���B5�����QS�N�0aܐA��<����}��=�X�����=�����1���4S�0E�<`� %D��T�����������	�FL3l��sƏ�޺���}�L}��>3'��q����#�O�0|��%#�V�]2��f.�7w�ܹ�&�]>����jmNj�߹s#�h^��CF�� �����k���/S�}!�Epr�����.}ڴ�ܸ����	�1��<�d�ğzo<|r���vЭk�>�{��ح�ν;u���/?͜��f�TV
��5wN��sz͚3`��!��8�wǮ�j��q`��G3�-e!*�� �ۥ:G�5H��,�h��1��N�&��>]���Un5R�f�ۯk�>]{��֫[�^��9gɼ�k�O��w'Pb(f�5<m�Ș.��	liC&ߔɳ�]x�p��&�s���Pj,k�82<.*��B�!f�C��� a>b�ڂ����jYQ|b�7�6�5"�>ka���T�4Jee����/,rZ-�Z%濸�Ǣ�͆�wn�L�N�˯I���Z��ޭu�����c��@k5l�O7�z��ߺs����q�U/�l��u���I��f]#����8�Z=v�ﹶ���o[7nՖ�-��/�kKjݶi�޿�=֕+�Y� #5J̣z�*zv<95V'���"M�gW�����KK�K��e���|'�[��|gA!��Տ��A����v�����o|\s��a>So�e��Z���\�Q��@� U+c�b/�]>x��_��\[g�C�YBxg<嘫_X�SV�((�[�J5c�������{����z�Bi1�^�;t���JJNoظi��5n�c���4��D�;h�Hh-���1��wM7��a���7���?}����]���ܹe�v?�oռ�O����}�o��~W.���F��o�sӆ�5��(!��@���������9���mV�b��/�IIw��6�9�	��
E\b����D2Y^I���t��7M~"�i��pP���+$��\��vp����Gٲ��s���pԖ9�OŢ�{	��}���B��@��!jŻI��;����͋���;�q�F܅�Q�N�3B�Jgs�B�OL�4iR�^��u�����n�t�کc�~���ӡ�שs��>}!A5T�%@ h˲�R��)�X#���g���V��6xԈ��&�<o�����������3ƍҧ��9S@{SgO;fp��]�0i��i�'L�1qެ)�gO[<g���s "�5~̪����{�������M>rlxB6��bua\�K���N�e����k�c�;��`A�T�@A�;�i"3�Ǖ;>DވH�=ki�n��>���#[�ضg�.����ң�/�zw��DإS����9�����%KM��y���'��0q��у�]٩���1�+�7���t1[����9\4�!�!�%N�r�N�׭G��������Q}C^��g��+�ի}�qC��6j�1C�<d̘I�����}�X߻o@�d�6��J(2'Y�fkJ ��`+��
�S�0���*�f��T!pyb�����C�Xa��5IP-B�!��Ӳ3�t��@家�K���b���Z�X������E�UV�O�NGD�Fڦ�?5o.���7��s�ܪ�~�����c�¦S�6���ï�^���Ƨm7� ͸@�p�4� i؁o�#uXR���#�:k�đS�i܌Թ�Y�T��]�9"�0�ON>#��c�[�G��zt��JLee��Fѩ����������&D@�<���u(1l���㶞<�2~ڞ˳ܼ����ؓ�Qs<���������v.��~6�P��YEF�Xg����̏1I1)Y&W����'U��1��*�OV�+,-�Q�S#��� >�@�O�>��>�P�5?z��B�h��v:6i�УW��u�Ω��<u~�����u�E��|K��K]|�`㟛t��a�̉�wo�^��V�~�U�ԡS⬝[7�:�V�J��
��5=!!96V���*93_6��~��ݛ�W/�eegܾwW��X\.���{�n�������ǁ����zg�P�n���r���E��㯃_�D�ZS�U�YşB�)��p]�|g1�BCo\����߉�_��7�	��b�.Q��D�1Cã�S'M�"�Юбm�mZ�oݪ]˖mZ���i��k�D��	.�\&����$=�����MaB]�Y���z���	�&��<zȬ�������߶f���][4�ש�O�~i5z��qc���}�������2y��)cgL;s�x�u���lߦ[۟G��n���SǏ2����taP|�H
K��U�_E����a
��)B���6�F'v�ݣ]��Z��?bT灃[w�ޠm�onM�ڳY��-��� -��t�ֵ+���ҡs��]��ٿ���[���2p@`��~��<``�.=[��2c��kv1e��,N&OI�r[afK�^�]+2���)�x�n�AC�._2yh��s'��[߷e����X�:�t�ѷG�>=���5p��� ��C�7m���͗"}Yh��L"c��4> 0~��.��W1���:��*%��x�M>dFi�e����Q��^�����Te�U{����F��u��尹]�Y�TR�U#�>~xm��lFX��{��.��p1+-�(�Jxj��m<zj���Z�mھ�O={tY�f�͞�_�%R��Ͻ�5����8�$i�N�p/#`�g�.��]�mm>|�ĵ']�.>�׍&L��wP�f?������S���G1]F�||!�����מ?:��S��l9�c�}�^�Ջ�z�J�t���w@�F�âD���N�8��_sL��s_�,~��@��ߪ�q:l�߇���Xi	Ǎq�e�S���9j+b��*Mzw����Q`HL|z.H�(W~�r�V-q42�}*-��}�����������9q��b�3��z��;�|�N�5�����Ǐkծ}��._��!4bρ��.0hX��-�6h�Q�ޑXߒ�hҲs�ރ{-_�����wOx���닖�j�ᇮ��ԯG1|`bBLa^���2��15!�͋W�!|N1�yl4j&9'��������&'�ry�Јp9���l�|�^ˮ��t�s��UDg[�z+bp���]n~%��>F>#33��+ײ��A�S���
 �)B
�漪	�^4:7@�!P���d':H���..�k�ٸ���'�a������s�f͛6��I�7j֤Q��U4n��;��UT�%����P,�3M0�-���u��c�GO�>c�I��L@P8m̐����7�Z6��Kkh+O�6����8v��aF�8b����Ԭ^����iV�u�og�2iĀ!�BC|��m���9�p���_E�U����Y��2LBD�I��dԚ"q=�&w�ѳS�#�u:�}�u��%5������m[5lߦY�.m����޵s�_:w��Dحs7���l�s�FZ�nݵk�Ν:���c���u�֫m���Z���r������s���xr:GN��~o�)48����6�V8i��!g�,���@-Rm��N�_�޷u��S�a��NY�k��:?t8u�O[�-4�k��|�� ]h<s]5]G/�{�-=s�݂M���]0g��Q9���B+�B�_/�O�IM�N�_,�T�j�% U*�63|1�	��"����]j6(����߿�^:\Z�����NVh�7/��u��es��+���\���`d������f⺦c�7���؍G�k0rm���[�`芶6��v�yՃa%�g����蚅����b��������}�>}rحҬ�W/�	�p-$��U���f1X�!�e(E"�E�L���.qӅ�O�3�&u9�8�����hY�a<�o���<,ۃu\�g��	Vl�����_[�����$v!���$EX���(*��v)�0����Ԕ'�e�%w������f��t5��YI��Ip�sY�'��_>����F�#�����	i��e����G�W.?mҤYS�o^�j��B�O]<����ͻvL�3�}�n^� ?ul�e`�����]9��������� p$L�T_�{4y�hh��[0����S�jP�Z�A�AVzVdxXx�����t�O&3#&:H�����9�aI��TOQO*F�ƀ��;��{��+��˦/^�.&�������[�W�tl��v#:��,�w�D<�|����Ǘ�����|���%"�E�2�c�iج2�"B��%�xԦ
�:��c�/�����]�8 ����C�������]��.���'ē�L���f��ٳ���s���ɺhz]t�{�V-���):>���63s(|�MM��0��ذ�р~t��;�� #�~�t"���K�,��,ɫ���S��l��_:r}T��Ǝ�>63aTZ��{ۘ��p��uM�K���	L�
��$&"9*����jc��`���������tӁb��M=��T�_"�U�ϥg{z����Y�+:�N���
�\U����]ʬM����6n��~�F&����37t���b���zz��Ӱ<<�||������z�����ogm����������3|��'�#m��jڦ�'��UR�T>:v��"RY:�Щ��/00���o�I�cR���5cH���q���F}z��eзW�޽���m����5�/*���u˱�D	:?�I�Y�뜹�P�{7l�֧�<�g'�r���>��$)>���#��͇�l;�!M"� B&����'zvw��DKT	���L���8q�XMU���%�V,�[^�[SQ�y�
��_>�UV䟿x���+�&��/z�+|��[��o�h�j�����L�)Qu��o��g|�=�|���'Nߝ��ب�[�<�`���-�u�~eC9�+���;�(>��{�~P��W
Uܖ.� <@ÿ�ܧiCR�Ϟ\U_$��0؂����p����3D� -�fBQɭ3v�6��������R�t���P�An�aG.�QF����l�]N��Ti�252~�û����6G�7u{�ihGf�9i�Ƕ]|Dk��b��&~U�V���$o�΃��=�t��ٳg�n^������n�����}II��+����˪�Щ���m�}���7���ߐ߾@���a�����t����'w?�`�2`��e�6._�c�ڽ7ڶ���.=,xT��dH�.U��������-�T����֖N.[~��3&],)���^;������-��h�@:��r�c�O��10LK��}�ZKg�ۏ��� 'g�C�w��1y-~+��M]�r�Y���k$K>���[N=~y��K0ߓzܸ��'�^���l{
䴼�t�;�Z��S����~GC==���,(P7sUZH�l���P�	O���{�\γ�E�u����LM���߯O�O�^�г~� ���X+��>^aQ�����Jd8*]7X/Cf�j	���2�fc;�W�e��J���4zp����c2b]����������`���
&F���A��"Ç�&'G��XZ���con��j���s�y��#��Нջ/�%�л��D������"��D�'yRe]z�y���m��3̭�|�ڛ�y؆�Y���6�1�mk�������������,����xzx�z��U�}�,�=\������"#�m��q��F)�Efﾺ�lv%MRG�a�l�D(���O�[�&*c���������kg���k��H�!񁡾.�&�}��ACW����1>Q���]���j��X�����u� ��+�o�͂&�W����2���V��h��|Ӑ6i��×��tf���&��%��.3���/"��`At�-�u�Pr��	"�k�;�{��aY���05�NF�O���BŽx�s�����_�{�}��[��C���9{�%�IɊMˊIO��H��L��7$&<+, 5�3��5��3*�7.+8yDx����a!I�C�3�R҃23"FI3&eܸ��#�G�Ǝ�3*<9�#8�;$8c��1�F�<���](.��=|r��.I�p�׷�-�x�!�4��K�_�*~�c�]��Q6��ĝ��;�=��}C6�}�p߽/[��_��Oݓ��R�ԃ9�*��
xY�T4#o�F�?�mA��m?��l��u������۵ǹ�'����>}��-�ֽ�ɦ1�����de?x�q�k�nٱ{ӎ�K�n�	�	�N���t��}�O�;sr��c���{e߅c����W�ܸp��%���Y�x��yS�͛�|��5��[�`��E[VM\<c�%k�o�}�����_<}�ҙӗΞ�|���K�\�p���'�O[�x�y�W\�v��ѽ�/�u`uU�+"�4������ŕ�k
	�Z�����{xK��)�ʮϟ�B��)����٭��+;>�ѵ������!��HCh�����"�����C��3������k�D�v��U��;R�_��8<Y����jyK�̔w0$_X��X������O�}��Euaq]j�0��cc���>b�{��է?*�^���7 �~Ɔ �И�����r<�Absu�),!$����[��K]2�{�-�L"�?}t�ج�@WK!�j=D�9�+.,(D���FF��ʄg�A B�A&�nv�A�q���A��a��{N�3k�3O���t�{��]���/�*��P��J�s�PRyl��w-���Mfѓ���t��2q���qr�4���w�ۼy�t��}=���;G[���a1�?�������mX�{X�whp`@Hdh�p���9�R��-7J=�ˮ��i���<�B Q���~�&j��>νM��Z>y�-�-���`
?�k�>�}���Bb2F��'X���w#zW�� �>����?6u�	��{���퟽�2�<}�ʣw��$�o7�2��N�`ߥ�$y'E�N��ҥ�t�*&�TŐ)���� [�W�� �����0�������)�с���7�
ٔ�ܧU�L��'N�=5aҔY�>1$2��+z服�ǮH�\���09cqb��Ĭ�I�$��4dV���qC�$���5~�����S�$�\8j��iK���FǪ�3W��|���Yf���7tl�Q:�dM����9jŖ݉CF,0""!#���+��((}r���܂�|qM��{�.Q�uO��;u���S{n?�U�o�p�F��/�ίd��� Z����W���@��6�{5w��-��ߐk��.:��	���+�-2y����nې7��C�L/��y�߹���Tc�G�7��5��?q���$�J&����$���/��X1a�l�/,n�������N��䛐���x�E^��^1�>1�~q�	񁉉I(����L (598-�.��)4�#:�+*
�����	���LL�K�HL��:.2fԤ�+G��9f��{���p|��m�n}��Ja�����a�1�ꦒ�����W��ξ�nUIU�O߿����]��T��� .l~�U���"P�Q�o���7@�����T�'������o1�"�h�t�{�F%V)�e}�U���Ӫd7k��V��M��D�*��������'/��KkR3F���Y@+�w�n��,h0�_����}L]}�B��/߽�KqtF�,d���@�UA�h��cϙ.k��G��Nщp��!z:��<h���1*B�`O�� ?�S�����QQ�Q�c��3��"�"tw���w��L�H &ƤOH:��+���j��=:�S��l*k�%�_�ʿ��"���\W@���U����{�����P_wG�@�0Wko+;��z�X��8���|=�}�ћ�>�`Ao�`_���n�q_0� #�A�}�M#C<"���B� �8x�D��Q��fy��-WJռ���aE'B2I��T4`��F��r�m<h@��S�\ޱM���QB"���"֫��k@hx�0��Xk�M'nU�� B��X9��Ĕ��d���7��z9�r���z�;���F�%��H>#�^�%MX�#\�?��ǅ="ԹP.��"�X,��P:��/�9�����jn����S\&�Bh��*�8XZQ�����	�g�{���g�&M���=d�Z7��.]����M���2�/|v@�����aӜ}�Z��pl�9��o���H{�av�C�����Yy����y�fF�I�4��������5��'��-���D�6O_=#P�RC~�+*��+j��qU�l:.z�ꅊ��k��}CM������#]����F� ��E�����]D�W���"85R)�R�� ���!��.��6#�/H	�e��3x!M�^�i�f,]c�����k�>�V���[aeiIiq�R��㉻����ܢF���W�f,��dc`�pCG_��(��/��'d�G�����������W[��6��܍]|y��L���{��0��d�m��o�d�f�6���W������;z�E���NV��sK�.z��*[ݦh��b��k��nٳ����n\T��Z�L�ֶ��[�-*J-�g�.�����������|�(>ѵ�њ�j��[��J>�$��m����'�s�]�E�k����Ј��QdJVs+��������jkg�t�A��DB����}��f�� ���ta*�^��.���E	-!�P"�["l��fo�t�@����'maT2*�1CS@��Ң~������-�0��;&�/1$D�~������������}P�gDbPhl�p�S��\��Ԕ�;b�kT�=�K���.ᓼ\�@@����6?hR��[�������4����c���QkC;� B_�@_� o_?�=�_�z��9Z�26�od�k�@�A}B���<C����:��s,��5m��6_{s=���Ћ� �D��dy%�	#���@��v���{� [CK���H�>����o�w��[pDP�`��>v>�����K�����Z�d���6�e�C��:򰦂�������u ��#������g����J�wQ�=��0�Zt���i��'S�E�+ ��JT�����SgO�8w���c�n\<��y�B��*�(+*�(..+��0�Ɲ��_�TJ�i�.��nk���:��������Q������{f�6��o:t��Hc�!���"�����M7s��2�����`��>��},�Ml�M�c��cLl���-ݒ�}3����6r4��;m����՛�W��/�K^���54i�|���O>~��E�����������j�T���#�`K޲D�X�� 4��n7i@�~�H?e���&�o�wH��늓��;r����:j9���|��5/�jߔ@@�**)+--�(+��(�QTW�VV�WT7��6��a�ꈉæ���j`�f���`�{� #�c�H8𥁙w�A����z[�:�:�eY�'��s0��C�0���: =��3���e��2��<��,�hP��P�A��~��.���)����ѝǷ��\��s����������������b�p�"��b�dbE�V��B�J��B�.�*U��<E+G��R��+?RT_%ߑϚg�pJ����`����ֱ�/EN�7gǬ��i��M�_4�cv"��/�ڻ�
�v�%�&��`��]Gn�ћ��������u'im�ɜs<p�^�ȥˎf�3[�2�-�~�ĹG�NM�lfj��r�������ɀ͌�Y4�45�4���8s�*���3�?��D��;a��s��eI��&����<iԐ�CS"|���X�w�0t��am�mg��h����������X�P/OkK'�A�v�ή��!��I!!1��w�ʫ$�7��N������!���k�ׄ�_���?�PD��q|9�'�r���Q:z�W���#�C��,]���:[t���rs��pqswr�p�7G������r��1��̬��e?{3Og;/O7�@Ht.�#o�|8n�ٵgsna+�b�=B&�L%��ږ6*[0�n#�ކ�f�}�n_zi�B��yoK!`<��x�� s��H��L3�о�����+$�&�ٟ5k���G�,��5V��h����z�z'��BT�>��qq݉��w]X���#W��Z�X�!կ�w��~!_�~��L�T��ju�F��]KK�V�QH��G1_,ዤ|�THf����ĮŰ�j�7]����E�&N�1e��Y�/�_~s���s����l���k�Zr}��K��^���Ҕe�-85v���.��p�[����h�ګ+7\�u�%����G�n<p��˫v_�z����Wn�˯i`QrKNcH)Lt+tg+���,�P�Ri:��?t���jk�7�%Zt�B����#���v�#�H�]��.m��:����V4��=�x��g�`�S�=,[��B�D�����{��P���B�HWI(�J�R �������ӹ�N	�����Ƌ��9�'���b�ɜu��9�`ӱ��g_�.�T��������{����g^�T��|�3�6}��ĳ����?����У͇rv��ٽ/g�����O�~v�B���7�ت:r=�XG��#�l)�-��nkR�P֬ۍY#׶葨A�*�B�nI!W�
����DEHTE�L_u��A�/�u���;4������f�.�S��3{�S�](Zz��D���#��Ef�|p�B?u�a�ɣ~J�u�r>�A�n�횺dɑ��H1	}�@��f͗r���y��E��/�xy����'�'�02�0247220����}���g�\hefngink�z��e����d��2j�{
������}s�Xn���hk7~hzB�7X���������Dx����� �--����52���ϼwoSt�x/[c;S{S{S�@��Đ��a~��!��m��)B
�/׶�����EH�p)��ē�8BK���s�Y��g�#c3��<�\�8��3�mo�Dhofhkjdcabmejai:��/����A+Ks���݉p�Y/k�~���m���d=�_ʥ�!��S��E%E\OAEH�P�D&Tw�<y��7�����|��-O�����l�ˠ�*BS�~&�FYy�F��g���s
���H!Y|�aɘ�;F,غ���:�[N��ҋB����IoE�Z���F��񠌺�l���]˩e+i�.��^�,��!G��G{??��E(�%2�B�B#W�������֖����f-߾�hmoi}עn�p�"*���V8��inInQͭ�/�=.�z�����W��ܬ<�����+p7�R�<!��[�f������o����K���_|J��}�����˟��n=�7��>l���|v�|l^=���U�@��2It1���[��f��U�hɚb5\�T.T(@�:�D!R�jsY�nQַ(�m�th�D�K�aH��s�v���9feN��R�܎�K>�OZR/l#)�����&�v�Z�B��������mG'𮣫�����C�n���U"$H����.TI����죺98x�w��^2�ݮ�s������+��?��U�J%��R�����4�V��J��B��s�{ϗ<Wq�L��S5'�T�<Sy�\��s����2Na)���J�3�B:[���)�6#���K���j��n�����j�D�j�6&��9JtCE+�����0O���>���p�����f�
�E֚ʷHMR֎�͕";����+�!�.���R#�ר���THh��*%��JѸ-W�Ȏ뮕��q��9��rq8xʍ�r�P�i�Q���|v���'����0�������������������������������������'4����^��~��L�A`*h��8%b<a���V�f�!��Ζ�����6��"��6��-B++/[[o;;?;'{H�p�nk�hmnkedm=���aL���;�+q�"���z"D��@�6ɡ%���o��sQ��K��ʟ��E�K�R��d���Aw�/�q1��-{O�7)391������ި�����i��������Q��`��Ш��!��q`�IoCct���������Q##�~�>��#�0���ܯ�>o���L)��=}GcՑ�	v��j�����6:�q����@��Q8h1��LS��,m��b�2�<��9�/�w�Y=����]FU�%X^G-]C�|`��QH�=*�e��BI��~� K�a������q�ω�g��?a����h��E"�P��ID�\�i��#�8>[$`�@#�\��@c1_�d�Ȼx���3w7�����C�^��{�:��#w�w^.�p67d�����=���C��R��#/F/:1f���n�zh�曯�%��ޙ��μu�l��b׍�'�/<*�k�c�RC�%qpd.��!��4���S��D�V�� -��:�m�lxR)[$�����[pE��� :�E"�H���t�TE�6���Nd������kC� ���Q��?���h��n1�J���u��#)$l5�-@��P
�|Z��}>;i�r3�۰qqc7/����]܆���IK�R�Iˬ��Gf��r8o���#���O��5l����N�ď�ᙰ�=v�s���ٮ�s<#g����������1u��k��l,Q��YQ-�X�k�%�U�9S����i� �|9
DC�]]A�ȵ}ԋ��jf)�E��|'���)V�o}���c��.�>����;������1_��WJ��K��T7#��|��6^�mCR��8[&�}GJ��'��Ň�	�����>,� ��?Fl�=�۵��k�v�݈�Sv^�v����'c�B��2�S����b�c��cc#�#�#cP�C��_���p��P7�� 1�EQ��1y���/R��5�m��l�mox��w��ۆ���{�G��������D�xEx{�:�}�\���,u"���I
�ڸcGa�/�S�F;[��#Bh֋�ͿD���C����9����F��&�-�1����ع���U�͟�`��Pe��������`C;K[+;s��n���������=|	"47�����̬��Y3H��Fn.����&��32��Y�W�Л��*���!��Qb\0b5�s�z�wL���OD���u�Sk&�Y;&�����Y�O�	�N���
����qp��>>n���S�l=����]�����SF(�����$�[����ut�s4_���F&Y؂n=!j8��t)��T�`AH0��:�9��u����Q7�S	uFtK�)�\�nH����R *w�@ ����w��0�"�HB�������Ҽ��ǯ��yQ=|�ȅ[n�5�-$�)����Κw(��-n�a���BGm���!fƒ}���aلN���0q�_�����C�m���3����-i�G�X�5�;n=6�5��	�Mf�X\)��.,���"��{�W�(��|�J�Dw�ס�%�V�� �X�]j�'�uJ�A:�R���4���^?a�є��&m�\y�9cV���zV���>F�%!I�˥G"Qt�v����>�6����p������3ם��O��������W,Ϥ�q�M�pk��3Cf���Α�ȡ@��f]��a��m ��/ؙ��x�,�����Eg����x�ÍG��Y�g��+I�XD̘����'��ƕW1��%5�Obs��9*����� ��)԰Ejh%�:��F�ZB7�P�*@gA�dU+S�NWu��V4#�
�,�K�q�H�<j�ҏ�E�ޡ��@�����,���[?�ȋ%��!|A�Uȯ�5c����P�V(Ф��l.dA��P��-��Q"�O��B�6���a�_��y_0~��5��o?p6>}ThDRF�Ȍ̡�����ӓӒS@�I ?��؈�x� ��g�5Q���%��4b!(���RF�ﰕ;.�ٲ�p��Obx`b�b�/`1� ��e�Ա�ϟ3qLZt䓕�3$1�OJ "|=L�L;x����!��!�ə	k�l)����2QN���	ל)T0E2&_���������/�O�o"|��K�	��D�!���Z���O��=s���KF|��̔�Ȑp/gct�#KcGkS[3g'Wg[7Ww[O =-aĐ��I�Q!�{����ƀ��IH����[TB��Y�c�ʯ嗑4�4@QC7� B�n��&����^�u�[H�w`H��������^�_W�w��'RUٍ�(�<=m�\����LϜ�8i�����1�<��]J� �݂.9!�@�u��.yG�3e���tI'C�Α�c�; ��@��,����E��P/B�*3:�gS�$B	T�=�I�={�Rb2OM����\���(;�<v��1+��.�<�`�/�]0i�Oh�1��-�Q�9���:�`ȈuG��!�7L\{�^��Ae{n�����-�/g��>�+�.W�;��.1{SNI'B4��-���J�B�^�BI3�i�D'Btߨn-|y3��{�*��](Ӡ����]��!�����^�f�.瓯W�+��U�"�����?G3\�?E�Їi4&��	��a5C1cñ)�O��=�U��uf�;5v˩r��5�7�<����u!�1�f��7b�����з�/���l�Ѕ�����Z��l�B��5�KX����b�1��{R{�qyY5���XRM��1����	�#�r�(�U��)T��S��>��JU 
S�LW����4�;��"V�Ӈ^2�`�.;_5��#6�Ъk�OX�]��zMܶ+���jŰW�沞�>~I�����52b���ˮ�+wܩ��7�n���P�l�^=n��6�RUk�̣��E��>��L!�3x���[Ol?y��ٛ�#'��$g�5dĐ���������
8y��?~�O�ő�T�!���ӄMLe�#rҦ��*6lٓ���c��F�ŝ?���%�Ў��><5>)"aBԐ�h�g��J��������>o��a�~nc'M|�_ـ��HR�!���R�� ���X�/�O�E�������#��\�t��=�>�����/�߾�h�fi
�0����~���������������������㒅3[�b!��������a��i��"��S�F.�xh��U%M�R���������&!ݘW/B�P3c�z/t��!I��,�����A44��?�䘀�� G���~������7g����G�<,��(���q�N��E�����j������r�����U}�(?�9�NT�2T���ge�{D��c� ��'�~@'Btf!et=�h��D

ԃ>Y�k�
�Mة\1�	���5�T�=+äL[;qÙ��G����҈q�G�>{�D�6t�K֚�g�N<c�Y*{P����/~���W�d�/?�9Wp�)%a���5�Ͼ��/�U�2e��xQ��@D��ԉP.DE(�_I���"T�7�E�'��N��@â�Hx�U�«��D�V����U$���m$�{����{K���-W�f��?�u�.J�*�a=G3i�A� �N�Xx���%�=���~�b.�9in𨵣������yG�~x�c��\��%�+��nY��1hr߭��n�Y9t�ɀak|3�N�t��+��//<��\u�k��o>-�,XVE��s,���P'BWPr �|��!@�[E��U������$iޑ4���OȢC��/sM��0mϝJ9F��)���G��:;l��J߰?].��?�4w��e'�1�ϕ��U���9�r��+C�^����5ȑ��kD��|Ά��V�F��zИ4o���wμn"�#��m;s�ԭ��7g����������������

	C�v��;p�T=�.ԋP��&х8�����=x��rj�	�'G'E�\����r�t�[U��M�M�	ό�����a����84-��:_�b��^�~���mdtԽ엕UT
ME�*A���`�!4�d����[�P����_"��J�i<vAy9����!�¬��xyx�y�A�*.�)d��vd�`a���h��l��b��f��	���xگZ>��E)��	�u���tr�I����vp�ݺ���Y�K������*���#���yXtc^ᴅ��|��⇥D��I�s�g�xjCΫ'������£��B=���DF��K���]��y��Ɠw��u�a��F~>^��|."�o��]�{Y'h�TF�s>�̃�s�����h��%�h"U�&s�="ԣ�*��ǻk��*��]�!_,��J�<�K� 8�.P3��@Ie��d*K�j�4�2fo���F6��1�3�;e�����:v�o����&~�K�
���6]�|��3u�K�b��%�Y�������+����ɛ�'��X�2}�mw
�EXA5��Hb�i\��D�&Z]���i��X�g�y.��/\"i�j�L���wG��DD��%{.�x�{��&[��t7Y����M��w����G�D�_5qS��q�f�}�N~���?�3cq��=1��O�1o׽K���:ͺ�/�o�:j��cR����siC������ \ظ��F�8v������Ҍ�|'m����U���T���ñA�8*���
O�D(Չ�/�E��D�ӶQ�*��G�`+M��#B��#M��ӎ�$���d��fDЅ�S�Q�zW)�H�P[-��s��$�-������یP�?Y ��\ҁ�?"e8-A�]����G�t�S�x��f��
�!���������;9oFL����ޡ@щ�/,raPd�wP�{@�>��d�y����"\��
�����Ԩ�fą͚0bdz|u�K��u�ȾqC҆%ǁ,�� B8����09.#!<&�;�΅���5��W������ܵ�",'�x-,��ŗC�� �ᯮ�_�_Jϊ�43��]t�ͣ��ݡ�%�3�D���������9)6>�֭��7���5�f7�����������������z9�{:̚2�$�������c���\��B<}�]�}�\}�\|��c��%�)�����r��tA����6�g��Y��&���'%�d&FЭ�m�[7wb�������Yrx|�_b�s��[���Y@B?�p��E�/<�az�OI��vƶs)�6EO\}�ZP.�1~]����W�vO�w����r�ĵ'�΍��b��g'��Eo	����,n��F|~y-�I��6����&�x*8��~�_t���� �2�
�J�*��Gt(4(hxB��E7gi@�L���C�Ҁ�A��u�CY����w��v<���L�1c���y�mW�5����_*K�}�#k�����	[��{�Xt!W����I.�y�d������8��p�Mϸq��lഽ�e֑�X
���Y&W"�T�L�E?��~���?�A�������k����/�sO����5Q�6
t���<�R'�nD�fgJд
�e��6��F-�9|��*����I룧n:�O�R�r�\��b��&5H�n��F1�����1ݭ���|��������6]�\| r�c�0g^�>�۟]s���ST}�q^���֝|\t�UiE=�è�2�Ȩ�]SXR2GI�i�|4�����#�\��&�]I�D�����.�B�m�t}�	4dEG�p�?�ԝ ]��Ruq�]<�{��P�E��*n�6�&h�����ת;i����ߕjS4�.�}�G��.���@���U}f�l�{��ߙ�Q����~��7Eec'N��vuu������vus�O�Bא�vw��t��0�����\��Б�FL��!���S9d�+!||9ڀK��3���;8��n���� <?;;�!^.�����IqHb���X����@�`o�`o'w�A����c�&��9�����E� B&���ղyJ6_��KyB9�#��������#B�\V]�:��LG��0x����1Xr����ƌ��g;����������������\������W�x����o\��`/+cx����N�>.>��Y	c����������A�~�(��$��w����	1��1	сi�!	�`bgKCO;�p�����h�� ��8{�$a�p���ێ��U3v�>�)�QZ�@~��ZٝU҂�o�?H�-w�<!��ѩWkO��}��V�U�`DﰢV���"ma)ѵ�(���r�?+�Η��W�=�����! C��u��9 ?��U�鐷����i:9�ti1:xr!�#��Q�c��Q�jY�w�LYr2���rM��{��֜��}� f��+����F52��S�1���%��7a��<��W���H����9j��q;�I�T
7���8n��+Oˉ���DHc�A�L�^Z����_�P��cA�v��k����nM�~e��{��?��a��S�����c�r����|��_E�&K�=�-���u��ssv]��}{��]-��NX9q����L��Y7�;��p��u��	ǻe|���	�7�xT�y�Ƌ/�&��x�U��]�C��ɡ'5��H���^y�yYZ�ME���N×�yZ������V�D�ǳ�4!�%%2$`A
ފ�7�Ej�$ҒEZ�f^�Q���+��U������RI��;���~�l�����Y�V��r6�1��V��C��T����.��'�f݉�-�P���Zu�Jѩ�u�%���\ܪ����(R�.��V����#L:���Sw���O�4%22��������������������-:A���ڠo_g//����T�7���Y�$�����L/Bh�� �E���v�v07�q�I������D8"-nHJ<�����������"%>pؐ�����h��`�c���4�b6����*="$3����+.ƒi�82�ƥq�T����Ehk"�wu�w�dcadm6�fPwG����|��]�|]���=�<P�7�2�o?��z z�G�{��X�=�����]}C��"�G���JkxMdi�YGCgM�l3��`��C������;fĈaY>ή�@��{lpx|h||pz�Oz�S��s"5p���#+b҂	[N�=�`�[�3�ϡ�	���3����b���i�"u2d��m�+�A�`�]x�� Q�%&���+��ނ?�P�翸�o���V�2oQ亮B�-4��] �d�h�.�v��-M�A��4�71�4dɁ�A6�����d�����ǭ�Y@����/�;|ގ�L�x)pԚ1.^,f�M�8j��MWG��>q��9K��C��}1k퓫��W���0u����+���3{F  ��IDAT�0t1�
KHe輿D�������*�u���mA�;��z~�D�RCd����Q�`[�{�����ՠ�Ϻ���.T�E*�gJ "��D/B��c榣�6���}
XmS��qH�x�q�{�L��I�Y��'�5�I��.ڙ'�����M���*b<�Q�h��}VQ�"&�pJ��1=t���?ɯ�odY{�oʦ����WTc��M�F
�SX
SI�B�k#��bE�@� n��*B��CԌ���o�eˋI���Jn��}�J(<I�WAdA�@�)�R��F��*U-*t5�f�Jss3z�s5� |�M��F�j�*��
=��A+�k$(*�\)G8���V.�;jԨ'N<x𠴴tҤI1QV�}{��c�n@h9p� ���~Ɔ&��z����"�RQ�2C��(�G-E{e�#Ao�࿱Y��v������掖��P���p^x�{\�_Fx1~hj|bLHx�T2Ф654��⑒��n�����z"Q�E-��%�_��\zDHa2����2�Y���<[Ne�(Li}������Z��6f��<l�M�,�;ۙ:X��4!�����~��>nNz��vEw�������ڨ��������D%G�)��X� K��'GkA/B*�eؐ�~����'���Jwqq1lHTh(|.bB��B��3#|Ӄ=R�\��,���88����	�6a��Gf�6a�֛�9�����S����@!Q3l�YO�Dj%��/7�.-!�����,H+IB9U$�Q��(�?�����I�8�I�~OW�h�U�Ȋ�P�s��D�KU��j����#��ew���li���e�ʈ��ZJU�KTm�Z���d�܃d_x�+!(kȚo0+�\�h︕G�yt���]'�����헧o�<n���s�^���A��L��u%�w췥xd��[�֒1��D��z��Z��Ȣ�bu[����O
��;��-�D���6�w���A����NN�n��,9:I���ы���V���~�@���ڢ"���g=k���6�?���u�G��OkN?��}���e�瞸_z��t�������ҋݗ�Xr��]I?��x��;�����J^��o*���z�k�v������®j"��(MTv]�c+q<-V�	��FIW��-�D�����(_�
�0O�抚Y�f��G����u��+��2w���g�-8v�U)�������,j�H�*�F�R˴JY�Z�?�j�mZ�8oU�[�q��])��&�vH�b	�&��E�b1���Y$ң�T�R*R��
�X���	�F�>u�����ӦL���d6��d``d<�Ф� ����{0����Ĩ���o`�wPЎ�����pt�Z"���l"����D�����(m�ָ����H�hרN��&������`a2Ȥo��{L�?4��<�$96lhzBFrt|dP������� ��,��񴏍�	���ppt�V�.W��Ș	ڟ����K�ItjuS}~Y�z�@G�(lYU=�eA����dA3{G3+##C��&�-�����w������������������#��`gganibd-I��wþf�}A��^�����>��	�1�U8 O�s��\p!�R!���08}������!aa#F�JM�t����rtp�t�	���H�61%nl�o��SD���~�}�����L^w�I7f��Ky�F%r�	1q� `@��W��;�b��{R"B
�_)�->�MkG�o���EW}�g7��d��*V�En����g�M�zg@M�Q��[>����?�mH���P�R��U������=s�����3?>.SE]Wڠh$���TQ�ɇ!C��ϯ���
	�<��Y��Q��Y�iq=��AP��6	
�oE/����0�7e.V���b%%A5�W��U`E�xq%N\EU�$�q-M\ED�����E���'�����)�Ū���H�)o���勎o����x�����"�2�����bmU m��("���[�ǯ�ַlM;����j��T��)�wJ��w��M�{kuR��./C�L���M��z~k#����R�TWѕ�$I	Q\��4r_׳^�0^TR�������4 ��
<���w���@Az|]�yU�ȯ����VI=��_Q���jH���+-�ַ#���r�Zq'U��W��]��H�E�V�H"d�Z��I��-2s��:���^�R$���>|���R|����!�h�t4�Z�R�L�.�&Uk�Z�hiV�p�QJ��u4˥ 9�H��ᨕ�����*D:$@.�t�ļ)S'�=w2'�Quu��S�Y��8�2�;�o����5�ݯ�E��}�0p���/��{�����b�
z'�� ����88&�����a|jVj,:D��q�Ҹ/`=����@o?o�`�@_�� ��Ѐب�����P8^n}{��IY�:9Z�Ƅ����ckg}�ȱ7yE8<�˓���9����XzDH�Q*j�JK��OeIHL9��Ba˪1��%��v�VNV��6.��f���&ƽLL���P<����]\<��<ݜP�ml,--L�'�a�^�F����^��M*P���F�$�U5 X"K`���c����|�K�R�1zѲU�ΈML	
�	
���NNO��>:%qTDh��G��]P���AI&.��^���(�i2fm��O"i�W���.��s�)�=a�n8�z�p��}���[�bĭ{.�9p�K����"��8��D�\�j*b���R`�^M�CϹkw�t���w����F�{}�?v��W��3Aԁg�f�_u�I��9z�$f�^���/��MDY�y�擸I�BF-�񪢆,,h`aE81P��ժ1��^E���YX�Ϋ��7��EMҢ&Y)NV�U�8�8V-�U�a4`h�8z�]��U�D �z�� �	��ԉu!�:4���u��������ǳ���KYC��&����|��Ed��5_9�,IM�	RlbJ%o�p[:���lm3M��Jd��I�[���*Q 41�a�+̒hh"Y��4�0lmK��T�S�x~q3���WIxSExSM�K8]�UNxYF|V��)�<�o|�ې������Goj�ǹu������y�o
�
J1���rLIecYMcEcS%�TAg�2E��Ν�����������o�N��W��W_VC��Sy�F/B���,n�w�NP|�y)?aҖ�I�G.>�l���w�/#p:?��ӛՌf%K��h�����	Tr@�� U)$
9�����Tꊾ�T�]gg'�x\�+���X�N]K%B��'�q꬙�/�{��aYE��iS"��m,��loT�����a�~�@�&��n^�^�����)���i"��(ԅ
!.c���c�Bh�EĦf�GO�ψ���B�cgi����y�C�|�B��"B���`�������T&�&����n.���)�o��|�ʵ��R���I�,t���_"�U�c�w�B
GDbIIl
G���:;Wg'OO7� W7/;��bi��F�"B/gWgw{'=>�.��v��A��������������,<:���*��DH��h0%х&dS!|��3u�|/����(O� �����Ĥ���,W�`�@;�@��a���F�[���x����Y}�����'U�2f��
���Zᗇ��+�	{���/�4	�٭_������9E�8�jR��n�gݢ�btN�?�P_A�YMˁ���g�T���"���N��L�8[��qc��c����N�����v��CG�C������ko �o=���]���.<.*�2^��
���4���VRC/�e��Ћ�i@a(�g7pK�D@%TcY�XF=�و��ᤎȫ%
��@]�d��@�����3�< ^&U���U�~�H�k�#�.M����[M�"}G��'�v��#A�� �bȾ�U_9�/ O�M��C�u��ɚK��F�+VU�5n#O����D�(C�:���z~�� :wE�.7*Аy*p-���1�Z���Ӌ���T�_M 
j�y���ʦ��We���g�O�P�=|Yu�i��������ge���?~Y��uU~QcQ	������������!�"|Fb�p0r���'��9~���zY4~���a3��|&G"��� B��������Ex�gM�E�o��O��/e�ψ�w�m���Z��Q*�+�D�����j�>D� ��t��-o���v�]��9�C�D�@��A8������ ���^
tЖ���U�i�;w��{/�
��bfc�nu�۠�a�~����o6����Ή���h��"l��
���<3���e%&L�9:#!#.,1��������>�v
��@E���0"4"$���������������-8�?"<8$�/"",==�qγ��Z*��H�l^�D���������D( �����)�Z�������/��7�������x����d�a� �Y�p����su�4�I�}���m̼<]}��s����"�+���5��EHf���:�@�y�:?<6�78����������G�}\\}�܂��6�r�wv��=e�t��{��w��#�_�S��*�/z52M󽚩�E���>A�ߪ�H!�@��K[�|Ua-�UY�~�5��k�j��?d�9��lA�9����];�tS���pB��U���o�鋷ݫ�㼇XZHT�Yp�j~%F�a~�##�Y�<j��pq%Mr�I�1���r#�WTM.��� �Ր�ki�B�����zfi���Tcx�X�>�
ԃgՑ��/�Q���e1y�P
.Y�Ǡ��<%�F����IԲr�I`����w�]��<�|ʱ��T�j�j�����;�j+)rz�*^�����寈ֻ������ H����L�P�BE�s��~'K����^aژ#���K7Q��$.�^h UX:P�H-�'��
� ��ei���\\E,,'���K1yE��� ��b�K�JKJ+��1x|-�\Agf7�bn�Aռ�~+N���~~ݩ��gm>6t�Z2W.�h�|%_���I;U��َ��"G5%O;8mý+�D�d���\���!v~|��b
��"��B�Z)o�UvVK[+�2���%��(q��'��3@o�0[��kiz^52�hR���琕��wx��:�NH�.�x�����V�>u���{���H1�#8���֠���&��F}A�}���Ehn����_'�ʚ�᩵DZ��D�6� B�aK��&�:����̘0j���iq��@Og �⠟��������}���� ��CB��O��u^eu=�Lg�x�G�\��Yb���
���C��@��%�L>��᠋%�v���%u '�p۾��l���ݼ ���FC�!z����>��3��?��'��������� �y���¹р~Ɔ}����8��:�����z���-�#AŒP)�?�F�zb�L*[�%36n��m��'�������������	~=?[�@G���cf�%��v�5�i����+�����6��)�!pL�g)Q8�$h&��`�?�~u�cA�{���grŊ���??��˚�*ں�,���]/�-o�e�+����o���T�E�����M\u�y�݌�#�#�c6]}RM�K�uB�v�#�,��_{UWO��Ѫ0�Z��S�c�.P���#�MܪNe#Jy�ˮ�0p�^�xF-�UK������j� �DL)��8�+bsy|.��g�Ib5z�M~�l�.�+ a�-B�\+ȅ�w��x��3/>�z����9G��l�qױ�$~gI>l²%��<zg���'�K���7x���.��p�������K��Vm�D���em4%4P�!������p���3��o(�k�Щ�6���)"0�x:�vDPGB��Ѫ�Բbi=���/�%V ��rlAySq9���	�WT�˪����Db�\�`��Gl:��E�ۑ2��U��{��$j���',�F��%�f!O&�)�U�B�t2;�;d��K�v�淉+�<�i��t��=�#���~���f︽�'�6��=�l~X�0d�-�������9��FR�����א��D�Zt�rl2{��^�f̘��B��uIs����s�!�v�Г����^�5��
�G�G$u��Ws���#�_w���ۏ�\�;d�gX� g�~�ͬ�m����44516h2�l���@SSSGGG�]�A��M�:,�YF#�����"����<��#0��chj���8;����X ��:��Z�YX�XY���Z8�Y9:X�X���������������N���qQё�˖,z��EUeG�Pٺ�A�a���o?~�%�_�o�D(�R9,��nI��P�@���]��'���y9Yٛ�[��K��},�ۛ�;YZ9�[ٚ[ؘ�2sCcKcS���p �G�Q?3��涱0��������u��sv����7�C�I,"u!���B�N�te
:�v�3��8[WocK{g�����m���<B]���b9�Z�o9I��#s��G��τ���z8h���I����/��$zz�H��rm���C�l���t._نc
�-]�21|)�/��P�Q�6j��q�t��<f�O֌�
]�VGWTʐ�I/=.�J����!��i��{Ex[U��5Q�8�}u"<Y�#��H�F��/��	jp|��M,ԂX��S �Y�ȃ,��`-M
�CC�[�|&W��p�\:��$j���\H��"�PR
OF��E #�K��������X�
*�?Ͽ����'�O_9e)��~����k2��9�oןսh�\��(��xR5��z���{N��Y{��s,����I���Q���9O��_�&B��&�/������뉣q�Ȭz�%@;��ay\XR��_��[Plt"Ā�  ��+����J����ג�g���~[܌<$��.�s�uU�ZJQL_���S�rW*���<5��,��k��	?��t-�F��3���o�_}�F������1���w�j>#M c�=|$�>�j��[�������"֌�Ϩ �j$t��a�/O;�X� �ȹJ��k%�^��o���]V��3o�+��^M���Nf�ۙ �ȑؔ��7_{o���,=p�����N_�1> !���w���������������ނ�pbff���aIE5��C�1T \�D����3c~߁6���x8���0 �:���d�h��d��b������ �2hajlge
��`;h�Ȭ�C�&O���WP[���2��ү����AS���o���%�_�_�?��M�2H:��Я��c����{���Q�҇�9��7�`����Y/ӿD����������������ffF�t;���NL�����ܤ��	�(����[�-�&�(l"�I���dp!
��%��i�x*�TaN^�቙���2�ptУa X��)��)���o�odjh��m��V�	:�h֤P� ��($N"K�g�	
OI���^5A�u����[~"S ���:�n*J���qd�@,U���]�r	K�p�Y���ڙ�	�*�����c����e'���f�9n��B2"��(}L���A^5b�HR�gS�#��[�#��uX~Q�%�u��F"�� ��� Vc9����Z,::h"��:2,XG���Ut% "lbʉl1�-`s<K�%�yT!^�m��D)*B]���ē�x>��
S@f�.\�}����+7o�>�ȩS�?r����> �n�9{�5O�[�g�ۂ����ȩ*���g�~��qM윭[nf.�u�u��3N�QIA��$��j������,B�4���eZ�"���dV��@D-�?���� �*,��Bn���h��d®c���j��M�3��S��s*��V�`T!W��K�`%��?(�/�s�4*�r��}ª�M�o܏�ٗ��{�᜵�)��k~G�k�\��L�R�y�D�V�����f��'����t�[���~��lC��
���/��J�P$b��K��e�H�{�u���b��r�B8��ә�l�^ؠA2���s�7��0zRT�p�����a1Qa������8���LKK��aM#	�j�T6�:ԅBA-]喹xڶ+>���F�]lzٛ�7p�6�t�<t��@Գ�yz8�x��z���z��x����;�8�\�q�53"�q�啘&���R�t�_����X~aM*B!�CՉB� K�C�8t����+&Nk�dl V31d��V�����d��oVo?/w_O7���ͼ_kcp$D�AP_M��4�׻�~}���D��_�c�"��Y �He�	4.�A<�K�'��1��y۹ػ��qP'B+�  ,?l��E��m�,�`�b
[�#s	d6X~>�¦R�4:\�����P"$��M���{!Г��T��0��K���Ӊ�-o����.�|^�H���E�X�
ϕ�ME2���S���yw�֋c֞�����'s�Z��Y<�T�${7yݾ�z<���6Oz��$n��l 	�j�U���_�	�#_0��&fU#���^QG/���70+��cdt=� ��n$q�bȂ�T�bh*�j���ld��Bg���l�����t��`���Q�A�6C($	��h�ׂaK0a��� ��oݹf���V�?~��1�'���tɞ�'��F��>vs��T���k!^��zѹ*NI�F�=jޮ��
�o�R��t�E��c7�eo��5	�p��"����f���"���H*�]��?�P�/
����2\Y��SU���Sj��F
��B�c�+��;qo��;�o���f�雏�h���s���u#�D�^������o�b�5�u����Ҍ�a��+.�$�>"��9����λ����I\ׄs�soaq҄ %��_k�I��bW�Xt��������oH�;���RE��3oTH�g����g��D���>�J�{�I\v|[vݱW�����H��m�v�]��̚�g�FO�����"�@E����p�^��P���B}(l��A�~#W�?�j��UQ!A��6IQ�>.�����~E*?og ��=,�����
�/�ܝ��=t�7pK���
\�dAmm}S#,H��@�4��Fo������C���K
A�t��:ԭ��k�1$��ӷ7lؙ�o�l8���ή_�>�[�~fFN��l̜m͝��:ڸ9�z:� #��]�͜-Z��/�M�Gz�2�p���KJ<2i؄�&zY�����D2�L��E�D���ɼ:"���������='�����6b����S�MN:H>5c�����OZ<r���.</jh$�I�=H��O��!��H��H'BX��n..t�%��
����eA�b�r�]�JxR���9����'w���S�h��;��%U��\5��F��'Ϝ;yﾓ�/�۱��}'w8���}O<t��ѓ��;Voܶvӆ���lرqǑkv`٬���>z�Z�pp,}�C���:?�:�#
����,��A6Q�tIY�$�P�l}�$zR�,&Jq�V�j��B��� 3��$lE ��+�r�� G?t�k��z���ȦH�U��-OL��$8>=4)s��ŉ#ƌ����۷_��x-�,���gW�>o��qK��)�.��f���K���I^��O�r����%n� �d���6�E�"�B��w�ꀓ�G��w���A�-�W���� Et�(��R^G(�ŗ�����EU� .=��%� ���rPS��o�V�i5$�L�̡�G�ݛ1}��'.�<i�����\�vѦ�ç,:s�:�D���-�vx+J۾�č��Jd���9��Q���*>���7R���D��#֟����D��wȜ�5�����/�Oz*C�h����	��=� �.o)���?�b]��k�EH��l�C|7����M̈́/&m�|C7�~A&�/�#J9�7����Z��5�W^{S3z���m9�����1��R��cC#�"��@�`������ ��%$ 8��?x��=���`��?E�6Q�pt��Д7�V|���I�	�	�z\���N;���uޫ��,��J�	ѓ�|�123���*)�����uKBC�,�SXX\Q^_XTM�
�t#9����@���]	������T��u�R�����<r�LxX���ݕ��EbbcC��qΎƞ.�Vf Bcp���������DO+og��p�����o����`io����(��������%��/ $|ہ��g��1l|T��"���B��TXmK�x`�*"o��ř����ft�����l܁P�k�s� c;?S� '�X���S��.�բ��0D.��F�Yz�����H����"�d�
�-����%�z�t��kw�?p���e�f��r�޳*���-odIqLaJ���Y�C�#�g��:n��q���4m��i�M?mʤ�S&M�>i��ɓ�L�0iڸa�N�5a����11�ѩC������!ᥡb#@�a���`=������I�k��m����u9�IZ���v�T߹-����T�`0"v�� ��ʰ�R��1^p�w*'���G���6���l�X.�);h�Z��eyӅ{�w����­=�o.�}d���>��_K�~f��~��0eÑU���.oR"5jdե��G�kP� �*�N?[u�.E�Q��(�"��H���	�-$qD`;H~���τ�0�w�X��_"DCaq#$��Zr#�^M`�"$�kI���/�X��/&u��I�C'���<t,�<�'"���B�R�����5��	5��cqj��IZ|�1	9��k��GE4�O�(���Y}���#��{��Ryƺ�7q]�ϖL;8�X~��ckn�*�l�K���3B��4�E"�	��cǣ�j-r���0o���7�캙�����5�����oC��˥7s� 5���o����8���&3g���78}�̵��gƥd�%�&$%'&&&��&�F%�D�FGB"�o�u"���U��A�h�K'¤���ߪ7qNR$X�/B���n�k(���s�x9�z���s"��"��ƌ�H18e�д��3Rc�GI�z���V	��ı�NN�<<�=zTVZS[��3��������/�*=�DȥsX6�[�������8a�� ��`��7O+d4�a��i^nf���pԉ�,��8���X��w�P�O��WO�G�;Xy[�Fz9Gz��{�xz8�yn�{4u�����:���*@]H��W.�+K�7P��A5I �"8�y5��7��9u}���z�ݱpͮ��v�V�^��ȶ#W��~y�E����EuTaI��E#�pd�~ξ�$�.��D4WB�J�q�?����P/�!��r. ���С�����w���u�����>�|��4t�},]7'9=+=m���GJbZVj&089-#1%56)1&!)>!%))+5}hF��������&G��H�O�q���K9~��Qs	�O"���/�c#	�&y�N��&�ēX82D��7/�y6l̲�1+V�x\@mn}���EITgk֬9�kc}���͙s��������J����?b\��I�_=�hxXXy�����wFd����9i޸��^9b�_ꨠ�㓧,j�uj���=���j	�rQ� �O�|ۍrq>�#�y�o˩�U�����D������߆�/�8�<1�B��/�Y(h��G/B]d�{DحC��aiJ��J��k��Օ��:r9�YM�c�z"i��#�w�������|B����tS;�G��^9qh��y�W��u��� Bl;�1bG� �Q�q�"K�4�oľ���мEx��|�櫅G��Z�_���������~��e�V�B^Q�ޮi. ur�܁��\u���|2��kA�<���{��T�h.��(-���#D�w�7f;BV~u!eD~)��U�?{�]GN_�{���)��'�dDF�EE�DA	�
�
�P�O��.ªZPQG�h �4R�"��*S�쟷�fddJr*¬�Ќ�` <�mXf��y�SGv�5�ꪋ�e$B�K�	��1,%fxz¨��1CS�O�/�$Fn]����e���}�|t����ۙ3g��it�-c0%�D������EX\��q!�Xl*����_�gee����q��e.�P�?c�`3c'����.��L���N?�03>�]���&��䄬�h� �A�^�	a>a���n����Ƀ���4��40�)ZC��S��Mz@�`Q�U$Q%Q 52ji7���>qcŎ��l;�b۱�[�����vm���79��9u��*:g\�H��]YS7v���Q��g|9�N��1cp��l���P$�(���6�I�dHr�J([[�Hg��$*�Ag�����ngm����3�R�aZbRJBbj\BR\l|\T\|X`�WtJDHT�����{��K��ShqI�/���/�Q)vgD"jA�>M�2�642��NZ���������+��Z�<}��wWl>XPV{p�^jS�;q��ͨ3n�c�m8��lG���CF�%D�Eg����I�<*2u�od2T�1c &��r��t�Jw��pOR�V`T�Ʈ�9f��e�o���z,��B�w�ʹ{�O�x5��>f��G�O�p�/�+?C#	/��E��.�����{�)="�8�����(������2LE���^��b��z<~���{o�t���v�	q�	r� �bRL��KO;~l��WO�߾��Z�N��������\��S�O�w|��c��0$�#GZ�#4��R�����J>s:�&���C��N;R��V���lAh�݆��H;�P��r1|V�b�/뒼Gح���.V�W�W���-���y��X��dq+(�&AGu��p�[��>x�|���ѱ��\srtqurvwu�pq�rs���������������ؼ}WaIUU����.ԋ���FM�2|yl\搄���� ��)�&�q
�v��ܺ~Ť1C�"��C����#Q�Ct�FM�쑕�i��C{�._:������u׮]5�M"��OJ�]t~��W�/�g����"�3X B�3��y���mذt¸�@{;�����ؚ�
t�t�rs��w}\�/�M+�9�m��iQ �`g�H/�� �W/wgw/'�������%4e>Y^'z�������B����RF���CⅥ$IM^��Я�u��Cp!$���.m>pa�޳kw�Z��$����xR"|�_�_E*k��E���L���E�?m��.��_b���士B��D��Τ��]��B.(N�<�H$�.Y����k��*���U��ѷl\=n���������R�����]�"���cb��〄����������( >""&"<&:$2:0<�?4�/4:($"��#���{�����v#�ވ���?M�0x�� ,�g΁�7G;�)t�SZ��8p���JR�B��I_�4���pI���=��'��(uϷ:p���1��y�������#�IHbӢӢ�2�3C�2��|�F�])��T0�s����`�E���\�=���As�B?q�:y��m�V�A1e��-�i�Ml��-B���ߨG~�~M�!D'��c:���w_��x�X2�{���S�V���rdA� �K1���&f9���c�$���gl=i�������\[[�z��S�W�ryRW9s��R���o���rV!V� ��T����Z�[iB|�j��4X�6��X�A��(�|k��5���R��pD*�KxP��&�~��~�-z4�~�gn�G������"�;Ys��q��l�� �����s�.	����35h6��m�v���>�!AP���m���]�=�7nږ[XRQ��#B���\���E:n#�0&>sxZJj\�ഈԄ O���Ȉ`wGk�>�V��N��>qa��Ap�������
�
���w͊�udgf���?>�#6�+&�/*&hӦ-�L��N���/�O�'R@��\ՉݛW'Bԅd*����|�)��������rPs�ޠ@`��A�����]�@�htBE�n?���������Т��y'�~N��=�½=��E����>xr	U�����x��[%s��Xr���7x��t��S��N�?|;�ҋ�KO+k�2<rL��y ��;N��~R����߿`�^`���ێ^?}�ŭge�J�
j)�F��HF{G�S	���PX�:B���U��WA�
��B*"�ޅ`A�P��O��r�b[��Jy|_�7�H,��\�<�a�"�m]ߢ��P�y��+�̊[�x��'w۔�;5������Mdp *B��U�:��DEF��,BT��L��<�ohb4`(z�.�៽��ޅ B�@�p\����k}��e7�KĿ�k�L�y3��#*6���Y��[7�u�ڇ�76��u$��u�yg�ĥƤ���G�ǅ��E�󨄸X )>!rlBJTBjx|Zh|j J��5[�)�����H�|*�)%?B+R#��Z{�c��5�C�]yް�Ѝ��V��IW���W駝�(����G
�&B
�/��Q��w"@�@iiSE����ST_XK�QH��u����7|�|�¢B�Ș��(���#F�X4wε�j+*�Ln�������w+Do�**���-�8{������_{U�j������,Qu$J��Y�nS�Zѭ��*�[��K���Vv*�;��-�U�Uk:4���v��P4w R-�X��O�D�]B�{ (TM�B�vĸ��6m�~��un�����B 466�?���������������� ݜa;GT������ju�Ϫ&�A�C�FƤNJL���"��[�Z0�������?�`Lj��@�� 7a����Yok'��D",+�R����2�����������/)e��?H9Pq�i,�_"t�����2���Ơ��y3#h�࿰ w/Wk@�}��}],��fc:���y?tB������q��E��}�ڵ"t�J����w�icݫ/�=�8�UsҼ��w^_t�ޑ�UG�,�{����yS�2z���]�v���}g��,x|����C��_Ⱦ�S����M�`A��) C�b�iLt0!�%ԭ*������BKiН��jݐ}t�[(�eb�B.Ӫ�-�\��H"�L����?��P �psKN��p���v��.�\@f%�N������j���f������0%6D��
E-�F����D��j�

�ws���u74q�� �Ck���4��Mx
�@��x"�@�(t}j"��SY��H��R@ξV@����c�ʸy�x=}�[O޾��չ#�
�-~p8�Α;7{Y�2q���/ܓҢR��S⃓�C�� %1:9!*%!6%!>111.!)*19,>1%y⼥y�س�ro�O��be�ELź�K��H���.yږB������k',�1c�n,WU�����,�C���2��"ԯu����D(��D�D�d�S9��",��u�/Sڤ��i�V9�B���j�Z���'�pwo��а��P <2:8$�x���Çd"��Gp��䗥�G���.a�Yr���r�����55�9�s��94d��l�d�� *��E*k�*=-*u�R���E�֪ ZZ�ͭJ-ЦҶ��-Z�ժ������E�mtR|@НCTU�T��5v�[=FE�`�������y�޽Mѩ�&F���.elܯ_�FƐ�||7oݞ_\^U�ы�G����\�eT�d!c7�Y�����:,365!�������֢���>������=���q�~p�r�D�^����(t��>�f��^��>���KK��1�������J�������iU ��r!XP��f�H$E�A�VV����Q!�&��m}�E�hm�ݒ�O�q�3C�����v���Y_h�yٙ�X��;zy��y���&���S��|�$y�ѫ���ٿ�!���G���~��^--��^)L���Q����v��K��｜����������s�꣣���\zp��Sw^�xQ���ZI������UdA5E�PEt������C��M(�s��.
����6��+~��%J�A��Ax9�r�=D����چ�L#�'�It.W.�$�LͲ2�nߺ��Cǧ��|&a�	���"�^;!R52�R�vs�vr����
�	����	����
�aD$*�7WC�{�/뛈XB4�Mx�@�_O$�wb1)LtC8,`�';����������z٪�s=���n�W?l�ɍ'�]��sp��['��:�����K��?���u򺥷�S�#�@~ai�!P�i��@zbTZB$Q#&�&�	1>2.>TGXbJ�y�MA��)�/]_�m܄9� ���0iu	�u��C���K�_S�����'���
<���yb*W�}�M�h{E�d�6⟋��)�\t�T����+^/XP?j䧻�J��b�5��aAi}��@Ai������rLi���R�c��]����<�ً;o�v��g�h���]P�gf���B�.)*�Š�Cw�EѦSwh)3\�9rv_a�R���[��7���s��Өe�D�Q�5r�J*GE�R�9�,S��5�Ju�B�V��M�lՠ;4���vkR7��V��j�6t/{5���T�&ѴB
��J�o!wJ՝J�۱gB"|��M~Aټ��|}����-���ӯO/tg��
�������o˶�����8X���	��Ta� ��1��03!.5>bHz,�m@�P�������bo��n��!J��"��w���q/W��h��_�`Tt��Mۊ�k�T�"��`�_"�U�^�w"*�Ƽ�rhGCš�î���V[ۻ��Z��{xy����;;:��m�_�%��qoW�Wy>.�^���.���N�ƽѽ̠gm�����������W��u�ޯ�{E�N_5��ϔ�ɫ/�������Ԅ=�����r���Ζ�<1�����	O^��z��ʽ���ח�__z��\���UO*�����x��&z�����\F�T�E�4a-�QQ����	RXA7�^A� �@C6W14�.��Ѡ�r�����U����G��x���5�T�WՀ�?zV�_�eB0��J��d�z��Q�H���B"c�ܻ�kߖ�k��{��ל�xl��v�\l�b���cc���C�}=�B�|���bCbP�\��&���0d1������ةs𷫨���4i$��'�Id�I�1��2�t�N`��6���ӹhC�3����۲�T��������ȶ;U>�-9�f��[o=9�k��;'.��z?��ӏ=/r��e�Ê����Hߔ�д�����2�#��FL�A]�~�V��e2]��n������z��ƫ`H�n;4yն��aĭO�q;N]��r^�"	UMt�!����D�ƣC�t�
`��p��dT�T?k���^,�d��F]P�,A�l$����+�¼.�yYP���
�s� ��'�e��~�5=�g�K��w�yۇ���K�.]�z���y��1��?666(((,-QQ���2D]8sR)�5�D�y�@�.���>��z�q�x�1�O۽j��Ii�Fg�dy�jI]}���,E��W˕Z�\)�H%2�JZT��2�D��)[4�Z��ݻw���jC-hO��+Z�-�ځ�w��f	[$ JT_E��bU_�����/T���Ri�`�BU˗�S,_��En%4� R@��-X�����ohd���SO���c��������DXQ��El����y�����cR�b�M285��)�V�����,��U��hMjhX�:�8����Ǆx'EBF�u�����
� ��ё�A�~NN�,�v�ܟWTE s�4!�P��&�K���,?��QQ�-B�;����Aa��kz�8x���xx���;9����چ����[���;���\�@~>��^.��M�� B��NF�vѩ�ޞ^~��A���7��$Lپ��H��P��1�����W�^
��Ţ�);�s��I����ۍ6��]�\|Xv�����:y���+��\?x���s77^{^u�SH��/%eWҟ4p�5	_`%9u��u�b"��̩��	�R�<M��Dʒ��J���֤��g��:q��=��Λ��$O�:j�����ŹĆ**�I���y����#[7n�("�T�x׬^�q��t&���.��S[Ohx��3m����\2k��~�ζ�>n�Iq�)	�q�`8_ww�@h�F���%ƅ���B�}�|!�����:����H�pE��McS˫��*��E	�Ji�`�k1��d2���37� ~ta]Y���fq����X̾G�x�R1w������8s�����c��=��`���}֎���2RBB\Ғ���_��̔X=�����p�����s9n�ZlW&}Z��STt�ѣ�w\�yy���Z����0�;Y��)��H��� �@A���������!�L�`��pd�L�A9jD�XW�uC���1�X:���m�p��:�@��ut'�R;DV�^��Ucн)��
�#=���U�2?~G-Y:}�t����ǽ��A���z�mmm�m�/^��2�Y&��$�1!M����9iϽ���՛w��9��쎅�'L�����]����g��[�HՊ��/�H�h7�H��4B��/VHT-��>�d*yk�H�J�J�Z���[A{S�B�(��
姯L�w���!�>���·]���w��7A3������ᓗ��v�e	�e	f��A�)��~}�A|����#��ݯ_?812�����+1�j��,���)q�w@TJltFRlfr<zL�u�.t��lg
"�t���jI�	���	���
tq��m��m?���_�QTZ�%�Ɍ���/�*���9"�����WRI狉,���iiy�7 ��7T'� ����146��p�u�ww�u�Eq��qa��K������a��Dhi���z���5<?��7(,��?�/u\v����-׳I�^��=g}}���T����f�l�(r�އ����1�w���1zǥ����eWn�<y���7����]�w�v�!)K�Ŏڼp����O�O�9t����K�l�ҭ���}�_٢[5MC�(	L�]eM�B���$H��Sw�H��|Ivܨ��^)}s���ie������wwo�4m�׹<&D��7KĚ���l�J�A�?����8a����Ջ�L�������������n���"�c||HQ/B 8��������͸��V��'��'/�طm��eK��Y�rΕK������"��Cd3pl����|��#�p����b�vΞ[�ri�d��s�����~�֓�W���9�u�?tm=~�FY����;^7EI
pHO��e��f��g�& Y�����x=�)	�	�49n�!O&~V���0�qA��;w��?��E��Z-E�y�H(��*h��+��
@�Ct�;*_�"��Z�P��P���� L��tܓ@N��;�-ŰetQUPC���u���r�M���^ZO*�#U����
�WP�����͛�:H�9o���y�y灍[w�9p8<2:kȰ����F�����IlL�������ıc.�>���Y�����O��9v�����٧�Om�~�̅
����.S�_��w���.��S��E��9��H���yTX�h.�䗐���H��>����q.�8�Wt&��>�B�B��*N<ݫ}�5�f=�����y�KE�k%��oX��N$k�ΙN_xRs�v~��E�1Cl=C��X������Ѿ�zD���%B�_�
,o"�Qp�R��w�*��aV��11���I�w���t�5uw2�p��n��e���������� ow'WG'GԂ@pppDDT\lBBb�ӗye5H��F��/�*�������EȓhIt�-{�� B/�n��7�����r�r�8�_D8��A_�-��7������m��0�a���J������}Ժ����{��x[:m�͸Y;�����\�?��5�ԉgr�TR�A�_w+��ڝW��>����ՇO/g�Ge��������Go��37?���������W�_-�p5w��#���'�.n"�UU!�!���s"L���k���5�|f��}��g�
�&Oz���{�v߹��Υ�w.yt���C��Ϝt��6�!���]o��%[�n̤R��"��H�a��=�)|����%�F&ǆƆ���z���S6��}�c����v�00����b��M��[����L#pl����S6n__Y[�֊�\���{.��K�֨[$���uXK��Ow���$��K������۩�ԍ
�Bq���+�P�#��Mz���G?��뾶K
-�${�kwf�"�ޅ@�,��*Q�ŭ n9�hށ;����S�\^�Kɴ�o?/�*~�i@^RW�@��l呼W�w�~���ᗜ�OL�LJ�赗���O�%%��ŃtD�a�F���ಏ�=͖K~����#��M�8A��-I"Vҵm�rMW\���HR�R�0TY;�my�>���)��zy���"���*;�
�x�@�-Pu~����V(Q�I�����Da��fOh� uLy]RMWӄ5���j��Z��
ﬣ�����«�� \҅�ו�GN_�;)=s��M[��^7m�, +[P~aTL��s�O�t�T�FѡU477�������X�кn\<�������#��|]��0i�uN�����Ү���/���^4pn=J׾�Cվ�����B���v�z���݌���r�X;��~o�=�\|�H�n���I����B�ؘ7�쳫�vԌ��v����0|�����5�A#���X�۹���_�$OvJ���Z���+p�c��F�Æ�0�rCx�H�næ��Z�L=��OV��et%2k�"���1."�"��E�`������b��h�lo�hc��`��n�p���2��0vt�ҋ��FFDD�����������H��x�"�)����E=T�7�%j� �R����+�lغ72&ed�X7o;k� �@;k;G{'WG7���������w����;���	��hm[�l�����94����������?�I��n��p^�Q��_-���q�`'�A�)崕�ۊi*p�("I�/ʩ���>)�z�i��@�W�`fO�?z��g��|�I���~0�a`�FԼ�+s�b������۞�d˝��
*\���o"dIZ�C��V><f|�{-�MOYy���5�E����wrw�]ޔwi��K�^=t/����˧�N+|�@!�dR�BB���S��)�J���4�J�Up�26K�bI8�1aIY�V��!�8C"C�p��`$:�'$�/\��� "��� ,��x�;�oܼ����×��7]J��A��K��{x�ͣv�uk��9s��F���ӧe��T��"�REp�e�DI�k@��tLZs�j��X�$�A�u�ٸ��F�8~�qɵˇ�$7�ݸ��.F�_��Fa��Č�` ����Ĥ(@Rr 9%V���`RR���'��)���C�n���w�^����˛�rW��kmU�y���-��O�,��P+T֋�d�DE'Q��(j�&�:H�Q�;q��<��O��N(���U�p��0���z���N���"�$�;��7	�m �����c��+6T�Ā
���"���jh
�j��������%u��E�����ٴ���;
����ν�޾ �\�		���#��|����Ё}/�?˯,.x��P�r�uc1�w�����;�:���=�.�^113���;/�ݩ+����u�-(��%=�n�����'0m��|Z��'ĥg�7B�}�S��9[�4�ȭ�5�W���^��D�;h�%Ҫ;r�'�*=��
�y<"���!���Z����\��m�0)ӜPq���V.�֎n��Ύ�N��z@W������������u55M�F��:��(<
��ԋ�/{e�ȥ��N G:��9�� l���'�a.6���&.6Ʈ����í�l̇:X��m��mM�V&Vf��M��E����Ď3fҔi/
J���@�R�p*�)��E�MT�)�}�Ĭ�Kǎ��`못(b`ife��`�h���P���C���CKC����	�
ϣ0b`>���t������CR'<%H7�_���d9�\1I\�T������f��8������$�+|@y�����������_�Dx=��ռ�W�M���!uƾ؉;�^�}Ax��u�=Z�̃�/T�؜{�VY*7u��*F]NdkX��-�a���aS`��}��$�J"u�Ĕ�������� t����{���=ul܅��Q�Z+HZ4:���A�_��h�b�D���\��>� \.E'BLx(�`hxH ,�â�#�(�ÿ�00����|Ӗ=}-�?���)4���n�_<��ã�"�u���=+����nK'B�DFկ�"UQ�Z����ڣ�֜/��@�v�)�3fΡ�[n��~5����ËE��޺1b�b������,?VH������� .����_�$Q�/�q��΅y��̜�y��>~v��jө��fm;c��;��jq��+��aA�z��~�}�~�kީ���}�Hl�P3����a˺�Rr`A�@�Q���A�U/�v��;��p� xkհ���J���.����i"�=��(*(*����Ʃ�¡P� \���r�q�ͼ'y�_�**VP�������(tHtl"�~aD���͉cG�dBe�҂g�N�z\P��ؕGE��u�ߖmڳu��k�Z=+)�fˮR���s������^�߅}����J���')����b��r��_tb}>�"�m���q{o�k��[.O�V�4�2�J���5��и/26?[}���&���mi��yǮ><Bk.�M����%��?j��^��{)f�\��$��Xߠ� 46X�?��
@���Z(.l��-�7PO��EXZK��GH`�0]�P�Ǭ������26�������:;��x8��,h�de�fg��rFy��"�p(@X�_`�{��k��{P�g�I{��Y�3@z{d�1e����ץ�UM���đ0~��۟?�l?^�i �.�֍�2
��EMT�����l߻b��P���=\.���^(/w_7o7���no�A�`onh5� `���t,�PA�ٓ�FN{T�-�*��$QU� "s��q
$<�!n��(pu�z"�������Һ'��w��}~�~�������"�g�<�w���:{m֒m�i��g�o[V_���?2y���R[㦯�Z��myO����:�����K�ӧ�Rގ_r�t�౗¤����<�3*���u��,˃]���5���<�{���gM�D��}�Eӭ�B�,רdj�T%+�ɓ0�bW�M��@�����`@hX��aQ�P`�)B�pq�غu%ᇏ����
� (pޢY?�������.��K5�|��C��h29M�D�LMS����`^%o�����[F.;���m�~y%\z�^A=�嫛�U�?���9�ٗu�k�zR�r�����E��G�������gΙ?[�Q�76�\��G��>���������}�r�s�V�{R��ĵ"N��j�3JK	o��5i�F����#�"A:P��!J�H�^��-�!��uȀ����{I�^��P/���V� z�p[�٭��r���./cHK�r����*�4À:,B
ki�� ��R8�lb$:�ɓ�����=T1>)���E��E ����9ݻs���G��|r������=)�u��KF��H��惧��uzך��VM�I=yV������@~���`+��
"����Y�ˣ3E�Ţ��?@�^H|睜r�)r�#���+�{z۝�7s��^)��������֤��v�6�ZQ"nnj�K�����������L���5{���Ǐ_{��ȕ����`�C�X|$6�		�`�3D�Z-8�næF���\VM����E�5Z��b'n����IA>�(�;����n���q���@'[c�B=h��������l�z�.֎�&v�C<ݜ㣣222ʫ��),K�S�����������	�)�;H�G��؝��fg�`:�X���������������t�������7;W[Sa�֗8� G cS'-X�3�~��	/4�/@�&$�EA) �/�t.�He(�&���T5P���U?|^v+��ƣ�+^_{R�4i��='�7q��~�:~����Yc�O_y|mn�g��	kǮ=?}uIH��$mL������#d�'.�����:��
:���`��s��Ȋ�sE��ݽ����w��>�k�����(>M0���I�5k;uWG�5�m!_��
�t.�K���AX���6�"ts�ڶm5�=`+W��>�9w����Gu��ޝ��_I�U��!B<-]KU�4�{����?�=Ѕ��ܒf��=mlyA}�}T&Q���V�`����v�ғ7Ll̓���"���ްi#������#b2'L�u�lp\����.Z;z��Wɪ#7�l����H�S6_�����
=��Xt��9P���\| m���.p�!��3��E��) L���X�(�o���j%U��J�@����a%����^�j-c4�2��y1]RJ��R����0�!H��48��xr�B�Y��0epk	ԣ��?�zt|J.
�'��1@��u5�9��KfO/|����gE��V&->x�Nr-���y��.ݽpx���Q��S�_�Q�p(��
хB��'F�?�[�b~���h����[�;��¢'�-�^���*������̣Cתo�ZQ?��YՕ=w����>�T��!����yۖn<q��ˣ�o�����@��C�htH��(�?�6?pa\�	�	A�1��l�i �xi���i��æn_�˳���$�G��"� <�7��p�I�;{dߍK��OR���]R,���x|r^?>+-9:�L���6q���l[���C�Fe��m$�Se�R B:_W����x�&����P����	�"*�D:s񊕸�GG�i�3&OO�Oq���0��fo�p���������޸��ѽc3R�B�}�B}]R�����(/W��IH�z�l��UO�XumKJ`ip�z��gs\�l�LLx��I�2�ȴz ����yQ��y��o=.������5�/�<�w�5�|^�S��_}����j���׋5��jD�V���E��%�IZ�5�ee���2\e�@��o~�>��sA����6s[�K�j��aQ�;W������s[�]_Ut���cc�����X@�� �ë�k����Cw��}�Z:|��XD��7u�T+K�'�։v�w�9d&02< �ć����� ��h>��ҋ0���y����mo���C{w,&6���z�e�D&Rh;�kV�ނӟ��tB���w*e�����Q�
߳�_���TFk%��������B�W��ǩ�ո舤ؘؐ������:�Q���������𨰰|Rj�D)��x~6���;7��ݸ� �x��đcN��M=c���S��^������˗��j���Ќ��v� ����ѣ6�k�=�1��Cr��ȣÏHu�_)�_(�� �$7^5�U�X-��n��ܤ�|��w��q�1���yF���CW����o��Ur�v��/�8O�y��??z�|��{�w\<|�~A�P�BX��:;�\)8�R�����:{�fJ�>&$<&,
^y569gnmw���G�۶����L:����t���f��k���w^�	(��OnoZ�",6��Y���v}����Ώ����Ӗ���T�j��U�V�bt@�~�>�Yz����t�ޢ��j�ޢ�W���;o���J��.��8���1r���wN�A[������w�������v��ջ���Y����Cb@�F�

�`�:��[=k7T��j+j��P�@"���ۚ0g���/&O[��$�B���[���y�������֔� �L��J�dg$�+1�&E�Ecɍ�oz�;��K�c<C�;N�
�A^g��y���gaޟ�߶EXW��"hT
�=u�Lwww\��/纚[��y�ԩ�H7���~�m��l�
�w��Q^�nKX�ӇvM����l��I��=]=\\|��o=0a��
��Q�D���"��*�C������z
��ªl�U����{Z��Uu޳�u�N=������O����l��N�>r���g5ǯ柽��΋J���"P1D�*N�N4�W�Iv�x!������~]����JnI"^�j�����Y��S�"�|��~�k+z�?iL֮��,^wgOg[�@ �t1����
8��N�7�Ԗ�*�/)~F��kԢ�w����N6�(,lAX�O�a\$:6�/"�B�m߾�����ޞf��w/����S����[��������D(Q~�@�|QԴ��*�g��S��v�l����v�Z���ݩTl=�5��(o���Ux�����V��ۙg��o��}{���}�΂���;:ڻ{Z�ûz�-[5���7�dNX�b�Y+��u�½��������A�6���S��'�-�:w�-��k��Tz�yGȧU)Q��=iO_{xǙ�$��
<�j��{�1K�ɚ��[��P�V�΢7_�Z�\|�<sK��UQ�VD�_5a��;/n�R'm�$-
��;}��M�n��Q��$N��υ�k޷�(�n�?x�\L�H[W/G7_O?�/��	�{������T��>Q[���d�6.�vf,�s�^��Ua���wO�۲y���+7��YuT��M��NxuP�J��Aq���ǅw�j��k�}CH��5���:�Zt��r��|���c��M�?�w���.�SN��4��V�	�N߬w@LU���S��/m隳h����n�}u�ы�s`�����cq�L�PLpȷ¼�2LA!@�U��ڦ�Z�����,C��k�Zqj֖��i��cb�X�@=O��P�����A�m�?�D���.L��L�5"IaT8&>W�<�S+�ъ�8��q�&prh`��\xF�.��S�?�j�D�	��X�Ě@�W �@��˟�.@����aΝ:-dq�4څ�f!��=]��q^t�	��a�8�����C;f�� "�w6G�ۀD������Ϝ<?g��~k9KS�R�R�rWJ��K��-��fK�Lȋ���>�]^K�72��2E�:�?|^��e��g%����9S�[��8>gRZpl��	3��_v�|;�ܰa�ޚF*8���J�H�%��;�r�*ƈ){�_�lw�l��8�|��eTʸ�9O�j���&>�
<������gϝ��.���hk��?|�����O�>���5�C߹ksB|���ˋ�7�D�� �z��s�p�p�  �aX����a�{Ǻ~��w���Z��s�ޕ9��(w�ܽ�B,˨l	�&�E�J�_ɏ��^�;S������C:kUsP�Q[��)ۓ'l "l�N\�L��{��S�v���X]�׳O+qQQ�L��������F�b���"���9}�T%[�l���7�ݺ}����[w��]t�ʭ��
��XVI���U���SWK�����s����?����ڸ�F��M7�*8����l!���ѡG�*��7�^�q�t�ڣ����jE�/H�)�O-?�W�����\1�T��L����r	w�/���Kxe�>���mwk��#�6��ۡRb��*F%�_���08�4.!� p!x�D�W�\����ЩqS�y��>h�Hx .:$2����Z
/����cEO��.�z�����^Q5Gցw���=���1���I���g��:A�Wi�{`>E{����;�6x����������]���-���tm?I��A�Ki��������~��~�t}R}�do~o����Lz��(h�m}���?E�e����
��_͚?�
�o�8�F�|PH����{(o$j��ե����k�"���׫�i���@��ܶi[�%�؁�De%$&aC��52+&�z���-�Oܱc�����p�/��΅���I�zF$��C�+�̺q�D����	 ������5X
_>�?E������DȂ��&B�*�m�l--������_j���]�����hm�����h��r���׃й���}vr��I�c3�R#�C��C��#�0^N "������iS�V��_e�*����n�h\-��B��-�'	������%�j<嫤�󲚚_�x_'��W�O_��x�z\NΞmO��޿e��K'de�:|x��9wo޸z9w��g�_��T�AbpY"C,ӕ�SQEJ�o��[���)S�m�kJ۔��^�		#�6�Yp�̑�Gw�.zr���};6N�0���B���c��7;gd�KO�<y��8�l&u떵@aXT���_?�;��C�hk;3\D06<��-�O"��E���{�9�y;�ٵ�������D̺u��ٓ��ݠ�z��o�d��D��N~�P2!���Vƌ�Ԩ����(����^פ��U(�&o��6v�J��W����x$�P����"|�ꦖ�矖FF�D�+����;n޾��B�h�֍i�#2��3�F�e��<s^a<�w�5 f�[�l����b��ܓ�o������﹕����-�	s�n�RV�{;f�/�hё��	�V���Q�������L�Y��"�?>��#�ݨ��.丧.8��V�>e�FN�ݠ�w�1x̚��땢땼��Ly��/~��یF.��R���O�B��DXCf���-�x���=G�l�{lԤ�c��7sޤ9��-\~�|�\��05*�B�}�����͗7s��T� ��{���Ew�z�]�V�e���nH�w��!О��[���l�zA"��tt��������Q(������_�_~S��*� �$�,�z�4�v|w�"�tA�6���C��^��P��3kѶ��Nݺ�����9�`:9;88ع8:��� �\=.>^^�������nOOo������^�V�(*��!��R �E��m�ꗠ�������T<.14X/�츨P/w4�0�����..�t�"EE�@_08.2���#w;w��0�y2�Lˉ@y!=fΙ]V�H�A7���j<�H�ͩkh"��\\����W��X쪚:gW333l&5!!<4�������������������uGCw������� �d6���������ww�F��y���m�#_3�e���g�[u8gѮŻ.Rԟ s6�r���jAO��w��{�<�QHL��dʪ=�3W.�y�q%�Y�Ƴʧ夂*��/w�=�t�5�&?�q2�w��KgϚ<jtfrfZ���g�\��k׮�O�+U����lx��b+t��*��۹�֧�9+/�Ő���m�Q�h�#��ՙ���o\utǖK�޺x���3�Ο^�`���k���)d����ܿ����&��?�-ͪ���%ł_������_?|x���cem<����a @��r�:t"�¡�IA/B_�}�7�5�D��ۗgϞt������6ɇ7�������Ǣ�h���2�2>E.���D*����a���ʡn���V*Fe�!�@�.���w�fM���t�W�*��>A�>�l)�#y:�-���2)k$ȯ�x<lW��d�������� oGg'@|J�\�h�j[�jو�����&L�:eƜ��VܸO��x��}gv�]��p�놕�~I���8.,k�_�^y�X�m�v��z���Y/�[u�z¤U �W	z�3��_%�u��"2��Zs��-�'k�����.��Ցs���Zg���>~�ܣ�_	?��-���曹�7s	r�d֌��~yV1vKd�lҺ��[���@%Ke�A*|y#KR�5�ED&|����.�,��{���U��.Y;e��i�W�Z�z��sWm\�a۝G�J*K;:5���6uW�|�w������^�4�s>-(i�*�v�Ԇf,ZE������n@��8������}�%�Emw���[�ӭ��P�:�}���ny_���_�7(�}+�}/�݈;>J��t�D��R���w��ވ�{g.ܺf��y%���_neeebbbinaka�hc�lo���������f��#������%+J*�K�ʫ	 `A
k`6�Du,M�����31�#bcGDE��b�
�B��8X[1p43�s�� C��dX�?!� �Ø0غ9XZ�X�ܭc1�H��x�b B"S@��E��g���DX��"dsyյ�...���(�:(����hm�le�_��MW���YAoN�����^��Cl���\,�=�~�[`xHƔgd��}W1cV|�p�)9n��E��ݨ���/���!����ݽ�������*f⊭g��"e�Qs�EM��V]TXI�z���I�w-�s�dP�Ӹ1IS&��5k����ƌ�|������\q����),>] ���ߔ��
�\�Ӷ����7��:��P�u��T�r��C;Ν�r���KnZ�tł9{�mY�`����*�ʛ5Z����_��۷owv�w�i�<֦u+��dL�8�Փ��fy�Z&��A�& Z���[
��	t�WƄ����p/���v|aG�R,b޾ui�̉�.�"�j���S>����}<FyK+�G�ټ[�J��V�>�����瞳B�n�&Bzϩ[U��S%�9�5m��Á|Z��=ۯ��[������wq���������f���b`BrRb
�� ̭,�ZX���a<v(%3mD���Q�F�����x��+6F��ʜ8k��E1��:s���b2W��tD���Z��^�BV�pZ�j�@-� ~�{��@U�D]��Fn��s�v���;ʨ��֮<�_*�r�؂��i�C��K��+N;'/����� �{HB欹��~���Av� *�v\|M�\��΋���%M�F��(���E�K��|%��d�,�����8"�Dŗ��\XQO-�%T7��%5R�H�R"���Sw�h��Z�4��6e��| ������|��r^-��PSYQ��ܹs���`kG-�!���_E�����h��� tR���T=���AU�[U7�B��듼달����W����띬�O��N��?}��U�N�~P��Iɜ��#��l��͌M̍�̌��56naf$ie�����t�ʲ��Ⲛ��F@y\�P/�F�����W\LjT8H�#�qz�;��4�!� �\�!�_4> "�=lC BK���="����Ui"[�S�?E�?�E�a��#z��/�,�!� ��Z�9��{� �L�ؘw�6q�3G8Y{��x������ ��f�2&�=��!��P�(`M���?.t��˅T�����U-P��X.�y���g���;��|�W�������7��gm>����k>�.$��g��VN?)#��%�Ի�^�c"�/�6o�<[�mdJ$.���(��#��:�i�Σ�����r�z��PBI�h�f�f�Iq��.�r/��E��*�ٵ}ۆ�WoX�|�%��,<vh?������!�A�V(;v������-(x��(r�+�7�_�c��Kg�ݿ�{��),�������E�D�F�^��[�F����~��^�:�߳�M˧�]�m
��q��ř3��r�(�R��_��.z����]��.�LD�˘2�T����
�������H��]1e'��Y��:}�,}�Z��3S��_���u��#F!�Q�Iz��3��?~�ԑ�Ǣbc"c�c�� �@��ii�#3���� Y9��Y�iݫ₪ڊ;y�ٿzݪ1cFEEEa����i�ə��ؠ����tD0n���d�B5�A����/�������+��;��R"K.҂��Y�g�r�,�$�ڈ�
�����`Ϟ���G��Y&���q�F\^ �X��ΔJ��_�w����곯P9���P����:�jE��>2~Y�yS�-edz5��(x�?E��c� �y�k��!�'���1e�e_�$���{�@VS�j4=uO���d ��|����+J��㗫	5�Ϯ^�9q�b��ͬ�Ǿ�Po�)¶�~��^�m��k��t��v�m�|�v~��������.x��?E�Q�=���$h��p;�Ge���Z�ccgkjj
�gd8d��o(�10�5+��DX/:Z�D�'1��
�a�4�3c#�b"�������{�!n�&@���]�z��F��^�a�kt0|�
u"�-�S�?�j�N�L�?D��*���]a��Y�w���)>5|����0Kc;C+cg[KwG BW�H��N�������ps���-��`b�n=���������芰��������bX�5�����,�y���{D֚�e�Q+�^-f�ە;i���W
s�m���P@���_=r�������x�����²�{�Q��(?+��0;KlRl�sg��5#c̘qӧeO�4}��m�VIT&�/P �:�����P(يn�jb�e�{��V~�G���l�O��߽v�_N:�����Νy��)P�J�R�U���{��^�Z_U��ww��T���8y��Ƶ+fM�0q�ht0������gA`;���V/B������/#��������Z�>���3��;q��M�������­��� B�w6��<)�E%M�S)�|�f��\7cg���BU܎S��Ҧ�&��Ӵ�{	.Ih=��#�A���_W1hiyu]qiyt\�^�q	�1���ؤ��䔄�d�]�:\�Ǝ���vq���4rr����bSSS��G�%ǧ��'$�f�D���]��E[[�
���GQw�������ki�(�����4���$h�K�V���)�s���N �ݱ~۹䬅kv�6��\+�d,�=q�Ƀy�[.��Y�>g��ܴ�{����>�`͉�5'o�;y�L~�3/ nf5�]I}']����;q���mۗmݹt����w.\�D�+�/Y���XOI�J�@�-�׼��/ei�8-���&QA���� ��U���M
�"�D�P�����+r�̕[��RfO�g��U�7E%d]�V�"w�o"���٥j���#��ʞ������h���"���.B8v���B����@�~ڢ�+7�������c�#�A41nf2��x����ե�y�}�K�-/��y]ZY^ݨ�PO�h�EXCd�RX�4Ѩ�'<���'F�ӣ� �G�q}�n`g6���&B
���'�<���L���1X��PO���E�W�V@���������_�#�2�p9S��e��&��Kh�`��hNdAh?��p1BS#؂@�nvV�v�>.ξ�~n ��G��������P�a�Zk6F�lz����0�=�����2�徦{��{��&�2�ȓ�.�'m�G���u��v��R�����O�-����z���`��xD ��?������G�p�e���޺u����W��fe����-8�{�v����]���`7�XD��!U�&�����LI'8�QDj�����6�D$���¢�W������⊊���Z�,���R�ΜR�I� �X,�˥�
i��K"6�~q���U��E�Š�1�vV �8+  ;:����1v��aQ�!�`�������۞ݛ��Z߿�n�Jy\ʕk�L!��o `@��_��e���R��,H�l��%W��j�d���2�o;6bN��-�jU���?U��.>�
ϞEV��h>��,J��#u9�F��A�����r8Bm�Q^Y���������6g�\�Ñ�Y�	q�qQ)i�Ow}�{kO���/�����
.Y�Ff�'D��&''���3v\����28��Qk�]�->3�����P15m,u���G�����ז�wRy�L���� ��ry���JS�����^�� �J��na�ǈ�)�^8�0{�('T�Sp�Kh",�4�154e�wx�:4m��[���eL^�(g����cG���LE��#P���P�@�:�3 ��;���7-g,!M�����EM�I�~�tp��#�mJ��6qҦݗ������ųW�eL8YP��̹1qՃ9�'�~��	�8EHx�ʊ�,Z�|��M�����Q-��!xY[:����v�Ը�����|�����A��_��B���$��-�"T��!h��m���qZ>�T����퇉�v��{��K�S�Daí���t"41jfnllhh8L_�P/�$����& �`e#���\C��P�%4aʒ}.QcQ�a����수�Ę�	��V^�֞N���pOZ7�@�p?pa$60!
�\��t��1q�6��E���w�ñAqG�_*�&�R�ML*["�)�7�@��#��i\~��	�wq�w�	&��p�BSk���������>.�(O/���/���twv��t�0�2�1bkl�jc��q���utq�F'��U�K]�w�W�}%�߯Ԩ,�'U�!�Q��7�����w�p�������� 7�@w�pV�@� z"1�~ho$���	[�a��WMD2��xUTz�A��'�J+�Ӭ'Q�h2�O��u���p�>��DȐ(�2 �PEJ
���U�"�WRQYZ4PUS�*��d��\W�	[(��
�t�
��H��<��Cg�I��EE�����X�@0ڋơb���| ��F������^���>�:n��k"�j�l5�ʹ�SƂD��P�|��j�ܸ|���3��2�Z$�I�p�Us�Z��Y,k��$�<8u��هUOJb����7u��*i{�����b�����?����B�񻅧H:��x�Z�X��<y�`z��ӧg���iok���ss�	���������i��cH�[D�������`B+�!�NV��nn.>H?TpP`pH.28,64*!8:�
$���+�e��"�0�-t<�S��G���e_߯G_H�Ό�
uhbLTFb\����!����)ii�9���S��8�����zN����$.���۸���5>���7!3)"9�nc`�8���������t��Nn�ow{����GpDL�ϖ�1���&�`����}�s�S	�(y���5��.sh
�½���cG��m����/{<a�c�Z�~���-���[�i͢{5}S7�E�sဦ�E����iT��Xmo�����V�Cm��KGÔ��u|�x�wt場iU��!v�a��>h��s�w^���x�E��E�"�]����`����a���0���Ǐ"��#��)�J"��L+��W�c���CS"&�1ad�ɣ��(�4���~� �����`Ѿ�,B�W�Bk�VaXߐ���%GF��}����RO%X?E�S��[���'8RC(�$p�؅R"��Kg̙���i�����|��͌M`�Y��;�x9�=yzyzx��<�|����������D����k���<�O	��GL݀�^;k{�G���*>�O[��^�m�t�y::���_�����7��>h�@X�~h?���Y�l���'�O��D�^�D��i�'Ph,.��ы(�[�Ȃo��.�ǎ�g�:[��.���K���g�7�����`�F�1>���<�<�HER�XoEb!_�������f'ffť�� ����/D��b�!h�PT�@�A__w_?Į��z�:߾�Ui$L���&��h���M���:�m���-*�Zb����p��<E�P��)ۚ�̓\� �����b^w���R�]�謔jT�mA�Bh�6��
Y�BB�K�
1E!�ɅL�PѮ9y�4Y9�sg����N���Q�����ǹ�k^<Xr�B�ËO���-|p�������ٲf��̴��(ХG����#ä�̤������9��I�$��E=��l0���H����rރ'%�w�2n��N��XtDfrΤ�ӳҲ�ܼ��ب�KW_8{iH�@�������D�+������������M�/���A@ "8���Y��P3�!��V�.���v�ђ.�np�K{'S;{{�Z
K���o�%�ۉ��&E/A�6mƆ�'���zƆ�����B�f�����}���k�M�M��1�@�_�z������}h��}ۖ�;X+��Y�����K��^�} ��<U_;I�u�i}��پ�&�lϽ\�B���柺S��;�w�a����_�TQc���,N��a��7)�~hΚ3�<u���;Eg-G��ں�Y��513066>�Mh
�B8��E�@-[�����������H*=��D��RKh|�ԵƁ��޾X���#��Ã��@��p�����[o7[ �x�X|=��H�`����M�<�l��m�^�� ��)iSK+i�M�&:�ʣ�Ģ�"���{�Q�u��J�@J��P���-���;�������

q���t--�;�[�E������x/y��E�nVÿ���������Z�|P/�WTME����l���QP�mf��^V��0� ���u���z�.���o  �@�  ���'L�r��Y׀�����{�\!Ȉ��"��"d�4t�����'3yz(,>8D�-�.B���P���q��q�F�=�!0"�bD ;�!�`t������{��=��o�*52&����=�k�:��"��k��]��(��\Γ�qP'�f�T��Hآ�r�(lT}"wB-�*�����Jys�T	HhVשD�v�G��T0ۥ�fUæ(�4��]׎C{b�sƎ���H��N�ě ,�n����Y�!�C�1N3ұ��Q�R03�ó��#��N��KM�Z�h��c�Ϛ��cla2r����$g�N1�'(��&d���X�娺�Jx[N�Z��}��������0|L(�3"g��G�������di<46<496��kΜF8;y��!���<܂�>X�_|؃"1�hOg?W[G�!�Cl,�X/??'7��0k�!^^�h,������io�logkkoli$ r���%��ۺ��6�����y:j��m��V0r�bn��3�ꅖ������&|I�t|��+�\��[��߻+!'r��)v�X�w��G+����˼�q�asg�X+�i���'m�Pt�:�?奯�F�R����; AGn��=v���=f��'��&��_�U������6{ݩ��6�=�w�̽�S���6�n�VfƖ��,�
,8������tذaffN.�@� �E�O��DH$~!���b�eh�����Ű�<��he:�  �:\W�����dmf`i?n<��h<4�����xp�=V��f.�N&~��	#Gdά����D&��#��O�O�-�餼��Eq)[(�q���ɓ��U�m�e���3f������e���XY[�}h�a��l�;�Y�XZ����9���`�Lv�6fFvf�̆��������;�/bĳa^%���*�ɪ�Z����hd+	<5�<�yZ\����4�r�up"� q�����������=SLH(�u.\�=s�|aiiyMM΂L�=�82,0P��/!�}˅�4��T{��l�L���"�H�W(��|� �J�jUo?@��,S�%
[�Z�}��d��Uiumdrz��	֎.X,V/P$��qX0��a�H��;��#5=�@&�����΢�<}|�;vo��� ��Xy������H�L��ǗJ�R%[�f˴|���|��#nfH{K��j�{�o�D��X��-k�x�r���YI�n�锼�dw+��F)�����7-�6�����FN_0?9#-9%`cd�z��ϭl�2-�.#�yD�����;�.f��`e6t���o��)�R7oWG�K΄	i٣���C�2�Ϭ�
��v�X����]M�6�����+��=x����/$5jd���+�UB�2kbzx�{��]Bx �s���sg��,�x9Z�"���P�6+g��|z��֕ា��j``��3p��hghi9��������i��P��K�_ݻb�3��x��<���-��n<~*j�`57s�;���bs�̭�����˯&�?���u���[/�ue4N��k��n(*kqҸe\U��]�|C���۴|��%���e��u���Y��Q������N��`���C���������A�wЅ�UиmWfￗ������#Қ���I���w2{ v�h�cֺS7�������s&.��E����8��������j�`o��l�pC��"��A�����.��ʚ?/�¡��H�&S�"�\{0n�Z�`���P'[��|�\�-\��@RD�����`?<�WOX�O8�|4�Ã"����\�^��5:� �Wb"�3�&�N�s����"�p������>������j���R�oh�o+�LA�����e�֞<�KDl\D����������������������	l=l���q� �ln�nv;3��)\�	t����q�#B�>�`=��Rŕ��w#�G`�L��I ,��EQ��_�+�w��������;p!8�WW�-�P88�Bc@,\�r�/g�;q��������D��*e�Y�Ň����.�"d���(��� ��cӭD��'*IT �DD�R�D.Ӷ�������oo޽�j��T��5�u��<��I٣�DGG���#CP��H �_�������  � :��?���bjn1�����X��y��Nٵw׫�5U�K^=}���W,(x���C��q��%�S��g!V�E(��1�=u��RA��}��mS�[Z�֛ߘ�)�Zm�ZY���HEd�Z�_��|�O���n�05��[֡���sFE��'�&��C\mͷ��# ���볣���.{W��}�=���е�2R�'M���;����u���?>yD6&��"l`ȁI�V~K���W���o�d�ڵo�.ۼ�Щ�N��>>>XlH|lxdX����_߶�D��"1���_�a��H���u��K��[T�WR��+p���^y@LJ�M�ǹ:70300b0|(�{@�3}���K�;���%�����J����Kd8>26�?��q��#y_���S�����u��Z[�:��L�~$��.8xjS�}��q�s�#'n��\ؾp��i�w��>~�
�Lu��������p���+��;�^�3b�Q��E�Rm7S܋_,l�8=��+U���fn,��Fl�t�D��L�ƫUs<\z�Y��3v�Z${i>A���_Ο���ą{�~�q癬	�B��p�Ht`0���	������N��INLHNN�����%˖W�4�U��9X�kH�
,kf�ܝ��酰��4�p�A�����u}.x�[��t��r�B"�Q^��.6��������ne�h���0����"�������޾_��ؠ���X-�߉p��ž�^��9�\"݉n��Ӈ�!`��v��C�YF�G��{�&60p��ƇFL��<"u��bRIZI֐�2�La����1� �@�����7��_C��[����[�؛YٚYY@�����篿i���CG��**.���'��t��!�w4�$B=�K�z����9������?��+U�J�H
�H"�R�X�U���3���[$��Ě���O��ڦ��а��Sm]|}}Â����1~`',��� \�M_��]� ::��[���N�6sρ���.�,m�n/�D.!�*�I�H�5e:�_�P���5\E���B�.���׺����RI[��������Y��ͯP1S�� ���&�4��ϐ��͒��|�a�	I!ظ�D`t/�%fܷ���C�8$��|ɂ)�7	x|���l\mog����y�/gILK
�Ӌ����7�����:	�Va����O��/j�fi�Uo?.ݴ��� ����_����zϚ2�O+'�>�=1.c��5K��v�3Ee�'�NO�N�ψ�%bb==��#P��/rJ��!V������5p�4p�6��6��1��5پiY�h�s�G���u���AD�{ZJR����Y�GN�~��mag�k������g���$����$�����UJ5����W-ɾBܷ��� ���Q��țGL����?y5�Q��+wso?�w��qW1�ߌ^�I��<��Y�o$�>i3�5��˪���Z]����ܯl��V�r�JU�%�?��������_G.;"�ύ�����n{�(_��B�̍N�۰�T��9�����8����c|Ѩ ��Ć`�qذ�0,�aU]#\��o���B-�q�����ܜ��C�%c����C�kML����
�wM�M�$ņ$E�'ಒ"R�C�Q�v��>u��Y��� 46,"����"d
p�q!\} �퀷��~����"������-`�e����g��wLtxZRl|t&���u��p�� /�C�m(������x��#]�~�>�fks| z��I�7�1��ˆj���ī!��H`-
�I��i $�WE�^~z�72�nb>��l��1`��1x�����@.[�
����/_�TT�5��t&� �Ά�L�-$qa,��'���٢o"���� Bp$Y|`C!�E���ΣөB!����ɤ?����ݿq���n$�?	:����$�������s�������t"D��QO//o������;C��=|������5����t��f�l�FƠ�
1_��.B��!BE�GV��/�c6���$�s�dܦø	�q�NXh��������[·�\�3_�m�\=������~��y�c@�k �����g�dG�Eed�ۻ�������5402:t<��q`߮�3&'%�E�E�"��RR��2G�KH��IF�'�N�[����i�N�=��>as;��C��ӼM�����BzFD$%��H�]:���ޕw�Љ���N���;8�N�0&5>v���F��D�D�<�.V �eb��QN�0G��ڶ`\(�<������,Z4s��uO�]�6"�����X��mA9vl��qi�^�����>��̧�uqz۸�-�}����7�-��yR[����o��=]Ԡj���3�۫��)K��M�u��F��D�I�W�����ĝo�O"������{�|���˕j�N>i���W,�"�m�^!�N<!'�ڹ`ߍVz�G��_To�%/}�*V��]�FN]����u�N��8�/0,4,��b1�!a�!� ��:���� "�]�oD8j��էnoܱ-)�z$�r�5������6��{�'�MF�G�!ctD�����������X�9">����o��}���'�����/�#p�t:[$�)���־O��3���œ��*[\��������1����p�p�����V�u˽�콜mP^���6�v6��v~NHgG��C �	$>���ϝ>�Gń���P���]����;���wՆ}q�3�jj�6�E�H�H42�\Hc� \��Ua0����A�!p:lȰ�� n]4�@�C�����X�r��S��<����������H�&B� ��0\IKXO����&������7���3�-����h`�*pX���
,	��ɀ�\�X&~��iUuŮ�;Μ>���uG�v�q����攕��Aw�%!�pp`�(X{�A��`���������� �ǀ t 2���Ĺ{�Y8?zR�[O���p�b�X)<�QvuH�|�ؚ-�`mK��l%�o��7����[��-8z;lʊK%�S���<g��;��(}�޹;��ש�36����!��'�u����A��	3â��㳓���S333�G�猀ӟ!<����p���0c#��&�C��f�$$'���&���$''���IM�LL���Nw��x�W5igm����ԋ���)�u¦�;.�tE��Vd�_rJ����P����yX�c���F���DY��E�1(dX(fƔ��G�����p��?1����O�eP-��uB_�����i��m���������nM���*��TD`���Mb"p�Qa��Q������gn��^y.(~��:E������7����N�����J��0��]= VW�����-��%�e�S�+��xJE��Fޭ'��~����D�vʪM��A BEG����G�=��t �"l���1 1E�go��]�+v��kO�+�RU��_~.� D���;%�FI��g�,��j b���o92~��#���zT2y�2�@."��c#"q@��H�BC�q��Ņy�,\����>nU��� j���ɔ*g���SW���H�M���"�¡�Q� ��-�;[�ReBNBZ|H|D@B8����9.36+9,>�?'5����-j��mE��аpgD��y��D��+j�
T\��+�~�opm��_��"��ڏ"����"����(�H��������G��r��7{�8O'k�����=��"��E���� �R�y;����5/���x�D����ˢR'�S��
����#0IT�\B!�����������#C�s�@._��pρ�O^�VU4��l����< �%4q� 
A@l�2�V�Н���D�E�����+�3�, B���J�M��~ݪ�����K�V9}�����䤸�7��vw���ob�4,,���6$DR`xP ��-�B�� lA4
��QAa�Af������Y'B)@���B�H�"���P�@"��<U7�{5�qkjZ�%'$�����$�B/�=+���M�Z�~3~���'�6(��5�=jT.<pm�/w�o�9[��b�'̎K��0&-qtjJvrzV�Ȭ��� x�#�����X����lm��I�E��DB� G�`���b2Q�Y��ˮP8�sW�N����k@�m�ur�����K�n���hߔ4Lr|������m��b�i���C[���
�E�ÅbA�����d�����4".jtF���Y3'��;sڼ93�̝6k��)SǍ;rdfZZJ����}(��������sDb�#N]�>�K?���ZY��������E,H�h�.BV��XP�٭|'j��{U(lnm��t�([[%�f�Z�|����*�@���ヶ�KK�oTi���zn+M���	Rv~aJ:������ ��!n�{ ��j ��o��=S�>�{���Kס�#0�H<��Ƈ�B�P��AAAh�=� ���/^��!L�7��ۄ@�S���J^�؈��(�ޅ8� ��p�$:�����1#c����YPO*=.ddtnbq~	��'eܾ~�éo �G�D�Ǧ̚���ID���._�݅?E����&��0u"|Y�Wr���&rYM������j����H�q�1�x�#l-�� ��6~N��vH� a��n'�5*����c"��C}A�n�d B��S�;��5",a��rf9QVAV� ֓� ��,�	�Q�C~h�,�a��ή.@�+W�"ܵ��aShd�@(d�t����Y<W���^� ��v%_����"��xt]*"||��9��E�f���x�ߥV��͞:*+mܨ�wo��6����\��N� ���h���΂�� �с��:�.ԉ��EE�{�X�?xR����Y8����	|��E(�F(��w���P�6T��Xq��uǫT��U��ڠ���q3v��M�pqۥbn/$~qz�-��g.����z��:qv\Ҹ�q�	�ӓ�S�2A"��"�%B#x��KskwWG/Gogo�!fz���D��a�^��q#�}��8]Cy�T�������7wj���f����9�nϭFx�#�痞���t4q43�q4w���`��E�X�"D�@��q�F"|�}�\\�����0ph�_9��[�[76�� _z�]�066������/HX�X{��"�����/��CF��7��*�@�]���vvO+���������� �������u�B�(��D-�|�V�nѭ������nYπ����*Bu�uϧ��P�GH��E��������-�&j�x������������M��o��_�=��=_?����g/��V�ݎ�H��D::� n>^�~^��W/w�������]=��,XW�m �\�-6���",�p�W@Č�����}[2M��@_�Hl���mR,�lb"�Ã="���P	�I�	8��P�8�or�L�' ���k?qt���	�����"f�]]S�o"+��^O��)9|9�)�O(�!��~�)�/�߉������*�����mm�fg͘8�����lg6<��be�eg�!��������5 ���p(?O��x���������o�@7��"g�Ш ��zaY���UM`�dx��� �ӥ�om�p#cS3�0Cc�u��Í���Q�֬"ܶk�㗯_�T�ՑjIL`�F
���i��L�4���[�N��Pח�E�*�B@ �g�ﷁ.�>2�"\�b	���$BvW�Z.�.�7c��1��"5�vwvhT
��	4j���!@o� $�#@��.Bw$
��jj�y?��#R�C�t"�He\,B�u��%R��[�:�d�`�]�\Y]�vo^]���*h����;s��*�~�Q)Gg�x�蝺%w��ZJ���]z�V��m�7ЌmG]��ͼ���i�G���::=cT��l �L}">���+$���
70750�������>�����4""!��0&`�ܓ��RE_���%4>!8��Z~w��S��+;��xy�A�KHHJ	B:9Y�O̰12 ]4��S�7���� B,�����F�`�1�8 x���y�[jdan�`����`iihmc	�`��Ņ��1#3�Q�1�1Q�\�g�-�6hʊ��EU'�������ngu ���z�
�-��#�����ۻ%m�m[s����_{�}i끧�eJ"O���}��O��y{��,��"|�w��u�������������onhi#Sv�T�u���_��V��U	�v��"���uqq�]�����fV�v�Ύ�nN� wW h�@��l�y�̜�����(��PDX�ɼ����&M����
�^Sl}=�������.�Lm�bѮQ8��p��0��7��6�-<�2�p�Y8Z =������ꍜ6{ye-�� �g���Ͽ~���O�li�4
D��J�,�ɇu��WT��9�X[ۺ:9�99�{[{sck��N�FΖ�v������h	�p�pw0u�7qw0w�1v��`=���k>^w[��~�����������Z�^�UM�j]/B}"�aaQ18!����� �L�L�� f`���H|&��V�]w���-;v�����A"�"[J��I<)!�D{ыP�u�UTl��'T�EB�^�:��5B�N�|�X �A��,�w����O]�=�w��C{wo�r���i�Ə�����\n<t�^��Nus�1H$|��+����_���#��]}P�t��k�ӗu���>���8����*�2��Rɓ�y2-<�C��`_,���!�0��~��>�L����O�ל�k��D����q�2sٱ쁉�/|� �
� Bۗ��{&l;.�M�r�#*mծ�iY�S�'�%�NI�IH�:2<%�����CE�E�b�q#s�ҳ���C�	�����������Rs�2 ��g�]�m��#�g8U��ӷ)cy�6is������:��.�b�8�LN��������0���;-����������',<4,��OJI���V�I��M����:��(V�.^@���@�� �Ň��b�q1����~>��I1�k�P��,�~�%�ۤ�0���ݰ���;z�,�+n풶t�Z�����Rm�7Z;ĭ��N�^�ʶ.�����^����� *[ߨ�ނ-ȅ ���R��N���F=���y��%�vO������*!.<����������������������������������E�E�1g������Fx�L=XP�D�#Rj��r*?}�>��I�����,4���q��f'[cݬ���fh?{<�=���y�"D9G�] X�������!��,
��E`���� T(n�̥���F	G���i�����\�ǯ��,�����D!K�b�KJ��ݬ,�\�\]�]lm��-ᥴm�� z;� z:X �ٙ\�u4�Eh9^$b�������7�!a0>���& znY=�߉�����񽸝�|z���YX[Y�X[Xـ$蹯Y����s���w"lb�areD�N�����y�J��k��U��E"��Ҩ�B�?,��YP'BxP
�^b1��6a޽[۶n����~~[WU�{��֍�6�_�a͊YS'�GG��x{#��ľ� ���������;���������D���_���s���v�v���F栱u\��]7�U����"�+�!�r�"0D*f���zԂݥ�/��N\s�	��S
 t̪�	�h��SS�\�^)8�����%���79m4nݮБ��m؟�5>����%����H&�9 ��7��7�+4,8>����u�	����â1��ؘ�Ȥ���1I#'��L�fLLə�5w�cҘӕ��TŴ�G+� B�Z����ww46�f��D��>:)�`t����������sC�P lAo�����c ���	S��s22b�#c�"bG "�2âS��pkOC3{+{� >*�
F�E��&�������qq>AAH\hL�TL�ғ�Lnt�um�@DԪA��w:�m}�����M���^�@ p!��f��"��:at��?����p��/��� E�{e�;����؂G� ���T]���_���	,B���@���W�T�V����qt���K.7>�Xw���4t(�:X�آ��K��`����
"���\/��Dԋ��¨��R�F�O�G����E�C}@tw�p�6�63 ���"��zbC=cB�A� ��P?;��V�lM|f�D�"�4mQi��^���M���ӯ|�������EX^]�����18��<�w����D;O+K��ݜm���ṁZ8Xy8Xy9�x9[�Y��������t���%m6���.Ät�����S��7�|K��4J�E��^{�D�[T����1�������3����R�����n���"l�puT�z����m�?�(P�^� x��@؂�uHX������R�^�Z��J#vt�|�����A���Y��'�+�=�;z����k�� Y������������#���`#qQ�Ȩ�(@D "":",:
������?f�����B���+9O��}?�s���т,(�5���"k?�*v��j���G�<b&�Y~(${q��UK���AM��s��I��56z�EG.�-j,W���Cӷ^}���5�b�&� B�� �.�V����~F�^6.Cm\�]}�!�9S&�¥�qGG���G\���ў���8@h\��oX@�����LX�[�忇hmj�
 B�F��.\�&-,����urs1wq4G �}���|\=}\G��غk�֝��sr�M�:r�ؤ����԰،����a1����h|�oP��?�����!5e$>*	��<"'s􄴜�I#G�d�~��2q�Iɣ��Z�+1sﮣ��W������[5��^a�Q`@�=Qk�w�
�Y!�z�(BYK�N��Vy{@����Dا�z "Tw�Sv���m_�m�U�UͰ%mD��V��Q��Y��E��U���7�`����p�Uy/��jh�����c�ܼ�,����/F�cӋ���Z8�e8aK�`��0�z��Dm�2+�┅{�`�2��G$� F��q��|(H�N���R�D���t5��g0l�ԅ����:����Q�L����~&���iaaI��e�xT�N�._SQN���prvv�D�8;Y:ٛZ���>�����!��N��?n�_G���
<�j��4jdg6��X����r�������5
D�������e���_�Į!�~!��������Dz�y�b�PAhOo/ p��(!H�GN��b����_����IL`A�BA(.�!��i�::���kb��.�q������fA�%z�"�v[N*$SI\W۪%�*����PQ]J�4�(ĺ�����^%���������GgF��O5c��E�.�4mɄ�`f,�0k��Y���^2z沬�˒�.��d��ݗFO_���Ŕw�����WJ� BI�7`�8����U,�k-���{u��[NT/��>�	�
(�F�;��3��RNG��t~5��S���R�Y��"���v�������Sl��9�30t20q10s20��n�������n?yu˱�������C��������P37sd̨��sV�>[�T��66�u�_�;;��}D��1k.]}%޵�\JR*6"4%3���B����Q�}=�o�I3f��v��՛f̋I��Ǐ@��!	��ظ1ظQ!1�A�阨��쐘���t|bfJH��S���d��>fڼ�ɳ3&L��5.v����l>pqњۻ���s�y�=t����䧳�Q뀨��/l��S�0���E��o[e-oA���\�{i��㣸�)l�Op�]]�yY�I����ߥ��I;�J�?K�>��?	�?�;ୠ��W�{z���C�^H�#�[=8͞i�7罨)���ڲ����mbieljdh8d�0xe(�C����M�A(444tpp�N�3�QqiA#�5�\�DѰ�B�� �z��4I��'��^|x���䑩q�	 �㠥����������%����������-!����eo��l��d�t���y��z�D����2JU=�Ɩ��^�T��џ�_4��3 ��,��)���r8L����R�\x��P 騪a���Z[��[Z���`B�����8X�;�x8; �����.ξ�.�ps�us@�����31p4��B!nn.6vNlR@pʭ��/K�Q5�WKb����a�h K(|^T���qA��y�{!��A�!h�@@@`���(����z��Z��БK���Z𲰬����@m á<)*[D`a2��\�C�J��b5]���2��,�
���/Ȓ*`d����	�[ :��gp�DE����t��q�RG§�biC#:&	�9�:(� >�i�i�;7	7�7f�O�ϘɈ�	�c�"F��e!�2�#2bG�F�XyEF��˞SMW0d�,Y�~�>�-�W�w�%Zj B�L*�)
�Le/]�,`�?2��,�;��=[�l��w4� ]���y�Ծc��㴾g���v�|��&NKv��mt��p�@\�Oh�Wh��˰	H0�b��p�/W�6�r����;O�u�O�	�w�wH����y�$e�\y���E���KX�zqk�P�V5�-��:v��4i��:��W�$��n
��:q���	���:�bC�b����LƎϽ��Z��k�^\�W�<3�'d����g��g��g��;��#�+8)*}J֔%筛�p��E�'/����#$etpr�7�r�����^������E�N>���,�w��4���VQs���_g�qK��w�-=��Z�D'��CݥQ�Na�@� T��@lD����R���_�� \@���T	�@�6��8�O��O�g��O��?m���C������N����Z�(�7������]�� $}Ջ�%�d��H���s���+.\�iXl�������������İ��bR��C-M��X���Թ��4�-�}TEx�D���5$
�uDZ�YB'.�k�Ju��	?*�03%61�Ur�qs0F�՚�Ezك|�	pá=#�}�q�	�h@> �����n��d�����&=}�PTN�ij"�:~�T��Ҹ?�����~��g�K�.B�^V[SZ]Ma3YB�N�l������=q�"c3G��2�������t�##KCG[sWG;�OGWW� wD��'��+����kc8��hp���A\4��E��z��F�&�ͯ-����5$~=�:��R�N������gQ����`t0�� ��!����U��8�`ъ�_>{UVZ�P�@�m��\H��)l	�%�O% �Q�@lZ���-o�
�MliGL������B�"�R��HU
eksϻ����:r=[̑�(�J�RD����yy�wH��|�]�\��ZΑ��/�m�ݴ�fݞ;5��~Ps�Q��'�'�k�<*����ڋ�+O*��-|ZI���V�<Ȓ�)Bi�?D_�����/���U ���V���#����rd￡x�U����-G9�T��T}lu?G3�׾4�巼U��j���%��N\z�6fn`xf�����LX�0qy�ĕ������Z�b������7ˏ]/�z"�'|�_�8��1 d�Xd�h��[�(7t���[�6�_���"!�;���&���l�i�$�����)g�[����K�^�8���w�ν8o���.-���7f��_��w<�������=�0�p��#Icv�dm��*.gi\����q9�&�7��{l:�d۱��\�w�ҭcl9w �2��c�L��y��>*��fgދ
���ʅ/5��u�H�'��E�0z������:�o�X�v=���ꘅ��������[s���_pz��G�������-��
=��r�(վm���9}�e]���i+g�[}�V�����
U��F-�!{�4�n��F�ޖ:m�/w�����W���ľ3y'rM_��78��ibmida8��`����.���p+3#`D#;+s/��[��m:u�I�IImI� �VMb�W3i�>�`���(��Ĩ�<��x��.D���D����������9�������A�c|�(/�����������]`�kXdHdL
?����eM5������P�h�P�>�����+��lmay]��d�4���&�&���(ڳ_HDT���������������������������������������v�v�^NN��.H� w7{CC{�mLBC���N���N.�n�����I�dH�@��=<*[/�F:�	��C�Ow��@�_D��A����LV�X�gߡ������eyQycY	P�@��?Sl�Ȓ �I�b�[9����"�6r��A2_���<F͖)�[��ɿ����K��R��\�pX�PΗi��6��U,Uq9|�^�P����çΜ8�ڳZ�"�V�dAÍ:֍:��Z^�����~Ae� �
H�R2���+�#��l ��*�r%�߁/����/��y
)O![�B�V*�J5S�FO��l�)Z��f B���/��Iu"�~d�>r䟸ʏ<� B�j�����{y�>��O�p� �.�| e���h{o��+��;dA��6�7�?�1t�j�C�(d�,�q��r3��b����������q0^1^QA��A�uB�%��7z��G��4A��H���Ƈ��V�	�E�Wo��8ru�ȵ~����L���0���/r��?�W�8*�I��%y�R\�2���G/r��4�?55% f2*��E�CF�J��M��2	�<�?~2n�oL�_�(���Ȅ1 �ı)S���MĦ�Ϙ�0!gک+��b-K��*ڥ�N��K��i�E�NIs7@�@Y3��$.qk������f�ң��,Qo>[1qg�:�����ȍ"����M�������C��rt���s��KMB%ݥ˦8w�5a��/��yDi��}����A�<�L��6(c����4zɾ�/iW_2���, 7��|1i⚭�n<{g��!.>��N��f��fC--���M�-��A(�21twuC�GgE�,s�MB&-��:7����YOd�]�]B��,>d�?������������`ieq�k8Z��q�5u�����|���p �f�Cum�P�NVT\�ȑ�#�r��K�j��H�&&��� @�l!SX@���[���-B	O'B&
Y|
S�D���u*{��#�.@����,��l�l��l�M�l,`�,m--l,̭ML,��,����2��`������ ژ��nl���b``f����������7�*	\��"��0�)4 ��{���������������A��7��>�~�'� :�^�~��c��|���IaeQeSi-���PRG�hb���e��i����+'�$����6�l��dH� ���E�2�������#4vce�˼��.\>p��gv?���΅Jvic����3q�gN<q����'��|Q�@T��r�,f�QH�R�Edr98 ,f�Mf�i,�N{ߖ������B G-a��dMQ�A��4j�����}�Q��"���e�l�;��]���������������}�U�@���Q����,|^A����b^�ż��+��U��Ws�~�ɼ�S�	g�i�� W_p�ϙ��.�3n��,� nro��2�JX�h��=,e�~�T�T�pT��,u�^�\u�����-�Q��>Q�,���
iQ���Z����%'���������_��Y�p���a%�A���+ٹ�|���2Ńr��*9�^	��c�鼪��5W^4 r��^~�뮾��VH�^B�YF�UN�WIZϻ��������%�8�V��],m��:�
؅p4�t����P���m7eӂ�O����Zߪ����/0�}��vA'P�����'*�zM<r��U���C�K���TzR9}�y-�CP��v�
�o��$�$��D(y=#���Щ����63;�Y�/��/��1�Ĺ+Q�X��tD�ٻ�Xۛ�;�;:X9�۸9�{�::��z!����0i����5��[gl�4r�ڊF~=�\XC�P�ן���/0��h������P���О���������n���B�`J����;�XU�n�� ?w7;GG3{p�K��8q~tԸ?E�@b��O�l��}/�D�S�6�-0���!���p��3��lٽoopH x�
W���B!\������������ft��`iigjfn0�v�!��������h�����&v��NF���y���.�b��#�بl`�Z2��Dи�'.��nΖvV֎�����^^� 7����������N��E����yQuA%�UE�����jRy��Q ���:���)�f�Բ�ulE[U�R6�� �e�Li����^�\9�*�")]$f˿����D��������W.mlxA��̻ux�ډ;6N۽~ھu���@-��%=f��\0>n���EgW�זR������O!���+�{����5/��8<�FD,H�
����'<T?4F/B���\.��"�*�L����U��*R���.5(ϔ
ξ��۾2=ly\�^��V�QA�P#�C<��t��g_��jl��jzٚn������0%�q�'���0V���������J���녜�Oh ��>p���/+|Ԇ��e��9a9k��zu�.y��1����\���R>����GM�gO�.�WL�����$�d����Tv�/H��6����ts}QGK[�$.��<-c�yR��0�Ki���U�g���pپ\��	�+[#G�LZ��_怞��l�+/�Z˘�w��r�:u����W{.?�}^�x�e�Ղ��Bbn�J	!�h��v!�i���)'�U4�|X�"�P�"�����U�L�)� �}S����Ϛ�u�}�h�|$�g�V�;6?�4|��36���[!w��� �*Un�i�	'}����@����-��n��|ޡK��ߤt�2�\���.?�3�P����.>��]vd���h���ر�_~��𕜩�	��� �/������C��"�}<|�P~�`'��'�?0($�;8=s����7W��g��G/�l6�x$N=�WNUL�y3{ű����f6fF��02�G1 1D@��+ �� ��̽�l����C팽���L�����=663*b싗��rbuC�\�`�D?E������K����,K����\*[B��O���q���;w����yLM�]��1ֻ(��
DC+{[kg{;W;;���ǄtvF�30̝̆Y����;Z�{za��qɓ_�q@(,�d��2j�������<~���a��dhfddnllabO�����Ő!�LM�=<�<>˗�޵����K�_��T=)�^N(��֒�,��&��������(��@� �s�zyZ���.mՋ�ϫ��D�/���r�^�kV,&��sɏ��ܽc��}�'X7���1G׌a�:�]�w�>z䀶���DM��0x���f�=R�n͕����������uS�j`	�[�R��v�?,�!|P)RʹJ)S�&���y�@���;MNw�N��8z�]��r�;������ͰZ R3t��9{���Q�lB�b�wm?[��~`7��E�Q��#�i�f�@C�*u4�N�L B��n�f_+�}�@&-�����m�]�Y�oL\}q��s�c7��Xu�X�2eW�u�ל����\y�!�a�����a	Y��ARL�V2�SB��1��hc+[9��
��n��-��Dna5�i������������x���a�I�%Y�t_�S�"L\;n��E��Y�l"w_���)�3z��ECG.B�;VH}IR\}I ������_E��*Zi��D��q�@�\�B����ޅR�?t�7��;�ᵿ��(/�^B�i�.S6��Gn:u��+���@d�oG�4�`~��q�&�㲋5�]+־a��Җn��w�h���~��j�"gn�KT��B�A�[�2Z˯�}� z�:g�s�v���+O��l��K�S��R���~A�~h�`,*���B1�pl0 
���#�#3}S�\,�l�R�6o���������E8f�E�Z�3,��F�|��$F��CQ@{�F$!=�>�}I1�Hl���|�otX`bt( ����IJ���{{���F�|�XS�(���'�O�l�����huuy�?DH岀~��&���GOܚ>sYtt������������������5����������Y�d��_0�tq�p�	��tw�40p37��1�u2s�fk;�������= 5f���3�0�ʹz�a�	D�@��"tՉP_yb�p���C�l�y�p�cC#w����%+v��?m���K�,���y���]M5��D~� ��֦?!�: $q����.m�_8��~L�\��yY �/]�����ы����kV.d�>��^]ߺoe��u���ul`���X�h�đ�׭Z�z]O1ǉ{��R[�go-�7���������RVsƜ�A)��*���*k���� ��3(dz�'��-��e_��K�J��� z����c�9L9n������� �X����B�����{�F�=�������033O������9q���l13�dYf;'3�?�v<Nf�y添�~x7u�W�-�R[���S]u΄#���$N9�?`[�ÿm��R�jP��  ����f��_������0�ߒIk��~�u���d��ה�g�����_|�>�=n경�SHuk>_����Lѭ7�繒�Oq�
�O�mE�����@R�C��L~��ZT��[b��EN���g٥OrJ[DX�N&���7�a���蝡�֝}�Z\�����ރ�l��L��v�$����eҩ����e�|����x7�p;� A��4������Ʌ-"ıۈP����<D"-��6A!��Յ+<���c�Y���n:�%�wG��%�ۮ;.��5�yP<�Ѓ�*$��a����/5HȀ�4=¬E���V��\²cWH���}=w��be�VŲ�&o:�iF�Af=7r6��s1����%�����/���-���u-w䢣�N>�}���9��;w�O������h+BP`����	�=�vNp����0a��of���g�㬲b
�bAb�sI�Q��.?�x��c���鞀� � �E����s��iBIn��;�tI�
Ɗ4pW�.��{��H���'a��9\^yZ��;w�%����w����\BAQYN^>D��C"���w���,���ڊ0+/\H�S�<�O",#rWo���y��+�m\���ξ^N�C?ogwWP�l==��\��@�� ����R�3��6aP׮����|�;y�Xy8x���FFN��<����7ҟ$��Ů��� ��]�\�A��]���vPzx�W,_�{�A���G�󞤕@|𦀖Y��'��o-�J ��
�ĀW$� YZK2n�b��MD��Dht�R��Z�%�K�y-"L�~����O�eS�o?�|�����GV�ٷ|.����U��j���n��aω��5O���O�����g�;i�>swSH��V6���YT%Nd�#�J4�[Jhta��"�n�ɾ(�nn�L<�9�T��;���P?� Ug��d��Q�DI��\��v^p�S�R��[��zq:E�%��X���l�)k�VBD`",cH��Bxc_�3��00^K�I���^0|ə��v1�gn���l�½O�9��8mә4�Ą�k#-���R����/(�2�<���O%�s�R�c�hhN�hhR5M�dr9K���@�cr����"\r^�|�t�"�\�4��Q�q!�y9�%Q�p����wt��7Xs�����̭����S:m�U������w����՗���8wS(�R������R�o��n���J-����AJIR1��YD�ӄ$��2�-"D](׷�P�2���3ơ���E=7u��$t��2ʾ!��Ȣ+)�����ĵ�2�Eܪ	�Hkv��R�a��U�6�yTL�@�N.a�����l�5{�����FF�Wn=®��8b&�⣬9�8g�m�V�]��B���o[.��{�'�>��hM`L|xB��ب�bBdB|$fAL���.����1�n	�|��˒�9�����e�����p��{S6\�=o���z$��H��/��-<���z��A.x9��0zt����A}� q1���3f������7�OBC�#B�Ϟ�*-��DfR��V����Z�z"�"T2����G���]܃���\ݜϞ=¢���ϙ9����κ#��@Ԃnv>�����>v��6�>6]c�D�"	����-]��;������ڀ�<\��ѹ��W���B^n13��E�e$:�Q�4;�M
�;3�v��[��"S=�w����r��=��6wQRFѳ̲�bƫ����"V]�A��x�DQ9_��6�����2�����+��.`A�B("-�����k�bC��ĸ����$Җk?X]V/��=y|��ɹ3&��������,����E'��ڽt҆�cS�\��<~pm����gN;s�<_��>|�闔\BnB��>�I��M�p&�>l�"q��!�m�>~I:Y�j["D�V,.a���#�Jt��4U�Y|��.n��=��&���	�/d���Y�"�b��2uQP�5h�ۈ#6��^.ґ�u-�������|eOa��+&�!B5��$r����!*����"�����>�\Me����[�8i��'L��	C�8%L7������k�m��ab�{��}�����v7��T }��z��z]�O/e�ɒb��אj_A��)E$�O 
Oa��SNJ+ơ�^�^�_���OK��C2U;g�-��1�����ך�����b���:rB�����,?k4���Q���{:r=�I�~
�Q�Q�Qf���2�A&�^z��Ԓ������RZ.�]L���!�إ@�=��|��/CWS�Κ����C�kKˊ{aE=��Y�J�����w��/4�7f�����t��
4�_?��0��,���w}��/ � G��W�7V����"�y{���kǙ�w����`a�oH��_t*�x��E&�D ���!�q὇���o����&~����/��
˨�e�<;�(����]���9�Oׄ>��0�|\��	!��'�|��K�<nHd�WbLP��`�k\h������];�v�6�o|�Đ	���~uG&����yy;yzz�=%'O��K,���\�#������� ���<<�D�~aN��#�������ܩ�rK������ֲ���9*B7[o[?���
���6g�3��xq9&�2&�<2�4�������������ۻ�9y%��rt�5&B�d�qa����:tlשhKu��,�V��^>�-ں}'��qJ��7�7�_�R���z@��(�Uf���\��y�M��"�#K�[E�
M�FCC�
:_��"4.��A�T=/?�¹S�&�|~�]���zo��Q���ع����7���k�^�;�蘱�֭[u�����|��mW��%��2m�ٻF�95f��~�����������x�=�/H'
�8�XP���Z/J�5dY�*�g�+�1��O{��	U��'���y��t�����(�_I��tz�9j�)��A�{W*�5R�R'T� B��A�$�DX��B��2d��b��\��[9���w�%ѣ�v����c�]���sF�y5��#��r��#�-���|R��T�d�M3����X�S�O�I9��A6A����N�DH()BE(��� ��`�%$���.d���98z��^΁����z�ē�W�w�c��/�H��ݻ�����.f�Wv�H}�P�0u����3v�#f�>�,[�8��8�8��IV	���s����HSK��e�<�����C-g0�$7�� �¿a��I�F�g���z��E��[��-�OT�>@�������r���p��J���o�+��4��w<]3_�n�U�X5*B��Y����W���q�Jҋl��u[#��DG�{{yx{�FGF�GF�������aq�=cz��y�ˬm=��t;oӁR����QR�*�qA��w�u�ݭwb|�.�'ƈ���e�g��/�I�p�p�����"��V�=�Et���#b��{��<aw��QnvcFO*.�P��_"��K�����a"�P�"�p�6��FK���}\]݃}7�_����;WN���؛:ۚ��trv�B8�F�FzY��4yD׸�@W ���׽������������/�0��han���[}�q��т,���y��������L�aE�P�u4�o��۵�vq	���2i���+g-X��Mγ\���gg�;t�a��2޾KO����$9QޔT�[}��2��B��IpW&Y.��j�:_�P�*B�@�.+l#Bԅ� B�SX��s��ef�?����Cw�X2}��)#M�l��g޻�̱�G�^0o<���{b��Mv��%��-�7xɁqk��?�bqc���ٕ_q��l�t�oK3�l���gU�a[�6"T˫�Mȝ���M�v4EM�63Tj��
��W�bM���HY��X�s���c�. �z�@��� \�Iu�@���*Bx~�i���a9S^�T�寋��C�9|��zȀ�����w��9a2��~��V&�N��i����R��av^~�Ý��|D�ߞ��f3�e�^�2˅�4 � jA�5B��p�z�����
�2�#�3��4!D�E4YU�G���T��3uM2Y�Nذ�/�U}g��1}�R%(�A��n|R��9i㰹N�'>ɔ�O[��nR�I	�(0�x�]nx�MLΣ�ӳ���zK��+����aǸ.E�*B�"B��Ho bU�`��]��p�Q~(�ϯD���Gj�M"}�P���;�;Q�*z�=�O�IK)��޶'�W��`;g'go?_7wOGOwg��������;�ǀ��-9��$pH��[�g%�$e�,g�sr�i[������vh���*>2�B/[�z���Ct�OBt�O"���b�����Cݺv	LH�=�{D���U��c&�S�Tai	�� "���@kz���_�e~�[[ff�82��f2���H�;�x89��y���Zo7kS4O���EGW'+WT��^�^v���^����i��u��@P�����������k;O3o[g?7'_?aL��/�@��8^]GXBb`!�tD��&��a�v&@Gt�EK���w��<���Ǝ�����f/��2{��c�qfo<:l����3�O]���S0_���̣��A�.�*��6���{쮳�H�I�J,�:�0�2��/Sh5��v�N�1�-C!���z��4uʄC�w.�=X�xΰ=G�?q܈y��-�?gѼYK�]�fզ��ΚM�ӹ�H�'��o�0rU�skf��%�$*ᨄU��}KZ�3�� �_EȖ�eU5d�ۣ�U�{�<s<MG���TkZDh�TW�ğ���{�+�#�F>�}�=ae@��,�g��=O^�V�XD"�7�{P���b����9�el�\"�n:����R����ξx��Q*�s_����6&��`��3�KyTū"FZ7�,3e�lt\�/'Ձ1�T�j G�/z0\��� ������)ekJغ�O��c���1���ɫ���*�M��s��e�d�*	'T(x�Wm:��>xH܀	t0?�H���&�%�/r_��I9�7���2f>�WB3f&��O�)���/� 0��D(���^��e+p�ΊZt(�Q�{���A�c6|���̃��r����������kncmne��lg�`mmcjkc`%�\���|�;�F���;+fʎ�e��p�t�� �+)㔕�`"��[T����㢺�G`@8����֝ ���%26�/>*����s|((D�����ũ]h�C��ݺFG{�����L��������b"$��L6���{P�hI���2'7;;;o/7gO4�y�N&6fhr�!�Bow4+��x8��8G��{:z�[8t4131�ig�be��d��e�����������7��k|^1Da����
��!���¬`i�	"B̂Mm-,�m��E�n��~��S'O�4e����o=M�t����YO����m<~?���7=',ͤkX��[{xӉ{iD���ɲ&�O�|���P%�x�D����Y�
*�4����U	%|caB:�Np�t:���[��A9r�>��.����a��KW� �v-'/����d�<)U�#�-H��C�����J��
A��@{�P�1��OFd�a�������)����#N�Ľ���!�o�j��ٿPH<���C���G��c�]��~ɯǆ�6瑴,i}[r�z̵�W
ы�l9�.+��J������:y��-'v���"����֋�Q	�}�C�r�/�w�.�u���7^�%3�����";���g�
Y�b���#���D��"V�i�Z��0ǃ	��ʃ�A�p5$���A��9x��VR����x�E�f��__}V�4��V.�H-��c����v����;�˒s�r���K_����I��I�+0�JEWh��K�D.��b,W;K ���D�&�-���������\����rTh�V�F�Z�����e����ZDHo�<g�!�w����Q�^�c_�>}]��;����3�d��̼C�N�L;�33moi�����������;4D�����eڇ���i컩�����]Zʄmn�D�7>�/�{TT��αa��<m!�@x�GT�w\�?�0!�\"L������wu2�03qt0��p��p�w�p�7nBY	�A��0���U�7"�3x B{{gkkk/OW/OT����,ۣ����!���կn����@��[��W������C�v Bg����V޾�^�n^.� ����^�ڊM�MDP�HT��=�]o7Wwg'''T{A�h?/�`��s�6s�����z�R¼�E�<znH�	/J��T�O�QW^����Cg����4M����U������UD`�J��_Eh��" �T_��KXBL�"�@lD���,&�`�����"���7��Cǖ�ݸq�����x����
����B����� �A�� t��^��С�!�̠���z���;�[#jF��<�1%��ؠ��ʖ�,�y׹���Ϸ�m�^���Tō:G�^���,��A?��hG���@N�Y�|�EJ˧��$�΢����q��[��l�*��W���� ����)!���$f��K���y�A]P��2�HA��,؅+��%hbU��%<E�k �U$���Q��Y
ؒyZ2�"��RNj-��	;@f	;����Ky�MM�a���S�ɯ�q�
^�g��πm[�. �S���D6e-i��.����O~�[ ����?��چz?SU/�nP�5+�ߪ��VR]?"��:�0z ��"�Eᮓ��R�ث��K�����ԇ�z�˖�u�hҩ�Y4����)�0�s_�8�>�����Ա˔	�v�����

(����"ބ��A����]##z%�94
�ԭ��02��Bpa�b��C=~a�s�Ǐ��+c0�b\)�Q������3rr�H�\t&B�"��u�����p��=lA�QZE��d��b������������?bgg���EW�;Z��;�y�8{��z���#���K���B�"dqx�S����<==����P������㢢�c�B�Ѫ�@��ߜ9�M�5~��O��L�~^@;v�M��.�t��u�w�:f�6A-"�GR��ץ�IK�OZ����-a������ ��qt��a�2xB�@�
�|�Ŧ0� ��y���"=�YF!p������J�(@ӟ�㌔AX�Ky" ��.���֢7��
�0���(�R��������'� N��&��ռ{o,�Fh���&I��������{��ߗZCjFbE�����CO���Z,�V�` � ���R((�f�2�(o�p�^�J-��#AW���O��Ío��Rr�SrJ�䢼2.�{YX����ZFJ�S2Ɍ\;��)�s
�":��-R�
�w�D`"d	5L���B���5"X�[8�����0���鰓_;��"ZV!�<-���,$�����.�z]�����RP�*��u!%��UB)$�uK��$��߉�XbɘD�/�Q�+���v"�;�֨�D�jA=(��G'����&���U����|}���E�P�3ȵ�r�[xu~��U+�U��Mg�6x����R@�k��"����.BT���.B��p��WPlD��ߙw�ɴ���m�v�jr1QZT�..C#�l�� *�!}z��˩�����t
�v�D��C�݌"�@Eh�.*­�'���3F��Ő���Eb��K���߶!����d�zi��2������xD�����nca,F����X������5��ÈW��o��_������}GS�v����Y��8X��z{y���2Xla@@�74O_#>���PpadHhtX�1ܜ]&M�2b���CG�~�2wՎCW�T3���?uY��zñ[�F����V*� ��x��֓���Sw^�;7/,f*��j� ��7"�`d��A�"D]�-(6"����b��L"��,5�Ij����{�9�^f�ӊY%��2J^	�/%��X)�����FDA�����U�,�DV�9G��^z�c�	������+�7�����W��P���>�������8�H�7o���G�VS˨б����1�Y�r�DX����3�I9��rfv)��h  ��IDAT3�����+����s�ҲKSr��7�ůs�^��.,M-E��e��dZ���|� �-"�ep����`ZD(V�a�!aG�*�-�ф��<�J���"�[��`���e��JA19�����,�d�ҋ�E�Ԣ���|ԅy EPcj~yj>>���]J-"�P��["��HS-�l��x�w��O=
��C+L
���R��T��?�iB��K�OK�9�
���S�`Wb>��+�	��`�1T�k�����d��{���s.9���j��O`PG0�	��,ؾz��xy���o���'`�Թ7�wp��k��_��S$%8c�Q��qkλč���1z��C�a���lj��^�@��6:
A!6eD������beke���1*�#<�%4�,:i�oe�4��&�!D�Q���0�j?���x
*´��2
�&�a��X+#������w����
���vrs���lgen@8��`����g����� :t07�ۥ+`ojfծ�u����l�M��\<]1�%��}��<�X�W��+e�S���E8��5�D ��'������L�����z��������� ���1y���CG��;�֣W+7��=ř	�&�����.`(��_��y��i~����7n���݇O��,+�,�s�4�,H�)����U9�,	#��z4��/� ����h��"
����#�s��l��3���.���t��XA`�P`%�ڂy����WZ�
��+�4���M\u�«&v�O>?�<=	��hC�0%W�p�_��OD��_�B�\��.j��#鲻����Ԁ0����D�ւ ������5)�"'���]L�m^) �`��BV>jDԅ���䕀Z�K�Ee��L)�D+�2K�2&��) ��D��<�bXh��c���>�m��a�@��
ON�(�	�-�1�T��.$)T@"�$V9��zE�d�a^1Ĭ"2�YL4�O/*�*��e�q|f!!���WJ)%�q4���-�s�J�Xg�ذ��oDh,��՝7�7b����f��1�,�7ə��F$]�lyD���e\��,��2��Y���=������@
�	�]������Ȁ5g.(x��@"&o�����w�����8�0�ྗ,�;��y��?s�T&�r)�2pf��Չvf���SzM:���%�O�]�1:�{@H������넦�@[�Vv0��Sǥ�U�H�~���8~5GQ¹Q��,���������9�F���c��Y�F;| &B̅�ą�� �,[H�gh�W����������������@���ν��LO./ͧS�l�Š�>��g����"l���h�D��Z[�[E� �A#2�):[�l���D��@7OGwO{gWK[�N�B�vvV�.v�^�~��������3�06$ �m:vB��ڙ:�X�{�8z��{{[���9G\��\��CI�!�CG�_�UP�����<rwwwss����x X!����EE�,Z�|��Y#�L9{����ҋ7��=vy��ۏ3��8�R����W7�g�9Ey�WE�B��ȕ���B��(ԁ�"l�`�1�`�6~@���T��B��g̾Ɣ��j�Y�R���-%m�x-��)t�@k�6uѵ��S
Db4i��r�5I���ɀ�&΄:3nڽ�3��y]��U����D��T9��)'r�	���|F}�����>����b�W��lP X0��
RlQ���B� �&DX�V�K/!B��YF��Q�I�
������ r��o&B���/[���q��Fx?�E[R("� ���D��3��i���K)@���0@�٥(��Ĭ"<D��YN��`�WE���H��|�V^�mxC�DNZ;wGv-R�����������2�:��H��={O��d���;�0$z��W����j�P��ת�E}�k�Sy7�N#�JdG��q��۬?Δ6�M:�?i�-J����ɗ�|2z�#wd�6$�ڱv���������/$:0<��ɡ�y{+;3;{k���:�!(мc;����O�c��C^Ӆq�+Y�� p@���2�'.�q
�<'�(�2}���N6�������C�u�����2����t�<����(.v���������	�N��vfN�qQ�}����eb�+ba6���P�T&��b�3e~��W�O�",��\&�Z���U��C�n1�W��>N����,��[[��Xt�8������p���������-��� ;S;ӎv��m��Y[�X�w�p4�p�1st�t�w��t=��+¿����>>^�~޾��h������@?oo_؂;'v_�z�̹�&N�}����<���y�E��"�Ô�G��yx��(�˸�<��,��6�ėT$tcBt�P۪@/Z�u�?[P^��i8r��X�-U����D��-&�DX8b��đX��i|�ÞhG���	 �X-�B9]ZE�|I#Ѝ�=P��ۍ�A����uخ2��T�g��#��k�ɔ#ǒ��W]��g�F���.;NS��[�u!�-EK<҄ ��r:FN-���UB���I���|Bj>>� �ZH�[ x <B�<���-��16�(� �'���1*+;�*B̂(���t��hq��h>��](�FG"EH � <�F�YR�(*��Q1���䇎c��a[XF.��ʩ"�$����B,��-����>pb�DX��V�"T�530NX�s���̷)H!3ߢ}�M?����t]q���+3/d�d����]�D.8�\�pT��Z�c���
d�=�+E����> �ab���'�4/EH��<����	�E��H&���A{�|:yK�u��r��6u�Z߈؀�h{W;o??wW{K��qʨ g�>����zC�>,�1k�_͌�<�YrĂ���0^rĳ�4G�`�&;�3�
�u��do��"B🃭���9lm,Mzv�2v��ޝ'��$�g�q�_"��K������Y�c�u�ϝ?�K�h{GS3�8'X-�d���\G�� [33���)� -:�`,ؘ�XZ�t�2ioe�ⴴ�>4��+����g/^bC�..Nn�.��`D///ooo��P���↮��	��Y�d���F��z���W���<L�,�n<I��BD:�Z@*�
�H�B�(����2����I���XZ5���l!z]��uZ�@�/࡙H[]��nb�A���?�� c�0�q~����[�����j���(����@�b�\(R2��Yc��3�ɫA��>^}��v,����Jj��f����_��@�B�u��R��gԽ�<#�.1��,��%�/"�3��B0tyb"�$���O#�S�I ����",��JI�"��P ��:� ��h+B̅�� ����ږ#�;R���hA��a)Ÿ��Q�S1��S"��������|Y���CF����x���L�̓)��<N�"o�]wE� E���'�e��]F��q&���DV5�i���?���z��8b�����;����h�g�X��M�{:CZ�CT2p��٢x��|�7���by�`cz���N�,�|����[\�������}<�C#��#��|=ݼݝ��� :�<�q��A�d����ޔ�G�M,�I�"d�"�;�`м��X�u0�h�bgn�d`
�v�k!v����%��=��;��+8�#����v�p�us�vsB� }�L=�{�aQ.��O"�~���Uk-�T���(:YƘ_��p�z�%��r��垽ڷ3��4qt0wrD(��-�m�\k �B'K+,.����¸j¦S;s0eG;���[�t�i������:��и���'3r�e��rv!�Q���)@�P�̗ɯ�Y�66V���v�6�����...���)�m����B��,Y9k�ґ�ݼ���̗i�)9���.��E�%���|"(��ʙR<KF���(?��-�������mS���~����;�\�-�G��~.[�ʈ���~R F�W�[P�̗k2�H�A�*�3e�dY3A��R�Z���-�ʮ���K�WS*��j��)�_ŨF���Q����DV�+X����-�j���u��%g1�R�B؇[���H�"������8Zj%�&����b!�[T��-T4��Αa"�Z�Ѣo8����T�t4!_E�e�����qD&Z'�,�1
pt8��S1�� ��0� |D��r*!@a+���a
�l���+��
\(���Ш��"�lw����	�H�u���V�lӥԕ�_�.�N�rtH}�T S�%	�&����#z'F����K_����ۃ�!�e����k��}8wO2�
n�E�����L��DR����V/ٗ���05�ƃ�G�>�ړ�K`h`Ll@TxHL(V}"&*$&"4:<$*,�@dDPh�O��N?|z�q����c��Z��dn���+"�
H��d��K#?s���SH�7v���/1&̗��������D��{��ChR�
L���b��D��K��KJY,�?��c�����Uk!�JM��J��+����2�E("ReY��M[Ϯ\��{���vff&�v�����.�	�t��t��tp��wp��s��u��E�Vc3h<]�\���<��-��-�]:ٸXX��Y��&��e$�0+���z�!ҙ,!D~�<�ޒ�����������������=4G'3Kp��_�O@Ȣe��.^1f�ow'�av1N�Q����<���-&�K�"<-��7t��%��E�h�K#?\��!��ͨC4��a���I��)F׶��0�W�+X��b!W^�S�
�P �0�~{U3��y3O�,�5 ,����QYM���+U�
5I�/U�4�̊��G��-Ă(��V��A���.rK"�w�R�!.�7 �~9S�gK���<;�@O+�fM�_E@8(�륪j��Z�AQ	.�fa"4^=UcU8���H��+��iL)�&&S &B�.,#��5��e�p*�<<�Q�-��O&����Ъ�8�5"Ҹj!K�~r�PQ%R���Y��d!��1�,4+�=�c��!�.� fm}Q&;p=eƦ����v����ţW�An�q�L[���u�ǌ^p�n&<l���&�^}�Ե'��9xkج�+�]�F�I���/������G J��r���ΐ��}�p�}ԁ�[��~i��yQ	�q�aq�X�������!V��[��<�<������:i��O���"��H��.�^tpٺ�cF��@k�c@� בC�N?bҘ�=�D���->
�{Bt�.�=�� ���u�����#~���N�0ftLH����?.ɡ��(�R�ߊ�˗o���Wkm�C�d:�uZzV^>H�pZEH�+���Uk�:8[ZZ�靸x����f����AD��`��rt�tr�p�ws�s�����Y6o������f��u���w�o�,"�N��5�_���ݱ�z�SSSS������-�jae�֬X�|��%K�L�r��ˇI�/��SrJs
�)�y��b* :4��n�|�cqp^/���Ml� �F�2�XJ�ѭ�e*��P!�ł 6:�O"d�tq �^��i��K���PDh�|l�}+p	���(T��"C���zT�2-t"�&�W���{�pY��J� cUIh�BJ���B���J���Z���mU K�G��K[����\T�VL�LU9ML��
SjL-$�*ħ��$V��Af���	���i@�����ӄ T S D��Ѻ`$6\�NN1�i�E(�7�&����(g��Y�x�.��A?�FT�.��)'sPi�!� ����Dh�`@ �f>���qQ"Ch���A!���"r%�_�P�1�k�r*�RȢ��S��?�v8��W}�����S�K�^z�EW7����M^��܎���&�e�z�Mɜ-G��v'O�5���=�!�?!o�X�_9~�ũ����X�f����I'�O�O+T��o9�t��m��0�?��p���_�_��ϰQ�F��ݢ�|��m�o���V".�I�\��;�fE'K�=�-s���:m|��-�� /gc��j�\�R�/Ι<vX��Ȟ�є����%�קgB�^��{�+�O���]Us�.5�E��#ܻ-��1#��M�SIt��/�j������`�LI5�#��)l�т<�,(L9�$��kBXD����3���%���s�:p!�������\��"l�Ľp��uU��*Μ�������������y@T�P���R��F�����--�}�|�|�X8w�1�'�y����T�˿���:�\�[J�SDD��E��{� Oi�F�iYA!���L̐�����P����'��b�r�r�Tɔ��2-M�&�d$��"R��*�HB�(b㠨D��7�EML�{*l��X�O��Y|-OT��|SQ��&աe�P�٭h5A�R ����sV�X 0U5Se`�@�:�B͗+E2�X*J|�����i�ru��jv���ױ+U\����f���ؕ���L�[�������`��j ��(��ぃ��8yZ4�[]�P�eM��iGoe��N׾/ޔ	d�V�v��˧E�b�:��O!r���j:��YN�!� R�x��.ĳd�05�Jd����PQSN��y�v�ܽ2"_(����-'
�O�R=QQC������/E'�2Eb�@B�I��1�4
�gt!u!�Ņ$p3�-t1�pE���I�ha���2�-�����k���]G���	I�A����o��"��R��m����"���w���S�{���Y�G��F��i*`)��|@؃W7��A�_�uo�w��..�nEsE#�K�4�����-7�*>i> �Z�_�h� �
d���~S��]�$��fǑ��� �ਈ��И��.�b�w��ѽsϮ�]�ccb�"c��|���w�u�<,ʛ"N~)����F��0�(\s�q��Kz�	>Ы�� �� (<�o{�A-��ƍA!8��� ~���>]`'&2pݚ�
�J/$����?̯ˀ�㓟�p�:��K��D��Z�z��"9%;��H�c�PZEHf�K�ήa��a�����^����U±��{���[u4���|��Q:�z8Xa̝2�V#`'��pt�r�t�2��w���.�MJ!�aK�	#���t45G!Z�z����z-^3o��9c�����y^���K�ƃT�I��R�2<Y���GI�&�-�5��R�
}hB-��ı+\C9[�M��sYL�����%�������P"�UU��Hƣ���l:�]�H�Ptj����]�&k�Ҧ���wܚ
�J�� �:D^��q�%,9UQ�־eț8��Tn���뤲f����)fVI�>Jnuͣ���s�=J#�Dr���SPxj��	ak/�8��Y���{q}������	+u\����	T�UG]Y���d^#U���7qt:a�'"��w���i����-¯���I��;����A�Wе%�
�%IXG��}F��*y�G�����X��[OX��i;�yКѻ/fh?�p�*a�E���s-؜����
�縲2�"���cpbE.�-�n�^��nƱ*��DT�l�>K5�/Xr�{�ߘ�:���+��*ޖD�ZD�i&K��2U��Y�|�ck$*C"��M����\P8hF4��"�aAlK(�b2�! ��Dz�QLa�P�<����L~K �CC|���;�j�'��ϕ@U-PC�W�k�p���F^�Z#|�1+���_8���T�bM�P['�Ջ���F�����l�Ï4��~GQ�N^�d�CV��(7��6�3���"�;��AX]ͫ��6|!h>�?�j����<ˤm�w�?26$6�+��;�+*6�[���=�w�ܽk������Р`?�~C�����Y)���fNz��O�+�޵��ӵgTL��=��o�o������Gm]��A.=vp'�0*Էk\8�,ثkT�n1}����׿W|���� ��gd��r�`vƳ���F�GuK@*�Q�<*�)�K���o�"d�9ϓ^���
�Mb��|!��-��;$��oǖ���?xp�b׸P'S[�vv�����������`������k �����x��z�x�ڹ�9aC�>A	a1��\��"lm�ML:Ztr�u���~��U[���p&��޳7�^��$e�J	R��LXNV���V�98_�T@���:���į��k��wl�7�NɿB����Y"�s뿊b2��ZY)�
��S^�򤔊f��sQE3A���t�'\Bn�e~��jp��ĺFz��$���*~�E�T���*��H�\����p�z��L��U����\A%��#��qȢ��c6��_��iX,��T����5��QD����7q'hrx���P���#l=R��@�5�%o�|D�y����T�q�������R�K$�+b�bU��M�dP��N��o��I�t|C	�ۋ��kI�,B#M�\~̼�,*c}-�0qu�S������8raF��W�L;w>���o�=�M��I��m8x�z�yɚ37�?M/U֖+jO=N����U|����+b	�-A�9�T�V���,|��
>uGx�9Y�ZU��Ӟ�Wx����LT}�W �K��ޔ��������	����"D�B��L����9��aAlK��;̅��j�R<�:� ���,������ B,�u-�P�o>��9_�� *��A��M�iE�L߈bh2��3����#�Qd��R]�Hfm���ɛd�FyE��Z!�Sp�j	��g�����âgY��{�B8����������

	�z{���fpX �0�����R�H+dd�si�%d����Ssqܥۮہ�u&Ą$�a`�.����-.."0��92�'<�5
���J�� x�ɦ���UbL����o^ҧWLDx`��> B\)�L䱘�_"���{k-����<{�_X
$�Y$��D�^�w�y�tM����`��fccnt�1�t���Ax�Z{:[y:Zb@�f�	�k���������������W`|Hdcf�%B�N��A��;�z;�Gz-]�`����gL��<�yjQJ-�HP@P�ʀRJ�UU�4`����G��mF��.}��T��xn-�ӈg ��2��R�;���)7���袶"�\�"U��'o��;��s|q=�`��Ȁ�wb�]�7b����1���q�R��7`�Iס�C������93x������I���'����־c�Ur]��{E�����:>a��u��>/��$`��ȡ{i��<y5K��h�ݦ�<~�C��;q�$��� a;����k���,���k���)�G�~e�✨�l�-�p��Ѐ�:-v�����w�|u�9��[Z��M����8�� �.|CP�#~]��Dm�6�G���^G���L!!��ԗ�U�������K~͑W�S���w�q�o��#u��:x�}��A�>!�������z��3ѣ��?�R�w�ň�G⇜2�F&��E�m�%q�-Y�=��L�5���#i�Tȁ�ʀ�{�,���1pءS/5WD�5]�-g��J-��l!l�L��Bآ;F9���*��\�5�6XP�2(j�"C�A�\Y��~�"DghW�V~�V~�U|�XM�i�X��S B��?E��m�PO���0V�mE��BI���-&B��I��W�dU-"�UԮ;�d��=g<�"n2�����������������������>������N<`�̒�"RZ!�*��QrK����B%�[����oOaDl@[&D��{���֬��I��[����z$`����с@|T@\�?�1�����<:̫[BP���#�tM����
�؋T���1P��5*������U���������t��i!�����������KZ6������M4�h���	�g�*Ј�������]GP����l�ޡ�������	���Ǯu���l@X��/Jr��y%��RZ�u����Jg&�J����78S4�E; �`l��,������Զ�)��M��w��g��G�>aMr��Io����^xϙ��]w>�Hy/��wܺ����u����=zC�Q[������\���"��%2#��?)ї�5�$������/O5�N8b�c�������O��?���������ӯ���v�z~�ce�A�׼����ܼ�����4�wݷ�<'�T��e�p`6�ggN<�1n��W
���[�.9N�*���VQ�_��}�����2zk���g�t]p���:|��	gd6oxR�3���k����~SF�IY��"�S����h�I���<d!����^z�c}ߥ�.d#�H���^�O�_���4`��Q���fE���������x���k
�'B�%�]V��rf궋�(�4��8-2gwR�U	���HԠK���Nی��-ߦ˪�gJ ��˖�++�#�_���Nic��W��v��-%]'_���8x��a{/Q׉'ݧ�=��#z����""~��F,�y<C��)�e๐	שUI����"�&.aKY�#���`.�-��b���;,r��x&��j�W�l�4h��?�P4�P��v�
�܆�������|���ZEX��"�h�>��P��W� Bam�מm���#���c]��M�,:�w�s�����w��w����vvD�����[ZZ��<0�Ș-��d�s�H ¼2B��W�]�W�И8aۡў]�],����;�";F��a�E��`D�xnNf�6���Cb�Ã��b|�b[DH�sI*BFK�_"����������"R��B2�G��(4iq��%��+-{��wp��.�`bz�����vs����;3P��	Z����Į��mG+So_��z��~ѾA=>/��g�3sK�+
h�8�,'�U��6��gcaj����9:]��]Ga�`��dg���n.�q�aq]c��� �7t����W�2o��y>u����n��N>a��VD��z�l�36�~��?����٧�7�����A]�m?Qp�jy.��,6P%
�T�)B���"�.aT�Hry}���|��KX��i�Y��uqk^��ܶ�u��T���Q�^��8j?�Lت�s.����Ѐ�L:�9�ZȊ���D,�6ţ���Eh�����=�t�=����'?�~i�MZ~3���m��;�U���&��7N��yBM�F�$�-M�0j��Ee_�����g�Ms6���U�h�dYǡ[Ɵ��W#���?�T��-y5�����ט�c��]�̚^�$.:�:tS�[d�U���M{�D���C6u���	�˾��甏�
$���a��A3/{���T�+@����j슋)��t��n��x&�?��u�Ui��#7���@�1n��S�7$z�%��;�&7���:�`�)ԣ1�5H�թ������:�یێS���>m5�ҒWuf#�Ͼ��@��H¬t�^'
%_�2=��b�w�\�v��K!.$��7�b;༶"�X��"�DD�q�V��!D'71E� [\Õ����R��Z����Ӫ�?�PxҊ���ȩ��@m ���@u@U��`J��N���ѥ5uc�;��3R���-U�?`����w�� <GΓW����|��NM�'��JY�� �^��,�ճdz����=B����f�@/��:=&Bz��H�_w��U'�=.|�O;z�z@d4����y��h=B�N�f�MM;�'���w�����l�CC�"�( p���B"�0�Mă���s�/?m��=82&!1]�/[�-:�i۰��A>��èPo,�6��p!��63i��$:�%�"CG��D�,j#�_C���?�#B*��s��Q:آ"�l���ɪ�ʡɐ�`k�Z�8.��b	�����6�Llۛ�u2�1E?�mE���������zvøΏ������2<@�1�'����rvvv��wsv�T����P��	wyz�z��y���n��]B���v����
�ced�5��&�0n��=���]x»�Wu"Yf�y��ܪ'�/����f��r�4��T*E���w���=z��$zK����04*6.V��5,��%�/[O�ZE.u�w��$�!�-��v�:y�D���o=���K���9h=j�س���H��f��8N<�{{�I��!�"&*�"�*�X�(o��)���0��e��v}��}�p�h1��G��F����W(���;_9�H��&ds�p�ꚗ<Ǳ[�O�h@N��ڌ�4���)W��/?��dK��n��zٳj$l��!뎕}��o_n5Av�0���d�J�ƭ~�Fzn�`3x�s��>
��s�k�R������d���;�,����1����ٹ|d��[f�#�ds�ߡ��;|��g�ǅb�	�y�+a�â߯d7:���{��M��]6�ݕ�,C����y�L��ч#gH�}��S��~o�늁�R]F�$E��_s�pmS��I��n�o' �c/�L���F����w���(�}b*kh�4�+���G4���9-�_!:�Wl`I�ٲ���<E��⛪���I]�UV�N�o�񕕺zTi�UU�E�<�"@W�A�����oB��_�mt��+� �U Qm�{+"M�GDS����y�ԼG`��/��{kx�	DX��wP#Ěʚ���ߔu����Z����P� W���j�A"d������v��J�y6��ś�y��BD�B]ة�	V���fffacm�wࠬ��������|�_E�l�%G�=��߱kÀ>]~'��\!���#�=��࿸H��(��h'��N�&Nv(`����H������ݟ�SR�pu,���"����W����'��˨L�� �?����U'�*��y;8�AE��hx;Z��چ���x9y9@\�Z���]��C��^ �{�2r!"d������S�np��1�����`p@PH@Hh@H���OhL����]�=L��M�1�JB��#���6���O6��x��u�%�A[��l�>��'�s�5����˔c#W\yJ�%�r�ｧm��D�K�$�d��* B�K�Vģ�et��K���ϲF߈��k�QM٘��y�������-�{�3�n��~x:�ʥ�v�Q{/����X�^�>j�BsȔÎ��.>��d@v���v��J��݆��}Y�{�k�돔�-�/�x���)��'�Z{�ހ$�}�3�����%��\��C��5�v���I',n{ ��M�ߔ�E�wU~�����kDz�?�0bü�偿J�B�2h��95lo���C��O�6#ы�[\�����)��o}ɺL�u�:~��g��c����t�z��+�7�O���{G���y�?BG���Ƿ����;|�LLƩ:��wc��^�6|�=i'��Cf��x�˲��z.s������]�k�8�m��Sy�a��ڗ*CFnɋ�z+~��v���f)r4Y0lw�'{o�J�y������25K�`�U S�dH�(bK$c�� �'�pyd6����,LDHۂ)�d̀��>�	Ѵ�4�� ���)�f��S��%�Hb7��u|�G��bD��(\�L��+��B��J!��`Aye��Ь4���}��� �k����?�/iDx�f"��J�#�.��c��_���*��R�kG�jx~0(|D� �䫫iRK]�h�\�V@���$S5I�U|���
j�
��3r�Y�yn�&�yU��ع��]ۊ�DmF���"�7`Pv~QV^qNAYv.��	g��g� �[���_�������Q����Bt����z��&° �����%��c�o���"�6u拧�y�����P���Y��o�_"�W�Ղ@[h B�J!�}�,���Шg0xD��h�h�	��d,�"�"B4�
���Q��A�Af&��&�&6�&�^#��&�}������\�mE���*����� 4�``` X08$"8<:8<��#(4��0�������GL\�=���_�u����7�f�ڼ�|��r߱{f��OQ"�ϗ�%�O�t:M�;x��3o
�s��������z�L�ZP�W���҈�jD��8wѩ��6�)j8y��s��mgs����I�Σ��>��P�u��#�d��WY�'o��h�Y��5Ȭ��z�����,U5�8U�܉7Ŋ��ς���O�_��ZNNr���k�A�[d���u�λx򔄌�Q�?�b��{whdi�K%�cw���z4aƩs�U�zd�R��Y��qC�i��>d됱��^ufޱ����5!��M/_�����vܺ��T#[�&��3t����sFm���Y_\�\qbΑ'�w��/�o��&�|�5m����7�[p�	Y���������O?�g��A�ק�ӗ��?q]�w=��ۼݫo��h�������3�3=���f��[��v������|i���A�����B/��=י�7����U&��"eR�����/:�*II,k �u<������%t��q�a[Ry"��$��!Bԅh~Z����������g��<$��O�Ý�[B��.k@v�~z�5��y_�U�9x�nZѨy+��&��=UYW����w��ib����;�^ڊ�O�|�}�H��1�#~[��G樛g�o:�}��	�6��c*>�ߎ_K1}͈髎_{I����W�:Y� Dq冃�n'��b���]GΚ�z�+��TX����0*�m:�O��+�Q���r���K�KO��������g�_��7$���!ʏ�֩����e���"$���\w���^=]��DN7l���ƅ�x�����>��B���"���`א GT��Naan���a�������ԅ9\1�N�1�-as�mE��H1Bh�D��Z�z�����%%d��`�t!�D�q�C�f�ި�n^>���^�NNNfV��,�m6�@�h&��`���ao��h�&u��`o������������Ƿ����{�0���_��/�a�(�k�����^�A��A�����B��Cãã£:���Ev�uh��SN�Lw��̋"���k/t
�����9ڸi��2?�!7-<��=n��R}�܃#��8�{!W9aݮ;9��\AUߩ���I�p�$ѓ�*��A�&��wth����`e4i%_l@'JHjY�z���)}K��ty5]^��K�AWE��E=E���4$e-I�HTo��x�[�ƀS�I��T�x�"�@��[��F�·p#U�{*�F�'��Q񉨀G�kE��h�W�ȫ ��oY:����:�x�e5I�#��Ս�[e}+���W�iї��G�#�@_�
�I���'_�(����L\����	Q��$��i������}�w�yKW43�ML�;��#C���AX�?�b�[���'����TsJ�\�er�/W�"����ɗ(t5M��*ˊNdK	,	�)�h+B
OB�K��<�T��*ӑ�E��-G��>�<�1y����1[oR�!�2����^s�Є�y^>l��-�b[��Z2���"������X��D���M'^�cG/���r���
�v9�˄�����S�V���.,}�v9���M���/��l��BoJc4N�t�^��N�c�&��H�m��+�rEÖ�xXVy�@={���s���)2xљ��[n��8MH�nܮ[�#7nLϹT=���K�v]�4k�op�O@���m�v��¼hP���rl߱CӶ"�-,G�3e����O�����~�2�������}H�'Ă�c���=�m���?,�6l1Z�`���[qw53�	pv����ٿ��@�!�S3ߨ�lF�,�2l��+�������!$�U��W���ὧF+�"D��yD��LW��n��9�{�u�t��nok��������`k�dm�di�le�jm�b�&u��CӍ�Z��X ����f���h��NvNm\,�]�]�@��.� ��B^ۤ�%z	�
�]�Bc�"����F!���!��0�?!D�Aaр�d��cz��uФ��}b�/�y2����F�:a�ugod�cG��S(���m��r��{��u���{��~SF�؟�1
�I���3V���$1�%z�����V�ߓn�`i��,9�A���)�3�:���W�K��FT����������$L9���m�]؃�+m���<�K����Th�ir-Y����d���VZ3ϡ'?=�BÕk�B�S�p�M,M3[����h�������
���Er�v�|cRlW�V�'�L��H%�-ǳdpG�(B4�|�?r47��̿ϪLZ���KČ�g�+��z(���j�)A�H�#��g.����%a��Y{ �!�<u������ub��]��W���6aG���"	3NDL<p��a�����ɍHq%R�C&�J^v���i�e7����������\u�eKk��y'3��v]p��)�AR�[��9�zi���Ł�W�z��U!p^��R���;��\��O?��j��=���]����l�h��jk�`iie��f������ff����?#'?-+�(B|[����x�}zLq�4ooen
��-���T_�pu���l'���V��,M [s�򊹩�Y'ӎ&;�*����<n�m�^���3_W�f��*
MJc
Y\1G �I������j!���3i8�l!�)'P�[�]�a��%+|���s��&f�m�;�Y�Zuloabbݡ�]'S'K+ ,�dm�`��!�{;���m:Y�Ot�6iom��ʺ����K佇y���rA!���%4�s,%2�HL�I��'�xx�9;����@@�������B\{�>��o�w@Ą����X�c���IY�&e�3�|W���DU/�i�0�ɥ�����f˅��r9���P�e���z�����,��H�
��@���g�a'������E�p!��rxb��@l�-���~�U�m���o�t�U������F����*�R%*�H��q��Y�|u����.B����䫫��ĵ��|�Dȁ{����`�S�x�:����Y�F���/����jɼJW��T��j<K����a���n�H+�?�Z�L8D͚���Е�#��<�$��w���Y�y'����������wȟ���Xw/d��ōkﱇly�>zw�Yq������c��=�?ޑ�;���;�L̢�'K�����H�����!~C���{�-lFF���q�o˫�R�l����'����Kߝ̩��V�;�� 	��p��\�7���?��R���x��J�����}^r�6����ܚ�hcd\���hO?�@������� _7wggG81uCk���?سw���ܔq�E��brn	Z�
�]����k.�N��6�� G�v&&�^���l�L~a륖Ę�V����HߨPϐ � ?{__[__�JL��#&�_fk�x�:3�MEn��A�`sU����S��_"������)mEXN��z��ų�/$v��I��vX&7[ +@�������ao�ng�bg ����-M:�6͌ŭ;�w0w>xT�W(l�хh:�"���!P�O_��{�;8����5(���}|�@�`Ate|�����D�[�v��=�}�&�֓7�_�d�R3��/�)\E͘��������rY�"@8��ĉ�tUeC���SVM�� 2O�"h�������Ъ7L�?=��^x$8Bd�b���جqx�S��v�1���ʅ?j�(J���Q�+�cC�?��?�F��
 �-���\�P�1cjG��Q},���P���;w#o܌�V�+ VP��dn�[G���8Ue�
<S�W�����NѺ��WP����t�т=�h����$�Yq!c�ƫ�㷕�eg�.�1~?�9�������Δu[|����]Y��轩W(�y���yWO����r�I�Ɨ�]�$�,EW�X�HCE��H���p�}�Ⴏ�h-�+t����u�U�H��Y5H��k�X�������g$O�:f�}<O�a�|<k�l
���GD��i���3�X{�:f��[%�ߛ�tKTB���؀������=z��ҥk|LlTxxhhP0X1((h��`!���F
g|�s�։�%�Fٚw� �@t����"�r���p�q
�o�;�֊��	`ؘ8����������Mb~�6#�Š����T&�He�����)����(�uh���/#���<A��ѣ]�m��L��d&&���fL�+�^�N>N΀������2����45oob��Ģ����	�����ܮ#X����/ >8����� 2~��%8F��EDA	L,~�<��3��ѣC'��f�p��U'K+�,-m��LL�YZ������N�m��K�����"#5_B��.��U8��_F��I9A(/�J�2])OJ���|�D�QՉ��LI�Q�R:t����fy6���[u�?v�����?�+� Xev �;�Ex�G\k�k� ]V.dI��R=Z�I�u�-����H8o�ɂX�OU&��z�|o�|��A}̅���t���F�Q*k�:����h��>�J&�Z8��ݱ��n<�r�̃+��f�>��5�4C)���QSR�UGJ�h���
�ha�@/�V��J8�
H��Bl��c6"�:������tܺs9��K�.]gO�p�T��y%�=�d
������Z�g�keM	�N��!ǲ����߉C��J�#=V>��D~8�1~��3ş��$dڅ���S��ޒ�W� ���Xs�}��5z֩92x�r��&n�����gxîk��g�W 5"�B&�ڝ����j�!����-7��]-�����]'/Z�'"�;z�=:&6!�s��D�]�&����FG�DF��B����W��S��]M_B��8��]I4m��3�-[�}ؠ~����a���>	Q��t�}��	��Aq�A�}����u����G1������a���9!01޷o���}<����]���~%��P��G ��<ٯ��W���_��C�(ʉ��.u�6���:,�+!!��ۡsb���uT������M���~��>������^�h�� ��@�`?� _go?g_O��ç��7%9���F/(綈�}�)��
�B��"y�,��=���D���z����Ԋ�����-l��C�&N�;~Ƣ~ç�~�~���;I9ϳ�O^r���O3�=˂[��<�,��^� w/w;��q!�O
��^f'�^�RJ�ۏ��6xjM&P�%��U�PQA������������*�n���k�_�tv�N3�գ"���P��^�������BtP�-X�O̅��F�?��� ��.Զ!��Ҁ.+T��TEs��a��7k?Τ�MYy��En��O\r�,~'�!R�Q#x��"VmSM�i�ʋ�� �5X��׉��N$C��6pN.�ZԄp�fr��J$���>o͉��F��:bѾE{�+�s/hc��.��k��E�q��s�[��R:�yB0�O�V�F~��`�E*d貋����zd݅�!K.����e����UH:������Χ��A���[��v!Y������ߴm��W�Y�E���Aj>!U�ȼE_$H�M�We#2{���'S;�۲�Bơ�I�6

�������"���ju!��"�)�?��(�s�q섵�ܿZq�(��QXf�n����������[��B Ыk��>��1�#���r��^��$Qd�J;�m��=9Y��<�X���������-�������!��$ReS[����3��)��%Yӧ���t	�/&BO'О������������<�{#�MҐ~��������
���		?n�𡳳28�yh�	a��G`��yyxA>^Z�������8{��:z�35kg֡�&B�:�377ZXX���[;��;�[�QA�}N�x�u�o.�����}tH�i�D�X�y��ޓ�w��&qʚ.36$��7mM��[���;{C��9�f��p������_�wy�⸕Dt�j4"��M��Ycz៺r���O?�����w�1N}�N=�����e�,i-�P(��!Bx��X�'Z� "(���!W^�Wڊ�/�@���j�F%�hj�@��++4"TW1U����������w�����.>�n@J:�Y~�y߀��	��d��3<��䚚/`>,`m�X'���	�:�P+�(	����s�5Ҧ�Ym��N����	j��Ua��SՍ�J4�6�)���H:YN�~������)�*�@+4����Z��Q^�M����A*����$n ���OШ�e5B��7~C4�W�����i@��OR��b����+"�U��мk�fQ�{i�7@�m����O����k��U׿�����GxDԌl���0z����O^�O]|��}`dlgT�F�������[��]��!Q����!GO�ݳkbx���>�����E���3h�%��#�������5.�_ϸA��taL�wl�ϖ�E�b�&O~��f7|������2�'�%�_"�W�߈�@(�����]��܎٣Q�+esfN��log�����D8قA���n��y{.�T�W�=��5��9��) �) ��/��/��/(4�ː='dgs��2fZ���1�P�]
"��㕥d̓gNn!�.�L-ZDhf�݅�͌c� � �����s���dݰ)o'���^d����q���̆tvM��)[�)E�%E��Q!/ed���P�-��#����&^��̊����n9��B���Kk��v�m��W����O3N�3?���߈��i0Z����`��x�W~�+>�_H�OT�;���+��� B��~eT{�k�m���[]�����@ԂR_����D(T)E�H������j��� BZ�q3��֖�ޑ+?��a����K�m=�x����d�Zzz�����=!�����a[��Q�M� ��A��B �3�p�T���Y�
������R�'Kk�w�Z^e����7���T6����Y"yZIYۤ�m��U_~��k�k���l��yg���7|���R]�-7���蔪�"q�L��ЄHdu��־U� ��Qkx����ɗU7����\����)Q��5�������T�5	*�T�P�ԪJ��N�z/�DXzd��Ԟ7�����A9s�qd\ϰ�����Ȉ踨�bbb�b�"�#"���h�@�V�᳋�Kn=��8*16
D�=!�_���C�A�7�Wg_�kOd��	�3&�	�r�r��q���<�O|��b|}����E���H����'t	���>tbN�����Y�d���/��k������ET�L�a��)����ں���>���+�|�4&�߬#�t�ު#�u�����s�����A^�����������'��NN\�,\<l�3�������u1�������r���*(c�_�0Ӌ$�����ջٖ���6�M;�4� 5��"�����?,"f�����,�7f�ݴ�<N����L��"Q���\�s·<��^m��Ù\�s�G�߷$����3�'|5Rī�s�D�(گOʥ�-�"��(Z;ğ�:�`��S�J��[e ����f5ZP��DȔ�ڷ��+v���ϔ�V�}�f�5�sߞco�����'�:�{�IޔHX�F����N�Ao�/��7�1b��O�������u�95�:�(t �ߊ@Z!�V�5Y�@n(U�L����J��R���+�x�*� "BM][C��Ѵ����$ၻ)[.>�~�e�IK�p�~�4��%c�m���a�Y�F,<v��M��Z����/� ��
�X'���8�J���+�b�k�:I�7��P�V�����bCJe�@k�� c��ZQE���^fh�TMhu��z��N^�^\�NR>�*?j��ZQ�޵"�6R��X�@���CTY'�$za�V^U)VȔ�Z�QJ�ri�H�$�#<=����S6����2"���a	�AQ.��^A!��a��!����Zސ@�!bA�/ �g߁`����  �J) B��N'��]ɴ�ۭ_\T8Vn�Wטαab���=��F�z`@\�eň��tu�;g��M���X�G��=#���ds�,�Ĉ�58���/�~��+��/�j��"|��G�A!������=������mP����p�fa��aj!��pB�����!���^��NƔl����;9�wq����"BG/o�T��R�sʙE�̂*�ܝ��oy�L�p�`撣��l�?lAw��v���aKP���C4�!�������{��C�N��;�ie᮳��>yE��N�2;/8��Z^��T��Z�(f����������:���r=��+� �`HtD������\>n��\n5K����*¶���ۂ��Wby/���߈�,�^����e���oȪ�[O]y���g��}�]F�/�+�}�'���kή��%y����!Û ������%5|i�@V/�W�RA�P�*ZJ a"dj�"���5 �2iե�Ev��:i���zN]����Y4�W4��k��]|��}|9����s�<��xmE,� ��ƃ�j����Y�~���3UT�~��Z����+�U
�\kP�j�5h�=�C$�S������FMe�V���hj��V�@�C1����"4�a�*k$z��B�!�PKtJ�F�Q�u
�N���
y�R�u��/MZw�AfR&���۾A1~��6�V�6��.^^hbO�Ww����7"���2zTt�>	1�1�]0�� ����"cB Ħ���B=��@d�GH�cx�������U�#GC|�����5-��D��JK�K���o�6DX��"�i"L�f�L�}�"���#��;�+[���֝\���%�nv����6n�V���}�ٮ�9����t��m�*BWw[O4"�J���uIN)�ȕ����ecf/=s핇%֜_����Y{��]�����'���m'K��:Z�t47�h�DؾCK�_KsS_/o���㇎�"L��=4kۙ������]J��Π�'_Q4��ʓO�x��n��w9߆�z��ni*������y\��,�Pt��cם�ᵈ��EF0�a�����n���P�V���?��*���Y�w37]�!Q��\�!����ｑ6uÉavf�şjr!�;l�'YB�����1�?���F�?�i W�xb5�;-(TV ������/�� �'��ɫ�+�h�*T��&����l�)k�� *B����m��j��lL&�מ����S��O��(��Ͳ�Hq5r,�"d��է3_I�J8��ֹ�-�q�- �V ���(By�P^'P6+�7��$�j�N���P�P�Z��Z[��
�Vg��T�J���B�ի��:��PQS�C��V�R�1�R����F?π�JC+�P�"��:�F-�+�5*y�Ta�괲Z��w��{��I�.�O��?q��0 8����Ĥ}'s3[[k;{[;���-ck�u��!�\�"\y>�U�}�&������ \, /���P_��wz��p�1qs���i��hj߷ohl�O`��0=��LqYjK���_"�����8��ڈ�A��)B�T��{���}��ڙ��Ci�ɘ�������\����L��: �`?�~�����>�.�����.^� Bo�����O^f3�bU1��05�'�����[��lbH����W'�p3G3kKS���Ḽ:�Y�7��hj�q���9�����M�6s�y}FL��Zz?��\�`���S/g����&�ͨ,�6�^u�j�P��Ȑ-O�a��O�*?�Q25W(!�$����?E��P�O"�ރ�!t�n��܅i \�]��D��'����*B��7LY���˴��?·߂V������zMݰ��ݰ!V�zE�A�d�B���|6��CP��b��.B���J��R���S�{ 2Z�:�}���D���- <�\�V  �QZQ�Vֲ�e3G�#��n�M<�[������h�8�����m�k߳�_Ћ�<�:���V
QR�Pd��:$�y.E�)�x�,�P��"�V���m��|m@o����BE�@U� ��NY� �UC���U��0@Z�<;�:��@E&SEV�T����Fb.�D�������p�pP�U��r�Rޠն�T��=�b���`"��BEhm��l�;���gKN�N�(��2�!��ze���)"\z:�<rxL׾]�c���ܯG���t,v��c�-�'�x�z�$B��L �LZD�'<6�/$ȧs\׌�b:E�eiY,�/�j���84������d�)Ä���eew�@k/wgOG_{�vh)	;3#h�NN��̜�- �� ?oǰ`O_O[��&�V(p�耊�����������/�?��㤂�"z>��M�>�.�=b�����b����SN>���C��gW;�K{k;;GK;'s[����`g8;:y��O�<}���=�L��8�ܳ�QK���~�ˤ�[.%�$��.ٷ���=��-�W��� ���t���~+�L�{)�X#�)�\�-�)�o�G�=�ͭb*�G-(�cq�_�q�@ѕX��t_�.W�Ǡ?h4(��'�D&¶:D%!V%��R=KZ-��r1��״u�^�`Y�{��{o�LXs2q���v_ʒ�u�;uۣm�
hJ�%� "�P�σ�?��83�e�ޡ�E:��a��J�Li�H����]�h��g�}Ӱ����"��џ,p�:�J�Vk�jN,��+��/=)�� k�>4y���׈�z��#YZ˩h�隸�F�M�*{�q+�J���P���=vo������{������J\xݢ�:��L�$�}�E��i��!x��b�A��S�z�J}3�5���|�(rM�����\W��A�X_G��`_���?tEͻ��wB�������-�)U�k՚:�,V;6O!�WJU����+hOU�g��*���A rmhֿ����QZS�T�4o��}��I��\g�UI�R��P�V'�4!;Ϧt�����Y���@D�ai刉Z{����F:�4�ED�'v��+��+���2�N$�aׄ؁����a�XΧm:��������^���N����n1�� �@ "�=��������48�&4�.2�9:�7,����3/��A��"d(*��}���r��j��aK=B�wr(T^Vv��IGWW�UOW̅�&h1B��ڙ�`���������������������=|d[Dh�;ao��su��*Bw�(������SJh�)Y�䂈���Z�9�7jV�����Z;��9��9y�9;9��:�Y:��8�ٹ�;���ioO/���mȰQ�F���>���7�_�~���f��+gm|�C�~�Y��U��}3-�Qq�Y���K�����3�T�K�B�@Lf�J��2q��<��G�X�LY�qZ��HZ} �c��/�k�'���oDHW4��kןz�_@�Y=&�?p;�v��V�أ��=�c7�t�4j�V�ދ���D�!B�[E�*���u��&lqabSR�7�$�h�q�b�Ղ�_D��I�?])l� (��Q0�
�LJRN�͞���$���_��C����=��-�ʲ�omD�6�,>�0}��]�^�ɚ�x��{7�ͭ@n��⦝�v�h⁼w�IE
��ÿ!z��R�^�T)Ej:�����?�%4Q#[�N]�!�7�ߋ�z/m@x�o�F��x�x�T��f�aV~�����j<�ZU��t_�(��W!�oA�P���HH�'Dр��i����ri��#­��׀��!�O��=B�|[���T4��"��������R������ʄH��r�(l��+I�/���.�	����je����� �N̀�����������ZG���3���Q]����9�_w� WoW;'�N��=���l1��;�$���� 7L�>�F:D��FG�G��=�(�H"����/�j�Zk0��	*�C��"$�� G������y{�b��}�!.tZu2�6m[�������i
����{XY�G/(�X�)BgWK'GwO7�H��.���摓�Jo<]ʑ$3��7_07�O���~����tk�D;�p'W_'wWw{kWOWO;wOGwg0���������������#��c����'.
2s�}f�[��LE����\=y�3�$���|�I��6^��1gǌ�$u��+��X|]B���#���d��-�C��"l�A�C�*2SDf
�C�HԠ��l�h+����Q�F10�8q]�����¡�w-�|}Ԭ���n�6y���}����Eg����	!�����k�� ��
4��n��J��@���s$���*Bk�Hu4�:}���%y.l#B4�v*��^������R^m��G�����#e��2jr�����e5��j?K���t�B���&��Ӝۯ�? �?�A������տI�"=2i_���}3��"��O^m��X�'Gi�W�Q��(�@�S�}y�M5{��G'�8����'�K�%�H������f�U���!7�*�x��Z��]��H�a�C��(�~��ۄȾ �?M"տ�7OZ%~�汫.\͖*�R�d����c��Zx�P2��)oD�z��~q�䍽��dߘm/���5�_캑���,��M�'�Y|��z���������?Iٰ�x*B��,¨���ظ��� ӏ�p�B";�,EE����7���q؀���Ĉ��u��p��r��s����rh+��0 :�-<��O�ۅ�D�yFGGGD�>u�����C�S����DUN�aC��D�����"�2L��Q��>�N"�-Y������rG�q�������ܺSax �>��~n�>N�^v޶��E�hm�`i��v���d���h��\��O�͇/��gn?����C�,�zx��3sW_�;fOϡ;f.��k�Z�. BGWw�V�y�yz9{y��z���x��z~~~�~�1~��^C��x�v7�l̒�C�nZ{�֣b���������d�(�(̦+v^y1c۹�g��$*�JtH���,)]��y�d��S������H�J�w��w�z�@I�I>(�-����d����V~m�O"4
��0p�Le=S�T�֭�}1�T|�V���9)��kϋN?�]��궳��*t��>li�\>�]�-u�R�X��WS�
��ī�=ETAע�:6���Y��B���.�Ѕ�q�����"�~�_��ʚ�xT ���q�YW�Ϻ~=�0l�{tQ�W�������z#�,Eձ�/�}H�����n\����m�
9�O�ug�5����s%s%U�Qg���"Ԉ�F���D-����oW���;���p�`��m�C���9�Yt��k��U�y�Ȕ�)�.,�E�yt_���I� q��'�>��BR$����P?EO?|,M��DNgiC'�M���_N���	���;a�R�	���<��iĺ�ٲ�y����q���!���Ï��/��������3y��K�o��_ڑ�n��u�m��g�8r~����-���`'p������ۃM;v®�GF�S3s��Ѷ"l�g|"t����h+®q���g�}]�a�_���F�޶A�A�A`�����Ҋ�)tQ�d�[E��Kp��?�_"��~hl���O�����<P &Bl���aq�[w�<uV\B���P7W/{kGkkk{w'4����s��k�J��S��|��`/[7K7[kg���9��8�YA`��k�~�V��7E�d8�3��u:�߸U�Gn4�@�{���O71	21q��wwqsus�`�ֈ���(+F����,X�d�����������Wُ2K_QSp�"����#���4�"Ϧ�sH�"���������U%C	K���IX<!�%�~<9G0w�1�R���H�L!X!ڳ�l�B iL��>�%�n>��o��'�?H�?��yER�\�.hB���9q����.]X�d��募]:�����ӗ��=K�j�"e�
���O�D���2~,��)C�в��a%EXUJװe_�j�)A��Z��O��X�TI-]^��C�^��c���J�]����k��m������@���M���8�2�n���̞��<����=��}�,��@���Ԫ����-G�Wr׭��|~!��|G ���P �?p���_t�w���)d��
T�F��wf�C�B�^��iiA$�W����hcHUEk?�j�Ȓ/���g���ney�ߵlש�r5E�2~��#ϰo����Qk.�{^BU���LY+S�݅0�]/Bx8T��I�<�\(����#��E�J��{Yʞ��
�B���՚�U��}Q���uA÷?����4jW�BɦǍsNM8�H�
%�>Gl���v}'t��w:���Y���q!!z�tWu+��|��17�dYB�n�
���>��]��!t�u E�X�3Ͼ�^-z�m��tM>��\&�->��j����\�~���q����)[v���G<#C"F��Zh�hke<d ��ݔ##�`Px䰂����F�o���d��WS�B�����45r�2]g�����Px΁+�!|��b��� Ӂ&`�	|>�;F�aÅ�CBBV,_��9<�II]�������Rd�L� 8\1����×o�D�����,�W��*Bp�n�ӈtމӗ7o�w�̥�c'����[61bd4h���C ���=�G�� {S؅ ZX�Y5�17��5��r�yU���)�UKfԐY�ٕjGQ���s���ѡQ;�M�gl��?�����ڪ_�.�6�"x{�{{z��s��e+�O�9?�u�������\)�^�e�;zc��xP`-��@�")<$M��T"X*G��*�\!�˥r8�)�,��o�{�P��=S$������g�u�W�w��,B�@��D�����/�b�Sc�D߸tn�����ެJy���2%\��_�\5Kܡ�kToA=�bA���;�CȻ��9-�^-�j�A��drT�X�OG�g��-�rkq֜X����dv/[�C���"�Kԅ���_!ໄ$@K��ַ�>()�p2i剴m7+���:e˵�R"^�*i��E� /1������Pc;��z���L��k 1$m���E;+p]2����144Y'C�ʐk����D(���R�X&�x�(�˹�v�M%����5g�f�}>|���: ��tO��2ḫ�x���U�˔����'M��Zr%�h*>r�u�h���$J�ބ�=��5��\Y�A�b�3�6b�5�e'������ю��S}n�Wh!�{�A�N<_q;;W�G������g^�J�_#�^L&�C}�ΔuN�X�2�n1���畋^_��lPԸ�c'{�{y�8���yx�9�:;9��Z[X������ aNA�~g��E�AQJ0��}�m5i����!�?VM���z:�xم�D��- �&���ca�������������� ���9s����~\UWц�}K�~$STd�@�B&[؄������`�y�:�����*Ma��>"q�F4�ȉ�GO��y���	�#d0`� �!s��p�1s�6s�1q�2���r�����|�����������������F,-�݃}F$e���sj���'��@�7@�w�݉3��4�MN����6���������������������������QW����EXX�+CS����r#.�TOd!Hl���r�i3S�e+	�˧�$�b��Z�m��qTr�D@p�E����Z���u�T�����_�~=��� ��%�r% ���xv��ٝ'�8w�Ĺ��O�z�܋�8,�.jmh;ࢵ�V֟e������K�$b=��!�	�]�"�3vֺ����)m����s�R�[�ң2y-���p�l\�k҂�g�O�' �O������ߋ���z�����𰰰�pp>R��ԋ�y�o�q��~x�YiB)� ЋP,ȗ��r%@�څaK�+��f^xU}�e�'�^ s��l��˥�(]P9�}��]�LE�CS�ѕ-L�a��*���6+O���B��T$�	%2�P��(������a󏾨V�ի3�}�^$�eR�]�]v>���x�h奬e�3�_��)��O$�%�Go��I��LS��L�zX���0��A��OW�I8�'E�? �W(��3���E�q;�'b5��.�1+rؽ%�/y�wQ��-���O_r��ٗ��o�ݿ�G��@G���o5lL��/��/�z���z:�z:;8�{{�z:{�:y�� �89����޾@�Yy�����F��J�{��Yq|ٺ��+�[���; ܝ��������� \u��z:�:��X�Y=�>��N&�v�����,;8[;{��;��)��Ӓ�j�����"S4d��g���\�~��W�K�oD����j�=v����;wxz��E8dȀ�0FCt�f���0��r������|�dd�hl`g
ϗ1�20�2��t����o�W��䬺�Ihb�
�	ϳ*V�2j�C��.H���2�cl,��,m,��XX�Wk�Hikncefeafnjbie������c�����N�1/!#�en��Ƃ:l�\���c�@�֡N�h2Ca�+%�<[��I\� �GGs�6����Y4K�R�)RQ�!�"T�
�j�P	#P��Ӆz~7_��W"�&V�9|�RE��RE����8�$A(����2k�l�ͻO��.�R�W��p�����r��߂L�  �
��D��^<[^�����
%�ʠ�yڙ�aY��u��;��ד��Wq�Y���w��� *��-���:�A���������� 82�B�<�7v+�,���k�=O��z_ͥ(?�T}\e'Ho:j����JM#��Yt�a�����N]�s����,�[q�Ҷ�O���>έ��������-Q�CQu�.T����E�s�w�$B@*�K�J���#����^Wr�-?YB۠��o L���+�xN�q1����Պ�m�z,���=�:���&�F-?��ҫ\jW�½����1��^�J�aҶW^#*E������s��L�&+����TbŰUG�d_�m���p�T��Pt���U��.b~�֝r>�@�	V����KL����
�28���>-"�x��_�Ho_xOёQ���E�62*|��a�Q�������D��_�?Y�o",�֟K����S�'��_D8fXȈP�a!��B<#C=��;i؟L�g������� ��`��p_3S��:�>�ɩk��	��YI���"dqD�&,�D�����8�~^�ίA`	4.��ƒXz�(�F�Ӽ���E�~�u�61lld��m��f���kgjl�bo:h 8��3	t����	p2���i=��f���`;ǡ֎ffN6&NN�7�9�eN}9��[R��d� ��O�b����?޵?m��+V]��fm0p���!�b`bcn<�d� �=|3/w�m����@"L�(|�[�]�̈́4�C ���L��!�!�28�H���94�MQ�lE!����S��m#����b!Q(���O"$�h��p�~h����/��3�$BX�2���r�:0b���g��9q���K�NZ�p��'37�Fͻ:j��)�e�X�,�^ڡ�)���~�-�E<�����.���:�pub��i��02:*��������k>>I����D��b�ջ���d����������#�x|�D(�.�I�l��b8��&A�H�S,�O��e�9�P#��-Tʃf���"�| "�o���� J�j�V�XY��Ӻ��83;75����)�>x+v����n��Am�����W��U]@�tEG�u�|�
��PPI%j���/���{	�Η��9[�a�_Im��>z*���W�'h�ү-���2z�:Ws5�z�=�����~Xt�ڍ��f>���%�nL\dӅgiHx$����ܓ��뽦�8��u�~*�=��|�����{&m8��zLB-)�E�z�o������P^�����E��@�
�)$�%gF�_U���}����@��#��;2j�����#�"�E#F�����[XZ��͔���2UX�)�]?y��ԉ�"���Ei�|\#���ݼ��_�xС�d'=�=&�}t���p�qQ�G�M<slج	Qs&��<&lL���w�\�c��.8y;�~�Ե�&VM=��'�$t&\��py B����=����E�,"�kn����o}.+;Å'�ۿ~��eA�V�>���C\��ma��`ol01�wބ�����F~F>�C=��\\L�ݬ��,�ݦ-X=lܢ�E�*$��̦Ȕ�|��Ks�]����u��o|�n��5�n[�����<40� �p�`�!�����"�pu�ܵ�в�'��->�(1�*��_�Ӌ��B4�E��3	4���Ƀa�1>��E�X����J($�T
�hmЫZ܉G���"�g?����@{@~:
Z��G�Eu��DoR#V �j����RcD�HTG�jhP-����s�z&DQ��i;Y�~.�w���/��?,Ȥ�Yt>���XB����o��`��{��JE�O�M�}����R�^�W�z���c���Mj���q�0Dx�14��C�B.�\>��������8B:WԄ%hl��U�i�N��@Ad�D�$a7N�q�͌3��r!��Qɜ�7ˉr B����l�W� �d�B����1��lq�+n]ΝkWn>�o�W1��XN^���� �����Uo�.�(����\������E��5Rq�D�ŗ�rdo�ʏ��?�_q�wD�Gp�t@�NxZ��%��8�{I8�t��T� ��w^D�~n� ������������1Z?ST�4�G^7���!�'�k�t~���A�R}�� n�F�{^�g��W�0��r�o9m�]P��+t �����'��K���"' ���F
���L���2L�� ��5 ����$�J�����I�O��~`$���n��G�;�N1:" ;�E�FHn*t��":�5a����3�F��px�G�����)��ڦ�����>�#B�̚[V�F�����L�P�&49���Ǘ5 0��2���_"���-�'5#���o"�]����7`���C���6���o_5��-�t�7pw
D��`�nop�3��޲�r�[�p��1�N�!#�������]�ᓄr�P��t<K+|]L.oА�X��<���2���`�!|[X����~��m`nj�����g.�K+I̩I+A��*��j4�
êA�Q:�؍��EQ8X:�B�1l�/B���z�ɘ�Y'|��w�n����9��ߊ%�[h�=|�N����"%^����N��D��c"�M��.鄧na*U,�Z��n	�n����������k�2,�E���A*W���*�ol�]�1����-d�L&��+����X���Q��ǩ�gm;iפ��cI\�[�����#�_Q�ګ�&�ܳcO��SYD�[�������_�p��s`t"���P?L�7X�D�V�z��i\�������I�P����يw9�≛.�p��:�և��%�^��>
�=����� GrI��''XI'���l��t|߮��(��ɨ���թ�GL[��U��]�1���"��E�����G(酷�V���{�J��-�S��־�Jzp�V:�ѵ~c�>�|����)��Z� {�=0(U��\�[�V�}������i���A�,S�����Z��	�?J{��:>�To�Q���S�7-U��RwJ�?h>��~�����3��}i;��N��� {_�� �:�
�������,5|�$ B_o?_ψ��a��,B/��q?�P?4�O��k�Ǭ=yNp�_������fNZ�`��0�y�Ɔ���=��S�1p�ǅt�>*�sL�׸(߉Q�� �;qT��[���۵-t��M*�t�	vu��)(��Sd�G䱸r�HEg	��/�j�����lA;��������|ێ�U��<^㴩!@<�6�v��C�I��[V̇���S��-�E�V�v@��>�㦭l"ʁk�
4��-Hέ���ЉK��5j�
1v��i�-m¬����+=�"����p�پc��U[&�Z�Q��S�V�ɭ!�#� h@��(VVT�4�uHb=�[O4��H� �b|`A4G,��ijm��*�~�A}q�gĒ��%�F^/M�������
�	�v��$0��ӎ��;����Jp�L)Ԁ��`7�I�HtU�	O~�D�^�d����>�Q�"s p�FI��b`���9"�2h<&��B�[Ŋ���	˯��I�WQ��־/hYQ%����x�{e��&Rzy��(S�V�,���)B��C! ��_~T6����>�_ X���{HY
E
�~t����+V	Zޝx��%���G�Bɸ�%�/K;>3e���� ~��"o#2d����K�V^�]�`Ϯm�w���x��W��'�.��:Y~=a̲��S�"�k�hm}��>�a�=B c�\+��YXP(��e����:�<a�g�
�pO��W����8�:G�����kyQ�q��aJ� d�_�ܖ���"���s��O�� �E`�)���oEm��Q��ǐ�ӥm�L0���A�����i�����'A�Q�[i�{��M����m@8��7_���U�!�:���7wϥ����ן������
BaDH p�ނ�UyCC�=��#�F�'ª��E�B.E�Z��v�
�������n۰r �!��k��Z�pz��˘p���#C�F�y����D8w,���>�&D޷!���G��4�"��x���{�V7`�܂�&EHgJ0x:�-�%�_��6&K܏^�$*�@���lQm������������/n�9�u�h?'Cwgg���&��E�&5��u>�}�m��|�M}�=���vr2"�q���'}{O�)�TE!��ͤb~ު��ݮjY����M��[/[نZ��68d��!�=�������.BoOO_����/]�m�U/^WU�x9���b\n��ޚ�VVQ;�r9�^C6��dq3]��5s$�<9��iⷡ%�&�GJ�\��=(5�k��o!�o�|%O�f
Z��N��+I�-���!�uT/�'��z�E��������J�?K��R����Ku�"�r�	&�� ���������Z.O������G�0_�5��@! Ġ)"���B�{��_V���⸤�W/�rS2�Q�����7����U�S�hn&�RXl=}/�I|z
8�OK�(�/���{�^XU��_��]�,6�Ť�����1���gѕ��ŅE��������E�D*��Gǽ��9$�_�4.�LgI���7o����:�̅��Yy��=�A�X�)��6�@̕�?����q�Z���E���C\H�"�\e���=P �M�BWt�W̛��������%:t����������˼'έݺ��;~�v��F��ы���-E�:L��*T�b��]��ni���#��Rv�.j�����o���xO���8��~#T�({��7u�D�F(��×t �	����g��$-� U�'I�[�0�x� ������r�o�p[z�/�����o��(�M��^��{��7��j����+Fξj��r|qJ)�nLz@�h?�pgG;{'o�@_�@� _?=~~ /�����ۣo4
o�D؈=N�Ӊ�ՠ�8O_0jX����q#�@(<<���������|��� 7� w��A^���#C|Fy���q��r��t����p���\�x���;}B}C<|C�J��)9�&�_>�K��ڿm?�0=��E���Dhkc?h�Ah�{����� /G}�%{��ζ@�f�M���������>vƮ��-���5���ᤜ\u�ūhf&�����_��14uQQ���bK��"9jD8D7Y�A`�!����������-�4n�Ҙ��bܶ#��:�`͉��s�x[�(o��61˛8��]�#��2x��w*���&^W1A3jɡ"J[A�pw��c�����-R�B Ԁ���ZM����r�5��*ZKF-Y���"��~���΂�EHH)|	�Ɵ�"
����4:(��!���}���/�����@�ܼ���fchT�����3r3/^� ����� �$�/&�iqeAuc�03/+�� .�e]TV���\�P��壗��3
��^$��7�sJ�_f��Aֿ�J�)�*�.�.�z����&?73��c���*)!13= NJKKs��22_7c1q�I�ΝǑ)&��+�  J����'��'�ܼ� |'��2�V Q��Vm��.b����6c˩�ŇϽ��e�����|M'!C�%+�dE{j!r��1w7�įH�?;)v����'�;oN{���#�έߺ��=~�V�1�^��%�6�U���/ �I���}��=�@�'�r�I�v��#�
�"J���Y�w,E_�-Tv�U�bEP�H�-�u���z��6 8ʔ�rU�Bۣ�v�Zt�� $�0�.��� �v x��~��-]��no ¶^�ַ���>�Z��Z�B�����~"h��tAW�C�n���Q����6��7���������������A_��������o`��@�u��a]3���w�f���d �ѣ��,�������KC;7� 7�p_W؅� ����D�����l��h��`��S����:��  ��'(���K��F�����f��"�o��ባ�݈ƚ[�h��d��124��x������ �An��q4�������������r��� �!vC��k-�C�a1�!�A*@
L�B��_�ƱDuxZ����b�����51725��/���:���h��Pp2 |{֖�n�NNns�-�=��	3�p'n&�N�����ŇN�̞��¶�)eHi-Z�4�|��Mude=U����#�E�k"�ʾ��Ya;l���S�����6u떳υ�V�@.jy�NM�lǕ�Y{�,9�`ϤUG�n:VM��n���Dl��'�m�76�x�o?�v�cPY�HD#����z�U�&�����߂��yYy�Ee9w^��/A��r_����qu<����C�6�$�A�՗��������j����W)��ཇw�
r��	1��T��>.�YEI1�y��������'Ϟ�54�,B:��`�(�f,C �����He >���w�X*�IDu��+$��f��y^�+��'�I�K���=!W�!Eh�kާ��n*�#� �ȯc^�m��dם̛)5{O^:y�-;J��/�D��~!����-B��aJ�¶"G�i?BV'M�A�	� ��C�������{	���G/B��F�-��X��HZ��v��]��Pj��T�0�6EK@���\kIO�գD��L�
P��Ot��l�Q�tiZ@ߨ�E�Q�ՠ�r!]���	�J���������r�ø�������&&f�ff&F&FCM� �F� ccS��0anayM��h�_�  �k���?D8r�_D�joagah:�>\���!��}X�7`���0?�Q>�}<Fx{�rw56r6�d:��|`D�������`�π���z�O�H�EHap��W���߉���l^
cimD����`mkgn�lccgnjebd8�`��������9��62p��b1�\���r ,B��NNFv��֮����v�!>!�sK�5MҊFQFVZϜ�r��㗫Pd"WNb�jь�ۏ[�X�y�XX�Y�[ۛ[�ZX51hnfdf2����kkm����h�<c�i�WD���,��£����O��y�Y�n;��t�o'�Y��ъ���;���,o��4qC��#ز&nk#����*�ݥ��~)�7��"v��B�Z����� �i3��<mG%�C%�%�BVA�[�|��ی�/�ih�O��"d
U����������#�Vpy�/_� �Մ����~w���&4^$Sr%� RʉL�P. ��򂂊���, ���$��+7��!*�*+kK��f�r��,,-��(tt��t �W������gd&���<�U�F(�*�u�ZfF
�Jx�Lġ�X�g���VV4�T?{�و ���nܨ����(TjTO� �p$G Ѷw#�S_gg���!���r�Z�Tj�|�~3%#�u��C��l?;w��#���J	���S��%�V EҚS�_�v�OZ������x�2q߽�㱅G�8}�����7o.����l3��+J��y��t��Uӷ�6uޮ3�v_�EK}P����q�ĮR��S�#V��z?B؉���2�]|<*�����"�+[�vXWm��R���E�{�a��X�E��!�n������ Dx-�5�izZZ�lhdd�_�4P���� �����!Q#� V�7W�6W�5W�c�p�]�$W7q��(�r�9n̄Q?�X\���m��M��� `A/�(WCC����Z��z[G�39�+���7(3��	���ĺ���E�����o���_�~��jL���).���P_���`#��^�@��v�N��Nv���ֶf&�C����.v�@���a��:t�6v�1
��v�v6`5��� ������a��B�B&�`k�YHJ-�H�*=y���{�/90����֏���������������������������^P��4u��qwrq�u�5c�N��%Ul=��yؒ�9{<F�>����	��1���R)������H�6�ōT�.D0�,)��i�t���F.>L��ȝ�Ґ��Эʴ�'X��%pN+���o��p����z��:�[��=V܍�)<��/�C7O�cW6�_'��;��'���,!����p�e���U�"2�*S�A`��	�|�����O��Y���"���9��_�P��"���̢b��߀����&�((0��������u���WO�W�64V��e j�={��߈�MMK��~���޾{153���3��Irʋ��i��ڄ�������KϾJ|QU����Iqnzav��7+
�k+��_&ggf���D�>Oy��[T|��m��%��#�$d��f0��8^�т~~~a1���hZ��7o���zzJ�=fS��Ǐ��q�VtBn�&Rt����X�v�����$J\SY�cVC
����`���+<I}Q���8�ڕK+�/+(�\}�<�=Ԥ~ߤ�E�;P���Z��{I�p>@;og\IEI� '��/^J��3>O�u�J��I!�CV���{�2���"ɺa)����V�X���;d�v��C�풷����^Yg��筴��[h;�"���;��{�K�<u��G�T�A4������D�η@�]�!�����⫻ŭo��lI;���ޮ7D
����ӂ8X+zw?;j��K1�_��ߏI��eai�'5h��6���u1&�������YY���EW�a��6�k��휧�F�7~���`���#"m͇��mL���������������������6��#�������������bPh�sP�s@��o�Ϩ	S3�*�Q��j�*&���W���_D����"d�x��_ x�;�9�]�`mmebb2`����f@� '{s;�� B�-��{��.fV.6�.V�~~�3�u��fr�X�&�`h���C'-\rx������~������gm�`�j��������j�����`�ho���r��sstr�s�=s��9+#��{�\y�Iar%��ֻ�\�G�P�%��/�vg��Ե{o�!��A�7���TA���5�U���B��y�"��G�ܱ����A���$�*2����"H��|Ge�_��o�6{׵ˉet�pM!s��������u�XB"��*�'���nj��#���|5�X
��Қ���/y"q[w�Z�&Sh���Y�y��n\��UK� �ZW������+�.e�U�&�<�.Hi@�]�v"+;���0=#PYU|��͘珪�K�����5��LL~ZR��2%PR���2.%5����y̓Ą��¼S��x��$/#>�AvZ"����i�%9�qѯ�ss��=|��*9#'�� �
ȯK .�oB5!1h,�H�rx|p,*)��+�5�b�C7H܊�[�ڤܘkiIq�n<Nȩ���b��.@A�t�[�	*	�M@�gb^��=w���Kz�������oߺuk���h���6��A�wU_���Y�y�YʉYH�'��?���GU��'2;�w:�}�B�5���͗}�n��
����e��<i_��?)�߉P$o+:��.��x����:S+Q/�_V� DUo6�^�V���hI糼z��W�	��@O�k��Lp$(�ВnF��b��iN=A��e7q+��;)wS+g���M%NЂ��� ��A6� >�L'F�:u>:;&��ʽX���YZ9 끦�%?@��$��"1b�^��UM05(؅�P���%6������M?r��ـ)��{9t%�]��\���"�QA>��h��nt�K74�5�����������\g���]B��B6�؟]�P���<�Ory��z��_56�K��Uc�����ήkD�h��p�z�:r�B��p�oFF&:�up�m-�L� ����ں9��ۍڙ;ۚ�ښ�mM]�����"�!f.���)�yE��Zz5�Y��W5�*)��HW5�h��eF�������������_������+�������n�Q;'��������,\5v~��%�.��U����Z���Ǫ����a3��M���e5����Md>�*@���D(n�(�3�8�!��q�W�)v��?�ɡL\z�N�XB.[Nek���kN��u�q솙�-��������[~N��y"��~���ӣ�iOj�L%ն��l��E��~�C�2�H`J`6�������j��� g�Sl\������Neru�.BE���c�H��o�9x|aIE��c_< "�v�Dt�����g����׮���jaA��'��b���:��&;;���;ϟ���z�<�Q���E9��|��nV��C{����:��Û���'�^:s���ԓw�G?�x�v����Č̬�/7��M,���SYX2E�6aI@HuH�BX�:�Aj���0;�������8�1���;fg�}}혗wN_�q�En�#i���v���`[+�CJUq��ښԗ�O�\�tq������O&�.��&�f��]�qMe�<r��D�Ф.|s�Ya��Cs�큒0_'�zy�w��ڍQG���. ڡ�	�G�d2;��= r��|Y?�ɢ�"k 
�eO��^n�yW@��]sb���y��-=�7�����wR(��LF�ϢG��E_V�fy�7�,d���o(��~��=��P����'�)�N�v�����f����Gb��5'l��=��k��5t���d���
n=}u��M�C�[Z��E������#��kju�j�9�F/�)3������<"2d�	�Q�Az�<}�|��,���΀`7� W'@������������^�a������~~�!��U0��z:�*%·	yT&�g�?��Kb�/�W��"���"��!�	�CT�¥k#G�������3747ddgf�lm�lc�hm�hm�lޗ���	,�d1���0�������?��� Kc3GKSG�!�f6�q�UYy��
ze#�ūǰ��(y�����jTe#�ڝ��!6�@uN�~A��"��_����m�U��6~^j!r�;���g�;9{�էy5HNF4w�Š�[�&��� D�EPy@�M,!�-i�(��-EX�����O��%�K�⺡��a��2�[���)���g�<��w
���Vh�S�����_��*B9\�O,�ʤ��#�����:�K� ��8���ªʔ��W���H$��y�e���2����7�5�JP�L��/�ӋP��JdR�>����q�⩢���ܔ���޾{��S7n��|����=@�����~�lVf�W�<����v�����/��>�� 5%��[O���L�q���W_%��ز�ֵYI��yr��8���ӻ�;��=y�(--ab2�ًW��x ��w�MX
�[m����، Y�D�(,�x��U<y�抚�'��%]rsǂ��Kw����P�j����le��	�oP}��n����T�5�� M~UQCl��"2�!<W�p4xcd!�5�>��B�	��Dh�=��:z�al7D�M�{��pw�#��]/��:��^x>�Z	�.>������N��.�|��u|� ���)`A`k�����ak�h��-^"y�6�j�B��P6�_q"��2����Nh�����\�.UC���|E8�B��uxѵ�ƷP�
�p�~�q�(��9�G�8�hrcT��R���/�C�v�����)�A,{����u�ã��\��y�lp����H3+�?3K3scӡ�&p&���E��0l؈�ܢ�Du5�7V!�;O���033r�����>�~h��ފ�l���`��0��1��j�@롃 6F�팇:�����Z�Dh�5,<0((( 8�aLFA�#)k`��R]D�������'�u&\��o��s&�6����;z�ܪ՛--��x���Y[Y[�� �[X8Y�;Y�:YL��\&��L��{m;���]��Ghff`b5h���+k��vV�!�/�s
��UL�8�C�YM8z�
h���s�=}�l���l<<�������pw�y{z��0y,]�v�M#'�NʪȮ�ĤW�8y'.��u9�ũ��s�Y�Ռ�f.�,AS�(
���mf��,�-�r������4r�˴��V;�<d1f���5���292W��+H�V����mW�l�\.�r�l�6z�!����"��<������
���
�*���2� �O[�L��D@�B�si"A-�(�ź�;��?w���䤂�ʴ�ͻ��H4UKG-�Z
×)�^#W�P_V[ۀF�4������r:��s�,��JǞ;{�BAө�S'��T<����U%b����M����m$"�ϣ/��D�v��	���Eu��͒�\w�����2�Ԟݛjk�����+#�oz�.]>W\\��N�9]Y[<}��M"�S��~z$����3
<��L�)����'żH�)����ąkh*�Ѕ�E5ȴ�W�����{�����؂z�\�5KՍn�V�
�vAU-p�v����,�
WM�6	(i;Z�N�2��F8AK����V+�P�yW�O�ȝ�ٗա�/;��jQ���B�hO"�)�=���j���Wg�S�lgu�NW��߀xN�����n�98�뇫�`k�-]Ԗ^R��W͢1��>�~�����gP��Ǽ�h�Œ$�g���K���]��l�p��4�U�sE��2բ�%N.4����oTk��wL>��W�	!��Q�n?�UN��$�Y,�F�{�&�}8��f��#w��iǉ� x�QCc��C��>O/W{[kKs{+k[K+[K�a��ss
��kk�kj�a����O��h�|Pj�pƆ��5p�6vw�����`�hc
��W#�"�\X�1lk:�������m[�hi }n���#[�|����ӪP�
�E��2�Og	8Y]#����_�y����EbDMSӿ��@�6�(@���]�{/:"r����s���������������	|��t���{c�@؂ C؅ {�!��C���4<�������k�����B|q���ۈ6�M8������B'7O;gg#SCkSG'k�@��㠛������rՆ�7��4�����Li#�U^MR^Cn�� �CqZq����,lű$��(�|�t�-%pdX�����]N�Q��U�xP��R�X#+j��r�MMv
z!j7���_!��TP��NfcK��]�:�D�sa��PG!cJ�Mdb����6� �EzZAe����4W2����<���PR��&�
�Ԁf��be�f�}*Q��oپ	�T��Ү]9�� ��v\�t��G���ܻg���h9s�8U���r��^����]Ǒû��Z����/�p�X����nظ�	Y�ݥ�s�]/�rٍ'6�}:v�����<x��P*���eͦ�L��+U��7� q�x: Eb3�*�\���}�C ��ӳ��*E��w��|_R����/KNG�<�n�/E�5�<�
���~�P��#�6�������'���M?p�ѱ�����w�`��;{��=v+���W[�>�v!�TtiZ����RH�;����ݒ��&� d�D�|�ZS��꺠-���T%�&�
1����z�*��V�R�U Za��D�'��.�FK���������6�����S���ܛ���~�{y'O1b�|��H��G��e��ЙT��S9���(U�8�����Rm4�DF&JgCӎ��l���@�h����+�Q�K/���d�Δӹ�
��f�?z����-{���������2wvs��� z�vV@�V���f�fV _o���a9�U�u�h�:��"����<ǯ��t������ `;`A_woW; ?{K#K�������#�N^.�ޮ6>���v����>�6��&N�� 5�<aZ@�H ��2jE��
%i"���W�����')=�����d�h�����R �݈"<r��s'O]��2���403�27��0�	v��@�Ζ��f��f�N�CA8 ��8��e�̍���,Z��
>9jĜ�\TN���Z��n���I��::l`h4���6�.vNV��2Ύ�Nv����a����v��:/)�0�Q�D�DPKȅu�r�
é!�hV%�UO�6�(��a9R<WF�ɱ|mZ%s��,�i{gy.�W)�� Cu�p�PCu5z=�	Yz`��3	(զk�F.ٍ��!�T�6�΂�E�/R����E���  Z�J	����<�:�L��<(ʒ�t'"���T�Uj���a�Jj2��<}B�rDJ%��%2l�������✲�W�Y���=���ᓸ8�t͂�+W$�$UTW�]0��훥e��7�}��.��z��5��p���qϟ��T�_���[ �]��Eܓ���Y3'�G��S�=yPQV�b�⇏�����ܵ��!��d��c{i��Ջ��!W�'N����f4zˎ��N�ሤ�&L=t�����v<Bޝg	/�r�=K �%]�A�7��S�ܪ����⼒J𔺳�ԕ;$��C�K�g�^I*��Tr'��E��7���^����V��7�=k>_�9��p�y����s7��z�����.�:r�މ�g�&�}�Jܹǹ��fx/��A���������7}���z��:Հ�U�o�m����z$5b��kN�j�^�6���U�ªSvr�ݺc?:�Ѵ��m̖�B��#'�Zp��1;!J'D�p߮�agm�����3t�%mº�K���{����5��o������Q��_r>��q���M�P*���O�! �*1�5}A��#DP� ��Y	�U�����'5'o��<t-<r<������khD���� â�"�BFDD��>*j$���72,2;+����_EX�L)�N����{îC���M��|\�}�|��\l�<A.���ׇ����7*2@OT�g�����9\���:�������#�µ�y��fq5F���_E�����K����/�W�gƽLj��"�3�:2@� "�n$�x����O98�8����������-�L-L�ڙ��EB����N�����.�E�l:��d��� ;��vC��-���f�[6m֪�
Rq���Q���w�@��&,�#�g�����8x� #����v��6��b�&�����VV����^�6m]�y��)��r�2�j���+0e�`����]��EX�f��5n#U��5�D�Ǘ�
x*��SB��V�`׋�a[/;?��+�y ���2���(�cv��z�5A��q����\H�$]$�_DN�fA@����E�{JW���MM� ��-S�'�t�2�Lɖ�q,�΢
Ē�6����s∬����R���M8��e�v>�~�ūVM�={�ر��O�9o΢eK�F��5��m�C'O�x��)_`���z͜>y׎-A>�'�۶u���'N9{֔�`�� ��S'�����k\��"C�/]12r��	~�^���K����u6<x����F#�F��m������c�/�>,�/8d���^����!��y��L�bӮ�'/��mue#N��Eb��_�6�c��U����3�J�A��t��ȸq��&"����$P�H*>�,{ϝW'����:���r�����a�?inǿ�*�bӯ�y|����;��ٳ����{��y�\za��ջ�����"u�J���~7t�A���jP��Zm��꧵�-JS�o:�Xt�㌽�N�A1m�ۂ�C�W���h�j-[���΅-Lm��m-]:eF �P#�+�b�@)��%g��R�P&�m���O�ؒOЙ��7򊘟"��>�F,<|-���ff�z�ю�ty����&�[{�2v+t��˳���D�\w�V=�j^x�bL�Ň�{�ތ6�0 ((0�?8���	
�9<|�g��4��b�j�����fJNx:�>bɡ���O�0���&��%2�'*�wX�������,�3�����V,3,���ǎ72d��P�����DL9~T�(���o����@X��4����p�q^%�
ͫ��{���?7]=��|���An  �L=D��@�uh���������p���eD����YP����������~�����
���fi���l2x������n��!n6C]�]\̜ܬ������4���rY%���o�4b8h&M4a`����\��p�@�C�̌LL�/:��x������n�D��uqvIcz~]~X�ũh�V�xUXa�_��U�5$A=M�Ĕ"�4O��å$��VxQ9:�O���P��x����K1p%[��.j'��Ȫ?��;�����z��w��V�$��!B���E��r�}���~�@J��5~��V���g��zY�LY[փ�I��V����	��!�%M&���+[I\��EyD.S_M��\��AS(K֮a����&�7y
`¤I�i3�Ϛ;gμـy�� @��?XrƜ����s x0w̼���̝1{��Y���=sƟ̙�Ϭ�Sf͞�9k��ٓ�͜8y�D��M;z�董G9*r����غ�L������ŵ腫��ԡ�\1����-������.�á�y��7����]P�ĉ�Ly�.�����r/Oե�+ �[��������^S�bK	G�>Z�z}Uq��#{�<lf��\8m���T�?rn���oƝ��t��������T¹��z!���׭�A��TYN�2a��U�rc�����X}As���Ct�����V��.B��[w���"�� ��lu��q�y���iu��!�ĝЭ��<��+��r~Z���
���6S��F����.����)�����^vSr�� �&��/H�29}%��^ Qz�'%�����5<��z�P�a`HpP�_p�oX�_dTpDXPXpPDHpX`p� @/������j$��UY��������%J�C�[�n���#�B�#���� BA�ss�vu8�o����N�r��-���A�@�����&����N��]Oڤ�p�|>1<����r䤉�5��xV��D��i| B[������_��*������,�Ǳ�("Q/���4Z-��g�`��fw��颢�ׯ�F����ieg9��r���!<Y��������lS�� ��L�b1���������j��a������1y��)3��U��,@=
�hD� 4�&7cHi�9��.��z�3�p ��!���!�L-̭mm]��aBjȂYEȼ
BI#�
-�D� ��E5A\G�#�f��עy4O��*�\m=�{����y/�4�Xґ��b[�%�p$
 B�����1s��4$o��g3�ݺ����o�ʁ�@{4���Ɠ�
O����Q���R�PJ�	b-A�Nv�o��Od�7��K?3���M�C�q}m}�P��	�T�ݲ�����r�$�~Rylpԋp㮝�Ç��z��[pԸ��G�������Q0QQ ��v���UO8�����)��a�A�a������������D"��"�G�FD��OP�������W�Ȑ������h*MapDRx�������,�w�9O��ǒ��X_��]���q+�o�.:WD�^�@D�=��ԳRR�%�wܽy}e��ۗO��]<����	�>����NK>�o���>KH�ix_����#w]���߀R��ŜoY��wY��%bh�ḕW���lj��D_&l8�{Q5o�v��O�ԝ��I�::��7|�;*�[��&m���oz$-�X<�W����>����s{5o!��YC�R|�� ��c��ץ+�������oY-��ĭo%�n����o�q������ГBnԼ#7ck�_��$�GN"�����w�	��J��ÂC`|��"B#�_�UW4TW6*��+����p�^�S�B���\�',����i�
�.d��;4襟Y
X8gR?�V.�sڱq�Z��В����C#��O�_[]G�6��Md6��%3��D�����������W�и�D� Cs�@׸��m-Ts�)FC�{��:Y"t�6v�6u��p��t���p�ˌ�a��M��b>��b(P���WW+'7'wG'7נ�a�FN..E�4Pk���:$���ր� �U������N�6�v�
�P�3�013"t��^�y��-{&L]�C���
R�[�� �10eXQ^RI��NqE^OW���u4YM��)
�R�����l\u�(ՙF�d�A��R��҄�;�m��-�W��f�CS�O[���*Ћ�ʑ��2*WN~����(���r�D�,hE
�9��Y_�T�>�S�����6����Hdj�D1��'r�Li;<�*��Z4\���q`���u�|K��RHK׮�t�3�����6z�ȱ�
���� �� _ ����{�y����z �	�<��? �������������y��O��/\������������<���
��u��s��z�C�a� X�a���Q��F���:������y��M�H"���E��RYL�A(�Hd@��N$�)�vp�o��/� B�G��ϒ��lyC����H�����Vn�w���[
c��X1i�0畣\�M���pvߪħ��l����U�/Ӳ��%d��H�I%�	+/к!�F�n����/%�@ �;��?�q�GE�O��;|���_�:� �"T������׏@��;E�IK���}�;|�u�T�'U���?����A��or�׎����y��7����.l���A-�������K�G"?��OF��Y�����_z�~�J�J�V�ҧ�����wC�����ގ��}U�XD������������{������.°ఌ��ʆ�
 ����O�@��$��d�EԢ�Q��&B��1Ã|�gO����͍'��,��F���`m�f�4LS��a�ϝ��a1.,����LB�2G�o���,�������<׋P�!W�hD�|��{}�����%�7g�@�^���Vp"���Ώo^�N~��`�`6��|���`KX�.�6�n�\��F��7R���&:��w6�ȣ	Mh|��L'G{�����@����	!�/^���E�i%y���E��
J	�_�����2�P��7�s�/��F2�ќB��(*%J�9=M�?ʥО؆��R#V����ġk�r5S���(�X��JJ+V�Q���4���Iz��N[DHf��l	�+%s�#��d�L��E(mku�r{��\p>r����9H���΄O^�~�5���L7c����Dg�2GI�KX2	UĦ�������R��"�uq�
�
��[$H���a���H@�0]	1,��PB��<" �`԰0�>��_80Z0xq0|� �N�a� �@y� �'�����@."���		����`f�:���`�a���2��+1y,
�Jf��Z�Bx��P�[a7���JA��-?��@o\�{V��;(p��+���-4"����w��?f���%���O�q���;�Nnܲ�Љ-��En��|�$��'�� �N*���Qk.�^w���G6�S���7\������,d��I�.�Ė�TM]��д� �ۙ�P�o�a���j�NН���=Be�n�� �v�Z> �lpɺeڷ ���%�`H`h��=���������������+HZ;�m�ֶ���v��]��K�����uC/�H�����4.�..�$4�P���n�d��i��������������������� !���iY�U����U��*.�K��}�4$pV��@��A �"}s�O
��
X�d����  ��	�s���|\]��]�"��O�:�?.���1>^����KɄf:���K���јln?�b�T�~G+x��a-5��������lϞu+��Z0{����� 6}%&{K#kc+SGks�֣n��6��V /'k� +Ӂ�f]���\\]��|}���*��@��$��w"P��"�s�E8`�`��~��Ik{;���^2j���sR
�m=i�<�{��Y��LX�����\0fUtVs.B����1�+�����%�#l��&h��%�$��?\/��9��q�f�ik6���Ri����g���U������s�E���W�Oݶ������/$��'�8j� !�#ѣ!� :pa?:)���P�aW�%d��RT#��<E.?]B:p7�������If����P����136
ԟ��>p�$��x&�ƣ�D,2�,k��$
�@��&N�������U�S�΀�z���C���F��<�'$$�����������󑣢@���������D����`b�d`d�y��z4�+U�c��6�Z�WJi\6�E�rT��������|�V�m�'g�;��T��Į੻�x|�f���R��3��Zr`���Q^��q_��oZ�`ɔq���8~쨉�#'��2�k��q�Wn<y��ä�B��Ge��,V+$~m<��b<b����X|D~�,���m�B�n�	5�B�c�x#����w��wLMA���4y;[���t��O"���Q�.Q�J�m
M�\�!W� �՚����S��P�D��M �|"��E��*4�
8jUu�FѦ�u��Jy�R���*�c��"�Oo�UD���damlf5������������V_���.������Dؿ�Zy-
���� DXI�5i���p ¨ ?@d�o�������Ё&����Y�G�|=A^n?p���tp? MF��G����U興��FMc"	�s"��T&���sA���.�~��u�%����,��q/�"đ`��!��bW5 ������[Y��lk�c���VF�f&C�,��-M�al��M6��V�C,MZ /674�j ��5�C�N:���������Ժ&j��	��?����f��?�'�:��9yzO�=?l�Ā�/�Kp�x�In~��!�t�����S�����5k�Y��E�>y�Z\��/�uqձ��v�i1fڶ�S��j����̃杊_s3���,���b��,e+Y�0�����Ç�u\i^2�*oמ};�=Xt1�R�� ��~�:�w"��E"_A��7���*�I{�ޮ^z&/t�����_�F���E���>U�m���h*h�ɸcW���v�;%��x�� R�<WRSZ�������\RYZ��[�r�^�>��z�'��^��Q����?�0(�߉0D�����~�7��������������E>j�T`A��՛wV64`ȅUuye�%%�eeŵU5�O沨<6p!���-Srj�������|�ϥ�g�s�x����'^�R/���A	^���	���2R�c�3��1�����~}�yޱ��kY��zv)������0��E�@����9�)�w�(l��ٔ'U�g�w�/���^�AG�kF��T���UA�v��Q䟩�wt�[��I؎�k��� B�a`v ��TZ��M��"�7�V� $*`�|��N~��0-?���C	Dخ�u(�mJ�VD�MⷃD�PH"�]��ј�R>������l�`#��������V� + a@@Hj
��E��A�aAt.i6�G>:<ltD�/'�a��8��w��+�(��Dxܫ���)-oA�Y�?�,�K���_���'�E<�F'RX"G��P� "�Y�D�Ehl8������l��)�hkfbebdcjN�m�#�f@��V& k#+3C���ƃ���e�5pr�rp�qp�wprԉ0T/B86��)��$]1O�n3-�M�xm�z��֦fV&��&�F�&�F�C�����8���z��[�2j�t;��k���{�%Ϫ��!fV	��E��eL^z|��3[��U3z�lJo,;t�zj�*e�?.�M�z�Q��a!����J�z-���G��i��te�߽i���t̲m�ľ,��*�Ij��ݵk׎�w]J"ld��B�%��il�������n�����ǫB[q���-���"��xߠzy߃�F��+e7�%O��[��*����#Ĕt�Y|���(\"��O�K+�*|����}p��/S���\�]�`�F,���n�p֧����7��� ��l����lڞ�_�[\��Y�[w��rK��"�
! E! r��\�W��JX��ިL��W~��@L��-_���ė�a�@�o�y�6�8n����[��Ͽ:~_�ĝ9N�j5e����>K�Fm<?i��Y�M�ysҦ���W5ҥ��T0>R;����Φ`1��Ec����}P��ң�^�O!����*���A�_'�#i���l�{����������!
u���_7|T���- �X����%�?C!\�I�j-\��E��Y�S�yG�	�@/���S��ٜ�Z����� C��C��2 t@�b "$%�WVaU-Z��I�AQʰ�K�~N;z�ؑz�;�GC�~Z���Ã#�C#C�r��Q$�t���k�(.�+��k������_"����~a\|"��"����E�Å(��	,BS#cgWGk���ٚ�Y�,BK����������������������h���@x4`ogagoeookk����VPX������'�t��6�t;,c�1��3l�-l-�E�����������M-��[S+��X1v���Ϩ�+��R�V���c�3+p���k��{X>i����X����&Շ�ٝ� \}�iR�KT�Z
�-!w"�'!%w^3�*b�	߹�6]|� ,�j��[q��{�Ǥ��:�d���'�=��˲����>w��ԋ���$B,��1 ��[�l	��g(��X\)�����[q��r��y�*<<������Եj���y4
\}�x
b��ב��T��UIi�O^;�,�B�Rq4>PZWTZ]�s�܉��؂���llA�������z�"C��~DT� �� l���'���0�����r׋^���� xW�s�	.`h6o�Ǳ/�.[�m﮳W.%�&բ�L
a=�$B�BΓ�`*� �$*�@����@�t�[�]��#�,k��]�˜��i�Ķ��x�J�,�q�a�髯��L��>I��4<yu�1 }����ǟ?���z�b|GД�㖝s�.j��u�zV��f���������c�Y]�a�X�pÓѳ������L���3�o�[��/���E����v��?e>�@�N�z
U-����Qu�4]A�!n��G�/O�i�i��y�o(�V]Zt�JteZ!15�>"jR@`���\~p���w�)@_�	X��; !)M/���
��n&���3�f��'�\8*"b����Nԣ���P�!lM��\�]���7����-,��-�CÃ��������Ga#qd,��������v\|2!����p�	 D�������mci������j:x0�������1!�-͜쬝m]] �g��.� `D с � �X��Z���Z�x�����_P^߀�����a��S׈�G` H�˴tk{;s+g������3Ȕp�DG;k;k�]�Z�;8�{8zx�\�4t�$+�������XX��א���W]9���X�ƣ	u�O��T8�X�4rU�e���{�d�!�A�y�͗�N>�������GyIhe�7��������$EIڊft��u�ib�-�69>r�ȍk�ؿa��M5$�^��9!��m��14@oDKЋ���N�L��ɒ2�rGKb� )j���Z(�5�h�N�]f0���U���s��h�=�߮x�>�dխ���=���DB3E��\Rymѫ�	/^>�sh���{�%�+�,?.����	�ς?�g�D����a�N��:~2�_<F
D����k����}B��@� ����aC�,�M��"�Ufn����w>x��ɫ����	M���>+��b�P� .��v�r9M*gj��)�]�3�!V'�~���_��Rn!���Oj�P�G(3�}'%���{��9}��9W�Z�z��5�v\�r���V�|r����	Ĥl��JȡELۓ�Ԟ�����aS;���Z.�ʸP���s.�̿��\eЬkk��N[�P�2lΙ�j5[MZt ����D�j;�x�_�
���3�V����$<w�B���(P o筅O��m0�@ɇy���t~���������}��4y;x~`�حߨ-P��u�F7�Zs�aIz151�
��? ����C���	k?����������������
�aU=��W�$�4sn��&G��4,$dlT����$2�?������������������Q/Bp�,�@/wG;W;g�~�
����`y^IuU=Z�������������_"��~��F�4:�'/[�d.O7O�m,,͆1<D'BS�B�kfm��` .ԕC���BG[[++3Cs�A@��headmij7+�Ǔ�Uz�5��55h����:��M���4K;[3kKW/7OW lD7g�l����	.La��Dh��6mޢ�qӼ��>L(�d��g�L[|&l�ΩK��K�N\|Ň2U+�F��S�����Ӑ��v�x��ܳ�]�D�s��-?T�G���eb�P�s����Ik_���ڽeߵ�G��?�w���g�>�o��\x�Յ|f-^ۇ�� @� ��L����z`2�l���T�*M��*i��[�>�Z{�r��s���?7Xt�n�#���.�c�&�
K�$SA2��Xӈ�5�	�-�%�<)�y�YWn]z��!�� �����Bo?￉X�'t�M?߇�Ah<"��^�AAz��p!����!���!�M-'L��Ɠ��QO�=;w���R�_�#�\C����
�J
D(P�jp!C&#�%LmG�6n��z�{�b�A�?����DiؒK�W������>�~>�ٵ�'���r�����&{Ν�{�ԉ��v�;~j����	/�ϓ�(&�p��
�j ��{w?�X{%k��K�t��{���WR���8as/�i�EВ�/�dJ
Н�Mʵ{oq�_�ڏ|m/� O��S�|߆T��RiLp�_b���{x��ҟ-�/B`A�L×���p	�bؠ�7�|�rN�>��E�#�C'M�td���37�ldP՟��HQ���޷�am�J���}ו��/n>L�������y����e�uz�U7���
A,B���SL�m�����'��d�, 8	zE��>���������v�������?������W��r��W�Ѐ�a��A�ag.\-�E��4!�d������,����$�i0*�̄�0Q�  B<�r�ĩ�����0g;'�AF�C��Ml�� ڙ��[X�[Y:ڃ�Kks 8���
ԏ��Dha2�S������������������/3

+*k���� �Q��]���tG�@uE�<@� N��ۈ)�3���ܟ��Ȳ�7��N~��M/o?�XGW�mI�o<[��9��h��f^zYy�u�-T�}DX��#�B�	��1᳗a�Z�PD�f�����5�O_���{����'�ܵ�E_t!U/B
O��N��s��~!�#���L����R�]Hc+ٲq�����S�.%e��I�.Cd4ST=)��z�)������-���O��L"��DHa��kP�������ݹ=.�i԰0+k3;{+__o��ɢ��E��������)3:��ut��N�z�#��ED��M�<uμ�6lX�l���K<����T�\C�B:��ȯ,��*a��Pɒ�(B!O�Z�&�O[�t1�_y]P\��I�-.>>i��*Eۙ�K�?xe{zv�e5i�����cGz���:���Ӈ�<�fA5�ab�{�_ϻ_�~(�u=�,8�����ԝ/��Y�2(�ܹ�zR�Z�"T��%Ws>ְ�N>ȼ�,G�b��qQ�[y|w����R�2UZ�����k���^��-[��U�����_!� ����R|>�7mǹ"vg��땔�+R:�-�ng�i�!�y�Pr�vr���ˏ�N]�"�����W̋�����gV6
�XOJ����\��u#��c�� p��`������������������O�~�X9�Z�s�-L�-M�u�nO?	��߸�!�UH$�!��D�kh�W�K�w"�o��MHH�Ǐ�>r��҅��-�q4��j��9
��l,�m��,,M�̌,�֖� ������� ��@�F�C���``0����ylRZf^yU���� �XU�T]���C4��ǃ����(P�Bw7X�..����������$B{W�E���Y�v����5����,dR.��\�(�'wT����b��Az#��-�`��UT��m5�%��OT"�Ji���]�?+�YZ��)$j�m8r�NV��	Z�mk�_~]H����]{}C��"|�.��k�,[��|l|=]Nb˚�\��"�g��� ��;D�s��ņE��`�X�o�H-)���q#�42�����߃�&�HK:y�ry=��7���K{��v�P��Qq4�>�����&<"<�dBb����mZu"��:��3߷��G������"�o���u��w����������(]����� ��AA�q�i3�)�&�f���fߺ}�ԩc��"37���&�,Bfq6_)�+� �R`J����V�7�۰���I��;�"�@Eh�b+'�9�{��p£��l8��uu죄3Aa�a�Na�!�>Aa~��:s���G�3J����/J�N�j?��'��D��#�
��/��w):�؝��R��:J����bD�5e�������.�ԥ�e[�&/�u�E!��h�N��y-Z���ɮLe]�CU�R5�Ț4�G S������x�P����!B�z�N��|�Q7v!��C��M	�o�͔Y��	!��;���ۂ7���T����f��o7S��Պ^�9�>������ᣦF��"D�%�>+��L�0z܌��*6 �����1<����~E����"��G��e����8��Y<k����7�>4�GQ&p�/�j�scp��<�E����PD*���C�rQh
��ܹc���/��9DW}���`cdcjjibbf2��x�	���5&m͇�Y�����`3�?؅��-`��F��k��\A/2%#�?D� 4 �w>1��4�u��wqr��p�����t��p�p����rq�qp"t��^�eǊ�[��Y����_��[�_�+n`52K��5xqVX��Ց�u)�ϯ�+k��:FK����Y���ʾ>�Fm���:z�u��ѿ�q.N��[�1��O�����o��6�u��u��
�{�Tjn͎ӏ�� (C�!�(��{�'��!R�K�S�n}=��Qw�΅l�~�=C$Y!1'�ؕ�OS�LX�Z�~z�Q�+oe���_�,�	*���"��Y�)M�Oo\�v��4[�"KKO�G �~���"��"�!� ��*�t��+$A�:88�τ�Fՙ484 (4 `xx���Pc�i'J����䉃��^�d�7W�X��bR�3X>O.p2]Q*�����TfWՍ���*�n{��B�h��g��v\+4c�q�T�\]�^Wq?)�+��.�	��0I�&L�4�����n��l���k;.޾�Zs�y.��3��z��~���\s-Y #K����\>�9�e��k�����:y�E�n�\s�y�U���ƌ_r����~k��UÅ�Tv��5����,�r}�i��Rr�@I���'�.�~��� P����]@��Â- �y.������b%R����]Μ��v��w�;�����Q.�����i;���X�::�].��]|���݂�g�;+0(r� �n��������<�cgg�hgociedd2p�``A
�>����e�py�a1�����>v��em�tELa�LMlL�ڙ��Zz9�����+.y;[��Z�	�s�
��
���h9�����b(��������W,�sw�r�FJz^zv)���Y�,���{�~�������E���t�2�'�j�$��=Ǯ\�����Ic'[Z"42��XY�452 �41�2hc6v��;���F�C,��Q���15����F���I�)�������M(@3�p��C�M-�@(���urs"��� �����9�� �{�oݹo��Sf��"9'��63���]�@.n$�5Q+P�*���m��0�A�6���Akid�7�;����G�����z]'ldu`y�8����8|%)��Љ�7�'fԖ�a�]~��ͻ�_:u'�U�,B�D�	\	p!ȅ��z���U�t���2Lp&U RNkq"&5��W���C�mZXf��_�s��$.O�n�/vJp5Tqerxi9�	D����Q�������7�ݸs���#F�[ۘ��;��������������~�_?���2�k�c�N�Aa�Aa:��'.[0oώ�;�nطw{�˘�����2 B*�B�sK�jW&�ʤl��%�玪�{�*m9��=r�}g�8w�if�ҳQ�n���>w�64Ѕ1�9������Q���x-^�����u����.�zx�髫�%w�R?O��8�RF��w�P�*7���sb�4�Ju����u/�!�N"^�S4��}~����م�tU;�������������lԒ5�ꃏH��^$BAK��E �hM��|��y����R�	�1����澝��R��$�z���x�����:@��/"IQ��!�6 B��Sc+t��>i�Ml/$��ljw��Q���A�jhڑ���s��~�n�U~�^���ϢFL	
�����������*�Q�������������������$&N/B�aV֠�������AS�:|n���^�z|���\����1Ok����n^NV�v���������?� =�"|�],�Ll��6�����7o^���_������!�H���������Og�h�f B&@f�)t>
M��m:w�깳��N��/���cgd�16�6ja4��x���` ��f�u� lA�!���l5��������������IW�鷩����T���H ���x�He<zk��b��4`�!ȅ��\�@�/>'���������^^>��w\�i״�KS�sJ�
k�kѥ���Fb�\�aTX�$N#�ߤ� �R�P\�Doo�w�$���{1n���	�7�n�~Br��S�q�V"WM�*��?�T�f��u��?|e����s��q�O�ՋI6�� ��L�Y,GL�K�<��sW�	tQKw5�>�GC�E�PA�B���	�u���h���S˶� ԛ_N�I,�{����]M�Vp����t��g�Қ��;.=��ة����]�j1�<��˟,��S�!!����_E���*B�B�"D�`3'�O��{�"�đ�[6�z�0+;��������BFec��tt"��BM������A�jc���$dߍ�άg�ͧ��p�xL���U�~���|+���D��/K+�̹�R~/��^
�NjÃ��؊�TLC�X*��A�_�>�!�?�d�jDý�gQ����w���TugM��U�#���joe�ݑt�js3V������z&r뭜:9TH�����-���w�Y��m�H�"�vpe=MDeU�b���NH��n����OQ[~�+@��yB���+[~!l����%�٧���.v��ũ�c�_��g�]MRN[z���SѬhΆkG�fa?.8�����q�ǌ3;/�^�.�p�Ep�؉�f�7a���M�;o�����̝1w����͞9k��)cF�Ӌ��VT7Vå'���e�Q
	%��g���;Ν��rނ/=A��nN�����Â}G���������
�7vX l��GN<yLȂ�c�}�ܭf�	s���6450 N=q�Ty%��_�b4��(�����������%��8��:|
0gG[Kӡ����VΖ�v&��lMu�ǘ47  �iAc'WW[ݞ2��n^��]�fkU=�h2�	KB��h<C c� ��x���Y�C�5552�065121�3����` x�����7pۮ���5wYrZa~Ycvi}q���X��U�5D�?����l����������ף��H��v��m����Fඒ9j[�m��c�nO��d��U�6��`����:�m�Y��*n q�)\$��!�+if�$&�)��T��\�!U��
�[h�V���)�p:8��H�:1�|&1�V�����*�@�\@��V`A�\Ƒ�d�$��@�B9��<�BǾJ�ON�G
�����dD��8�/B��`B`��g��@=��D�D8"<�t�  BDMy}eɓ�7ϟ9���(-=!�(���T/�:T��EɓK�"q�F���k}�]�+�����k ��wf��o<y����<:|���#��:���u�ɛ�&�����m��Y��/<eͽ[�'�Lȶ���|f�DS��h����%�D�؏��M��^wge탵���.��H�ţ����@�u�o�Hm�*e~�f|z���'w��_���"(ފ5Pv�p�;�#�P*h��仅h�7�Y)a�ƓA���xN��W���e�!� S�DHV���o�7��yz����o���TL�~C���(]��D/�}1�Fe�!�Yg�_ξ���꽗�������.#ǌ5��;f̈1cF�;z��q�G�� �=��?~�ae͟"�]X�/�g��3�Ƭ;���ԑ�#��F�4s��>~ĺe	��Ę��W,� A�gt�ߘ(����&�	�<6hʸ��B�/�42�}��q�o�H{v=��ى�A�n.��MNI/ $1��D�K��U��߁E��g0�*B G�`�����ֶ>>v۷-xt����Ey��ۺ;u�hc>��|��`���PKC=S�OM��p�@��K��m��n�������������kԄ���$5�D�n2���1$֡Rt\�������f	4��zx�ҀG��P������i�uw�aSvIc��L��y�Z�� �QE�U ��&E�H�������hbu�����Bqz�Y}�V����#��e2���Oe�����E?ϼs;�䉻��\غ�܎����y�*��蹻7��#$�Ñ#��FA�"Y|4G�ኁ1l,E��̗�����<H� ����m߰���E�f��9s���ˎ���e�̽s;:~��m{��%�l��+��$B����2O�.�-i@V�d$=q��ݫO��
������t	������w��"�[@ԣ��
��C�:���7ݸi0�$:���G���b`��e��#�vn۴j�ƕǏ�s�J~Q
� �����D_.��@�����p��K D��"+�k��f~wAX�DM̩*n"��hH7:)%9;�ғ�G��_q�܋
Rj�,��uꖛ'�+�<}����/O9~�F5v����o�wN .�(~��,KJ��7���҇�+��-y��>�x���;z|wCC�@��h���V���}�O��|]���װ,9�S~�����h�b��/�"һ+����G0�|4t9�����/��ꇯ8��}�R��+:�r�H��ୈ`J� :#�IALT�{�(��l��!��7S��Pw�7�&��>��[�'�>��X2���;
��OA3�\x\��H�n	���������5,lDTdTD8�9�^���������������/*uӿ�"�n�ZtU-����Ms
^8z��p?�p?�!�E��ΰ`�Qa�������]�B�ؽe�~tL�/��p�����af�7�ǌ	�]JZ��@m,���`n����VԀ�+�"��_C������!���D�%p��nn�@��F{��^������:<���������� ���b��%`���������1`tTp_��KŌ�zW+������������3b䤑�f�!�k�2�5lm�P��(�Є��Ehba��_ۏŽFF&����.�VnX�z��9�ӊs˚3K�
k�%0S�_K4�ŀF�PO�S%H�
�k#�{I�4�� 4�WԢ�����t�u�fƽ����(��JW∼�b�1|d#�����	q\�@���G%�Z�H+�%6��,�-�p��l �P! �P�"B�
���Q���&����R�-dv+[��	/��Z�I��bIZXȂ\��)�!I ���RIUaaivFv�s��]<�<���K������U������a�߅�����;��u.�E�hk���d>t��^�JLK�;u|?p�G7_g$b���=!��*�:�a*@�o��5�<m']�&����JɊ�,�ELrꓴיu��<~��r��Wn�^��zbq�����۞;�Ӫ=��k��U�z��wk1�O��t�������mh(IO�{���K�O�t	p�i�jΈ��oX:�ك�d�����ˤ5e����?��|��Ԟ��G���� ��6Sd-=Tn'��a�/��J��ћ
�]��$Xp�R�������J� -P�]C���Z�:3�ɹWB)ә������=�9��wֵHSv!����Z��72CG�����u;5�r)�j� ���G��Εw�e
�͠��R���I;����] ���� Յ���"G�#Pu��2Y�L�J"� ,d)��k�[����t-�>���$�� tqE���:�8��/�����wws���A)^RXPHXFv�٭���3�EU��iT[Ըp��hw ߰���1Q`dhH@­k	X�~Ŝ�!��� $�T�C�0��u!�c�PT|�+U�k�:"�@!������8�O,�	^  ��IDATB���?AHd�AH!8�g�V��;Y����ܾ�����B|���``mf`>���� *m�A�lM���`�� X�KS]yA���C���F 0[�#Z���ppBz���Ʀ?/�ΫE!4-aC+�n�Q�B�z|��Ҩ�����?���!�=s��KF���aa��|bFգܺ�Fv-]��T�������4e-S]�j�cw�r_4�_�x��=�q�w��[��2~�^T�l��s�5��8�@�H���5����2J}-���_^M�o��9��VN3C��ɚ��&�Ǒ�8�F�� A9�/�_*@���z�j�H����*�p�j� jkoa��!�{֛߾�gK%zk[�[J>�O��O/����N�9%��MI}����@�O῁���@�����,ڗ���@Hh�k��J�w��C5�E�ey%e��,���2[(�b�L�RAwI{��L�NT���I��?ucA��Y�=nC�C{�KKR+ptANQ%�ơq�����dU���ٯ���(���ճϪ��.�4}���*ܴ�W�/�ܷ_{~����W4FKR��3'�/]�h`n:f҆���%>�� !'����_~fh>�M`}�n����F6�M+y�%sa�*>CC��]j͋�ʮw��?��7Y5қY�t���5��5���t�*�I�WMϡ�x
M�	���L�F_
��2��F�*�
��o#TA�/d�v��])�TH!��߹*mIsgȈ5�S�T�����������w���ҏ�231275����c}#BÂCv��[VU[Y�k�u
6UT@Ex7�f�9����Q�T����jѼ�{��ܴr��)����)���������C�\<��ɝS��GF{����X��j�ϊ�'����;��2��q66�ί-ο�e�Dw'[3SCCh1&[+[Sh�~�#산h���qí�lL��4��^;��!Dyzc�S��d<��'a=��_w�/��G7�ӀA�u;P322���N�2{��#��z�V�Y����)����B╇E�u�Fnw5Mݗ�q%]]AS�7��������d����R�V�*zW�蒽��1���/�.>\�|���+��<<y�􅳗lY�}��ëVl�Μ�p�u�&�9eќջ��{�Ivz%@��
�+A�B9�/��u�Z�%�d"Q���M���<�������RPE_V5�V5V��"��^QW�k�Jxt��ѽ���t匳��#���"��#���K�!����FD�y{�W���=u���Μ8{Ƅ�+�9}����qyB6��$Q+E��BH�I��g�f�];�5���ݫ�]�r�ĕ;�¤��-�|~k~q���'�%W0E�9ҏ�_O}�}�ޥ�gׯ92u��e��f�By����&�v��T(�Y�k*����<{e���[O\��^�Y�{�����*�H;�}�H:̼"��9k�%.>t=�^�(�(��J�Zy�V�zjY�F������ՇV�8)��$�u�k^�T]�����?ZD=x����*�:�w~��C�J ~�¿F��D�Q�5J�F-���@�^���'��QF����ƹ��-��V֎V6���V����&��ff�6V.砀��C�mٶ���&�����*�>K�X��h��c ��n����!Aq�a���B�AQA���@/�`�{�"��9��U�@oX�����=�@�*��p����3���X7������vU�'�?!�W� $0x��V*'3����������tDL記`Gsh�x�5l`2������������>N������x�	x�`}�8��r����B�ꨧg��iivVMeY7�6���X�@�[>W��$�]�FfV�y�bePp � ��ފ@hmm�#Ə�<a�L aҳ���&-݅��:f�6L��q�r�;�%y��yRJ������bfT�;cgov�����3g��ͧ[�d�{�
�b���M�WT�g"���d vhL����Hp\��p5��D�{��@��<��휽�m<p�^���V�>^ϕ6	�lTr��<Y_� �I��B9P��SDO �Qr�J�P�+@ �HD��)2Eb�P��A8"9O*�Ԕ�Ք��$"�����i����,��n�rP��0R_zx��z�8�	�z{A�������_������.��O�?u����������q-� ��
�p���{��ݶi�C{�_�PQY������^-��/���mХQ���EO�n���<���)t������9wwL߶hW�֣�Ғ�y��(��}���#��>Lk`J~�ɿ��p�N�Ĕ��6Ϛ�b���{����x����o߁b�q����{��߹a��	S�E�ڰ�ҩä����g�o]i���;;����gl�;e��i��pdԌ�$�6���n��{�Dr�گ�߽�$D���ܲR�#RCaԝ��R�̾���/Z�˷���' �t�@(�wC��7�z' �����G��P!kW�:e�n��[���
���|�ܝɳ��E�ut�Dy�#�0Vv0cS����fcieoky�ĩʪ�����ܢ�*�D������O�հ��p􄈨 ]@�����XO�+�/*0 64T��0G{sc�!��&n�V�pk���/�r�v��A�{��z!m<\����6����.�n�>�_O�>������?�?�!+����fo�1��	��s43550 ��Z��+�ph
� ��A���`��M���H���m�W~�
�c��knn*Wg���cG��:b��;OrW�:꼻9M��OؑKnf����1c؜-�M�L��=fV-�U̜�Oky�mn�lގ�W���J_S�
���^"Jޒ��
jYTd�ϰPlDLh�X߱#<GFã���킽a�^hO/_k�{@�5{N�N+[��d=G�"P��A�WP��B��%�I��^�?Y�L�X��C(Q�$j~;4V������"��ʪb ��L?��¿��C�[{��x��j+�p�i)�߾�fQ-U�e�͍\���T��dm@A�Lŗ�x�N��G?]5S�FV�
^��^�}fۂ�l^<%33s�Σ�Ο�~w���c�w���}����.�t�Fr|bʥ�W.?������v$V7-�������W�RN$�?�u�2�6�(���͢�2Om-�q���qb�K�7_�v�����\Os�^�@R'T�	4�%M	i5B������C�n����*���G������ļ��o��g���<&[�Wȅ**���ݛO������|�,��@^t*K�_Aا�D�"���S���Ұ�u�����U�vǍ�>t�$��Xw'�����������T���� ]\,X���,'�(=+7%-+#� ������&=�;�O������|������A|�n0Ks���h�B@  ���!��l�q��F!0(������y@��:�OB���?A�J�hPHdVQ�w�������&�� ����v�M��X�@��W-LAk0��������A�?Bau���X �,l�,ԭGX�k�y;��6��b���`#}�������CS]�`�����q�'Ď��^�8t��y��<�'�Ӻ�����m�/<���o���g=���̩彉��}�t�-������[��A1񴒼p�I��c���FR�':����2zWHk��K;x�̑�N���~�� ��=�/n��C��!l��8�z.!�Aا Y�2�'9B(\��_zE�_?�,a���
�DT�X[��GL/�.��)|�����k._?{��I/w{k=� �o]W�W ��F�� ���~���?������)����cV,��n��]�6>��v������,���F��*(��� B����z �({B�&^;R�tjϖ��'�]�c�U�-?s<6���;�W�9����|<�奄����sw樂��H]�����E��q�����Gj-.|�pq7�,��⦲ӫK/-?�\�t�t�?�����ΞߞR��b�ez;��ӄk��.��]J��r�Қ��j[�ܑH�/_j�Tƥk瀃�޿��Ety��iO�����c�VA^.�A��W�ʪj��:���	�PI����X�"TvC�����W�E'�O��K��[ /��ݼ�h��C���_�r��3b���E���{zzzy��	
�3k��+׫�j�s
J+k@9X�v�� ¢r\��2� |��pFO�����3*:|XXh�������B荄�|����նB�! B�� ������D�@��<|\�������O6S9 ���X����>-M����-�0 @ha8 fM(
�sp�[��������F�}[�	�}�|0x�����������7�yF]QasU%���\[K���*B}Q E����|46��wrr@��.�PHSPY�m�A��tqqA"Qa�Q�ãb'=�(���}����z���EV����^�s=o�S�n�L\�\#t:���2z���K$�_ne7�]���$��}xX�8g�aV�<�����H� ?׀��cM�V���O-%֥�9�it�S����Б��H�(��S�f�Z��x-G�(k�B a��I o���"��#�O(�?A�a�P��Z��k�B�L#�o��+z�*�p��e�ߟ>c����B!=�0}%�~�`���/��m��@������>Pp��i׮���������WL���d�H5��!(
i���v K��3�K�\<{7#k͡cl���������?�����}~��=.m�㨯=�ήiy�_� ��BJ���51���~�[�oڜҢ��Ą3ۄ�	EgVU�Y�ta3��������S�$�^}��Ƥ�;������w�'��H��<�VF�ń��o>ml�3�(����{-���a�5_�nnj(+)�>mRʓ$1��e0�FKC�㇉e�c��Փ�,mɊջ��I��^\�H�-��rP_BE�� �N���0Ut�7�#|�W�N����SCc���1X$���˫o*>���iӷn�~�ƭ+�n��=��/��-�-� �5 Ku�˔�@��R���:}gL;i��ᑡ!XoO��-8�6q��@9�y� ��!��X��w�!����rwB�<\\���UT3B�O�U��8�»��Dd�t&T�Th��f�y����y��}�==����������F����к���{�b� HW8GC����VfC���BcS'�x4]������#&#���� ��"�Ԑ��I���������n�8�ͬl�.�.($�����O.�W�����	�
����|������<�<���?[tx��Φ�_s�N���X�D��ZWԼm7�8�u�W�w�Yw�zE\N�������Th�w^����::�z/�6�GƖ��*�n�9�yd0�i���J,�p�G0&b�������j�P_�/������U!E ���&*P����X��}A��S��uc��B_�z������q��s�N<J����PX� '"HwWP�}������ż��a� ���;F��c�"�T�H��mڸ6�qbK3���߂��d:#=7_�P��r�Pg!W���~;f����žc���%�y��TWY�@L��`2[��\;�������5�I����7�:����ˈyt��]�:�j�j+2�=H�u� �p���w6�9Zz�@Ʃ�׎g^>r~���'�g?<p|'�G�����5��طxǮ�[vM����B���-O�E�~=r����r�����(�����I����f[Z�::w��>}�t�F�1��<�p�*P�с��#�:@����Cs��v��/ 
�4/�_o{��&���\��}���؀��P���áI���VB�AA�! ���~����VJ��B�U��T2�a�ll=�����'�:i䰡!X�+ሰ��[��rP7˨�n�Q !�r�� |1pO�.��X���������	��c�n^7�/,n-������&^+��W.�������������Z���
��Pܾs/��Ba\��,�������mM�@��X8;@���@--@og�
"�l��k0A�0�07��1������[[�� ������6UV�ʫZ*�[*kZ�k	�u- �V ���7,l���"D ]���H���8�@kP@�O�9�"A-�g��Gl숨�1!c<-;y+93|ƶ}��ݳ������Uǟ�Xz�I����j���Q��8��������m�ǭ�4qQV��,z^CK)m�`#Q܃c+O]N�t�2��gJ찌��7Nn?�s���s�~.��h8t�18��Ż�U��EK  ���� ���E��(���м�&����a?� d�z�KHn�ԕT��g�;���'O���#D�\1pz�����s��*�ߦ����!��?�������{vm۵s���;TQ^\VV������@E����Be'����&�_��q�I�����
�$��p�+�ya}a]i
�"�^�������#yM9�_;���PI#�U֊��.x����_k+D�>*$��|�ʕ
XT\]ޓ�ۧ��Zuu����ݸj�򅗏�v����[N?XP����~����t���[O]{h��}�g/�\�W���@�\X.�IzVm��4�Y��v<�����>K~t���#���K���72���[�R��pi٪+7��S���<94�^ڮ�P k����!�f����~_�֣l��<)�%�*(�p���B"��0(�?A �-(�/��RR�gaIesI9�I
��v����`�!a��1##Ǎ��z#����ۛq�4�[9�@3R�Vb���B�,�ps$����	7v��:q�v�qs���q	�F3�!,*��7
~B��՘<N_�C����0��-{��=k�����kSc�+��h������ +��ɵm,��͍�y�x���5�@-8d �脾"16hbjhjfljjeddok�u�nn����i,�n*�n,�i��ÃsR���+�~��'�,���X�ĩSfN�030lԽ������Jfl<;��]�v�*e�;_��rVvK;���dRŰ�{�x����>���ɤ��N1IX��ou?,č�����VG�;�AGx�zz��������u6	D��^ؠ0&�#r,(%��<V�7��,a[���@
r����R<
_D�I	Sp0�_�_���B����^�s���سi����\�l>a놄{x����ԁ���������!�!��w��E߾?��/g���>ytάi?@�`A��!G�!�|#��DU���*d�� �%7�s�_��_޶p�FQcEA������*%dK>HԿv	_w^O{� �!/oRk��h۵��.P�_�i��twHxԆ���>����囧�^=o����Iμx�qvqeim���흙ee��<v��ދ�v�;�r�>�g��$ڗ{q�8����XFgQj��|��E�ٵeŲ#GČ3�ࡽ6�6bh^a^^a��5�G���h͖��|�Hɔ��d���D�&�e�\E��o9y���7�Ե�o>H������a1#�MEr����b躨�"�/o(��U6WA����G���0���������t��,,�@]�@���x���`;3C;�Av����-u�x�ؘX�X����b�|��7,,"� �y-俁��џ�O�?�w�B"��L����]���ݻ���}��^@;S#��w�!ut42�T~��H	�#��:z100e��� Ch��A����\��,�a�󜪬��������ʺ�����F�a]S��KW�k��N0gw7��Z'���vsG"Q($	 tC���h����9Ѐ���	����o�T�y�t;��v1�*hm���R�y��(�u�qߤV���m9M�|�'�嵁r����$�*'�5��X��RV�����������C��Eb��N�>N�An�#�\�N��@���@8s��e;�UQ���$x���%i�H[9�G�)P��堄������B]�� �U��#�r�7���"Jnqz+������k���ɸ���`p !����ǽ?Z?(ҏ./�_������!��[�w�E߾? ���2x�0?7����a��m[6$?N���,(�kn�3X,���_ �}��B���#k���`(_P�>m����LТc�#�.9�'�H���rS��KW�:�x�ҩ�{+	���V;�ףY{�T���sw�:�NI#�i}�����t|�u��z���S��+K�<L9����&�߱q����5U$qy+�*h�nen�w���|�[�j��}�On9�����6lnb�����'�;�q��3��1#Gƌ������;fX��'�FǄ�`#��Ō��?e��3���q֊�'o%Qe�t��#W�d*�?@�{�P���IAU�\�-�vI�/����U�ç�p�ƽ�{Ii�Q���b���!��
κ9i{o���6A���(<x�DA	t]4��:��OWП=e��g�]>�����Y��ٚ��,��0/����������l�[�����0,��m��n텴�r� [pD
��:n\�_�b2�I�����r� $�$��H�]�����L"�߼i��m�����<�����������@[��`��ѝ���v��!5�_B��22bj��q@xݼ��[R�S\�[Z,��+�i(��/oh�o&��|����������F����,Dy` �0G��`�p��-^7!)� %�2��[I�o�� U�-��RK��3ڪ)�����Ʊ��6<����F��%J^����\��n�%�����{`\=��Xw������������ o�!^�&�n��(o�`{w�g���NY��� he)[�r<]�S��
4-,a#���H�R!]�a�;���6�.��"'R��д2��`��-���y5_&c
Yl!C(爔l !��O�|�{��[w/ݾs%6.����l��p�`��-�
��������>���/����O�������qv����������ݹyӺ��&�9u��(���\$p�6��_R���)T"��]L`а�j�D�Ӽ��}	���B�͓h=�Ng���d%O���ard���IY	�i|���'4BQϋ�w�|Xr*�i兼�E����Pǣu�w}���c�JavzAnqu5q�'��Oz\T^M�kdR2Gɖvl�{T��2��n�c���9�}���M����v0���wʧ��c�~��^~�޾�~��X_�/���������?
<���7mѡ+	t��H��)�R%_��C�H����X	~'А	����OݮP}�J	E��Pʻ��k��_����=n����7dݸ��?$6<j����-��Bc���������^^X?���Ƞ��C�N�s�]t
T5V�j�{�ɩt4zʌ٫��7($��f��l�v�ø�;Z��r�3�65��t����aQ�AޘpO7G7G37�����u�� ���Ζ&!�ޡ�!{v�*(l��kil��������[�'|��H瀐�,�F"���u�=���1{�����@hQj�ۃ�-�@+.�B�͠8�ڛ�56��Ah1
�Z�@�e�����[��l`.�c&��}��_\�R�#��Z+�- ���5�-�-�f2���xk��������������(��⬿:
465177��]�r�u��O��(5/5�<�WPI*�g�4p���+��Z��DS]G���h�F�|��jk�v4�C�QI�03E�
��+\\<QnO�����?��d>�3C�������cl���7�p�cSo�h�2�@J�x���"׼���o�0�J�RÔ�kfv��=lM7S��K�t����__�+ح�� B�LaE
�L�/����o^�����N,^2�����Fc���!
��@��o�'���@}pG3#'�1�����'��9}��s�r�3pu<>G(
Ă���n�B��:U�Rh�%K,u!U�6tΞ�e�3����o^-�Yw�ڣ�|���kY*-���|E��RAp�T)��޵��l��N��l�>!�O��5vh���H�E�O�Kү]<
�Is��	���q�Љ5k7��wt�����'g���X��UT۰b���A��n��mS�D3~�v��7��,aA(� t�g��X_�=�/_��.?�G 
���q	�r����bY�M�i�G��ҨTݩ�t�#Wu*t�+(S�)>
۾�ڵy��qk����z��n6phpx�afmw��#lN�.�07���������BS�%="yxM_��@���>N�>0oo'_o�td��Rl�Gd�[��]l:2�}h(v�аɣ⦎>iT���aㆇ���8�e���v2qwǸ�[�!�]�,ܔ���.hmh�SE���_R�AHbrA(6�� �+׭9~4�fmgfmobj>��v��7�9;Xe���ɼ/� ��A�,����m�%�@5igg� �;"�e��\3~򳂊����fbEske��@�%�֑DB3�v�v����p��������f���[AK20l4�@xxy�]�i��Sg,z��05�@XTA(���7�Kq��f�"n�I@@��H5P�>M��P���-M3����"�^��_���g��Δ�W��b��Qo��� ?Ow�aa�l1eg��b㏆{���}��]|<�&,�yv����M�&֋fvO�U�������� ������������в;���IQ�A�k�э.�0�`�>�!�J��
!W��T��-u�8Ș��ݧ2��޽q�|N�S6�XV�c�h�p��x:a}Q�8�WPa��B�7O����!�����3��!,-�'�SS�ٵ��0���*7/;+�9P�/������?;8������+�s%�H���W�2��7m�ͅ�>iP�x\����U�������<������W�J������"�I�|��ߐIT�h���ڇԷ��ԍ��k�J�N|�z;7#���A~��ü�\{�¾�HoS�A���|��p��5w��;}��f��v扂cQ^Nnѡe4��{��ϗ�N�{��5
��
��[A������c�<P�@A�������*�o�\���<�*h��p�Q�K э�h�;$�Ni�Y{�>о�B�R�|%U��(?�տrڵ�mvC{����n<(�q7��`fm9�������z������9���������#$4<@x�������:��J}-�>�%��:N�c�՛Ď��!�AA(?g�����=4�v*"���
�c�#��"BFń�2zh��� ��Hl��k��S\0:��m��(GCc�{L䄴̺�Rzy-����!�������k��%<� $S!)��6�%յq�F2�q��	�
���p$���sw����h>�����z���x:{  X4��tspvv�#\�\l��v;kavy}	�P�B�l%U�5$P��Lđ� «����0�;t�q ���� CCp��C�t_�|��5��L���*B�����jRe=���Z��73$��w $�G�ն����f���"k�+��Mlu=SN��$����H���}*��I���������Gv�6Aۛx;[y�م��B9i鮋��/hRճ�6p>DNݚQ/����g���k�<��L�r����y�G���t�*zH�v����v:O����WU^[ $���J3���K2�J�KWN���� B/�"���O�ǯ��@��/��vx\�����.Y0rD쮝[��>njj|���	�ť%m]��*h� _��P(���xCu۴%B-�7�c|מu����vG2gܡ��'���νZ���;�]7�$�%�v�ۜ&��GeG�5-���������Y엟�^I�������)���<zx��E1�Ϭ]�j��#�h�[	g+�9���"��#4c��O�2���/'�?�x}��v�ȅ+����N�����y�{{�y{��ѕ�__� x��_�o����~#���1�z�͜�P����D���P�Kq�}�mo�("�;��_�����;��N�3�+�q;�ė�'�\�O��uEy�Z�401 uy3`j<�4f�&f��ֶ66v���A!�"����^K�8O�����-q�A�{�Eb"#���({?/��H�Ic��Ң��sgp�rs�E��xD�Ć�����=6.��f�dRM!W�T�?��.�=N-/�`�UsZ?!�����cs� �� [	�}i�П�X9:��Z!ܝ�\:I���<M �S3Op�f���"=��%��[W�9�W/<@��u��B�����6N�ذ����5͕��"��D�#SA(<�
�Je\���o��M���q�P�G7�ڀA��z]ܐK��Z�z�艳Ss�d�g��6�Ւq�����`!�.�'��ɜ���V�cՓD�X�3e u41Q���oV�<g�n��-`��*�Fb������^��H{GCg+C���������h�����l���/���^�пL�U+ֺݐX�In�Yx0y��������6�����~��3A����*:h�6�����n���𤝥5]�v� a]K]AE^+Ob�[��3SҒV�Z�u�ڻ���[0�d��b��p�]����Q��%ȿ��_���O�B_ooO��ё���zp/���=�Ë�O'ܿ]WW�iS�\.�]TR��h�C(TAE!W	,T 9�6���륿�-��0�4l�Y�9ӎ�-��\������&�\��-�i<�ˤ����h��4/3�پSׅ.;<�HB������q�Do�����Gä�d�^�znӍ�ۏ�\� �Ĝ�#o%�Ć �$��r�a�����>��¤>/�O+�Z��\�{!�Ί�;�m��KW�$='J�,>	�ND��������xxx��C5VX$���ǆ�	�<<}��]A�W1�>3�zX*h�U a��2��z����j�*�٪n������o����fv5U��;��ۿ�jh=e������|��Ϩѻ�zt�^����#�G����7C#���2<�`� #�!�������A �",�n(��)��-�ZKq��nr�6<4f���/ ������z{;��&���{�x>�B,\�x\��3�A��A�����+�GF̚<<���|����OmR)�3���x𰰨�Q� �5�=�?/��lj�B�P��l+8�0zxTF�3��i�à`o �;��h���-�Wp�q�BvF��)q�hGs$��n�����`�v0�5���1<�_��T��Z�RO"�A��G�����t[���X�!(7.^�d��c���V�O-|�U]RϨi�W�uK^C��T5�V6W�� �D��)yI�t4��8���!���H�6�-��q�t�P5�����Hw�
��p��r0�bm ts0F9�89��<C"&.[��V�c�\m>��'u/��}�6��q�˜]	k�&���/1���7�$�~!�_S�����/�mf�Y� ��n 2y�o�d�ǩ�o߹r��U���XGX�,���p��^CVW��V�'?N>y����IvN&(
y|��*,.R�i��=B��"�C�B����|G�֞�hG/���6i�3�k��=��7�Nx�<=�x>b�ے3����_��v"*?d�*�l��5�>`͉GTMS���_���Й��E�n\سkӜ)SBW��r��Ε��:�18
{'�ڎ}�7l[{�؁�{w���ʂ����l\y9�iɡm7��E͞W'�>�X:z�)�it 
jP'�Q�F�GF���D�s�y�ña��>q(���8����_��������l�+���
�T��/~�|-l����7~�Ρ3�{���dB%�kɎ�#V��?��aťڇ�c�ֵ��]��u��������Kk��,�!P4��XZ������<�)�l )�i*�)�BK�a���=�|CP~�n�Q>1� ��P��1~�w�������&x9x��{���)<�"������	�E�b���ėgk?���B0^H{��Rz^�BO\Y����O��?AH�z��@c?�̳�9��ڂS�fr�G�~�����6��-a ������V���.�55.
nuu�bgkbgoa�`k�ah_�_DjneNESqCsq��T�" �����ר�����̀�Cz��Z��͜=΂�Q��=˫z���i���]���6�sk���kZJ� ��-��MY�ۑ�QSO�Bk�ӄ 5$>��nf�Sf-��aTd!
�B]l,�"mM��&h�������8t��e;W�7ggR�H[��V���Z�1G�g_����c��m��/�O�o=�A}e+�0�/2HA���!�&�vb�����(W��w�$j A+��Jo��,>��*���@x����'�_�v6 ���}�et�F�C����/�B�S{��C��� aTD������Y�|��M���*�߾}d�y�
�J��sE��8���mת����6O��q2?p������UZ�Z����^k�>iE=��O���%I�$K��[�m�V[��ο�n7y]y�W ��筢����vmX2vT���;7oߵ~뮍�w/[��ѳg��޴c�ًW��<Ph:�dpnWE%�Ӊ�Me��Z>-f��ZA����q�N��g/X�i��K�/[�|Ɇ��Ϝ1k������]��mb�j��G��?�`ﱇ��'��[:t�������itU�nf��rR�Bv�/��V�G�a�/�﵉��Љ�[��j-I�gf�S�d�����߶n7����2,84���ro�?B��� <v�lu]SI�������G E��'�L��ذ8t�g@���?���*B�Ct8&:5<�sX$&2�=���T��hPA���`�ްd��E3�o_�9n���w/�%L aC���#R8��^�˷~B�����+-lmmm�oZ����� �!FvvF���~�{!�9[��"��]a6�u#dM,-�mLm�m�ڹz:{��2����j�
j��Jpe��J�
�?q���������,�! ���ll'N�6e���c�</���x�i%��2�P���|þk����M���W�$r{���&�����,���eۙ®V��@�GGC��y"�Y*���bcnol��Y��tG�@�x��M��h����Y~e����k2�?G�8U��z�mm�k�ſ��$o�x~ל�'�k<��dv[ҥ�O
��!W->��I5o��!��"l�5��D/^k��F�^<�{���[W߸uaيy B��U?{��}��E�S{������� gN�v2Ҟ����� ����
�8��u��������/�g��k/�^B
���^���#��	��9gɎ�w���ty������⤸��a�ϗ)>WI��.�
qw��Ni|�4��ٳ��LO/۴��������qFM�vR��gx"�G��Dt���
%MB>A�k�ӹ�;2q���	�����8Twu1�?��艣�l�t�*�f>.rt
Ix\��3��g,;�;�+z���T�[�����!�s9��V�d)�2�_*��u�7�q�hm-�#Y��y�����'�.;�q:�Ax�M"��8tú�w�_�8z�z@`���l�B##�! �����MMm��@ъ���<x�DiE]~Iuniu^E�e��	��a?��(�P�_������
�����h;�����a������v��� Ģ���������8�v4聰v����	��"�:������&n�L������O��?AH��A��	�Checmekiiejn1�� B3�V�м�fC@Q�:[�l-�,��X��I�AF惭�M ��N���wXrfEv	>��1�������������(�R��|��e=��� �z{�Q�Rp�� �A�Ɔf�f��;~�ę�&��V�8~��cX����B֥�u���O�����R�ۏd�aD�-�j+���'֑���:����iᨚX����+�U62	t��gّC=�(W�p?l���?���;�c��V�J1 �o`6t��e{�^+�p�j
�o�n��uW���ߡc�7�^�do��WdY7A��=���œ����<)T��×|O߃�㺅XE��|���0ɕB��L�+B)(�b��j�@-��r��ZW\��*B�6�	�����^���-�(x]�^�������m����v��~V��RHħ)�{w���z^VR���S:���r " �H�э��n��*�R�Pup��1{�n����h�J{�L�3u��D�賶��q��KaS7_}�>eCJ)�{���m���v}=������f���^{&�~��#9d��S�uw�Y<G�^�Hg�ޥ�5��{�����
��iB�''4�b������/Ly'M�����ml�J@R�(�W��F�ˇٸ�iy)i�)��R�S���ݵ[WwG���{��N�Ge���KIye��JZa#��,n�t���L�Fi�:�{wPA����}��K��z�
�_�x�,�]�^�z߃�O�s�F�6h��y�%�׾�k�y=���!A1���-p��j����������	�p������~A^�{�-(K�)N�-N/��,��.�/��>�8�af�2�����C��tr����65����01 �!LP.��HX?�|�zaV���VP � H�;
㊁���^{���Z]��A��9��ڦ=o~���O�?�a+��ֱ������&����c��v����Bs�.�� �����4�:��5��_�+��Ղ�_�k�McK5����+���CL-�u��]��������\\\F�3f���S�dW�x\�<y۩��F���Ͻ�S����]����1{"w�'�
�^!��H�?A�U�!��dsm��*8�v@@�}P�QC��'�:g���bݭ��m}=�����=|����n��g˷=ı���
�d�/yOK �⡡вN���*�,��j^�!TA��R׏@}���T!x��R�JeSD
�D�e����G'N �ो'��|�0G����������5���ڱq���������[=����B���:��]���
�r䪃��w�J-��������M�|���j�=����l��M�-�-]�ꓖ��0{��V�od��,��Q��Pb��:Pe�u)>��d��W��ͤ�Ė7t�;�����D$��)V
U/9�n��#G�
��|��R�5<��MU
mN�;��#Y����$�%��b����>pԸݯ>\��`ּ��'/!ReU�
���Q�̮���5I�~F��UB1�B��Є�/ي�m��W��KL�<q�Vܣ������8G���^�bwY�^���bGd�ʝ�n���9u�VXh��aqHW�������'�r�pw�Ơ}}�>^^nn�p8"08�����>/��*�մU1 ������(?l(&0�3(��'�����haj`bd`i
 �0C�� !�P� z��NH�%��X����a����an���������7w�x����O)��j�Y�޳�|;����
8cc 45bjNߠŕ,�zg��C�h:@�bm�nc �7dN$���o �h�!���Y�:Z�ځ��������������X[8��A����a��i���R�[&.�0v�<����3wq��ξ�^(_�'cܬ�G�Uǌ��(��YOQ뮎�/�r	<e3[�ZP7i�*<E���X�q;���z{N7�ބQ[�
�/�������� tń���yo��W��^W?TS^3ڿV��uQ�XN��uc$���Đpd���BE�!O��+"e�D �qhB9��%W�>MKJL�_�aٹ��n�_�6u,�����A��z���.:�����-�'��ѿ��=�?�O����!P������Ѓ��%>�����K��}��(00TmU;���2�<|�zB���AK}�%tj#��)��ږm���\Rט�'�E�[俑U�3��h���r����&���ަ��PV�V�����qymY����JK`|�P>��o�H�V�����6;z��K���7�/l���W��U�9JS�f(�4��&{���eJ? �L!��&�� E����.��- ���s��\��i��2�@���%��̑��M���t����W=� �!�)�4�8W���W��S�D1a��	�'o��Xq�鑿�n���q&��x�|�k]�:r�]{���O���
�zF����`Ã"B�#BÂ���|��"2zXHD��S��.���C�l�0%�in=�'h�����OX�����H,�`m5������>T�e}�]���_���l�`V�f����A8j����E�Ԓ
j=��'pZ�l2�������O�ۿ����W�*	�M� �L�%�B�t�1q�2BX��#t�2CZ��Z� �t�����e�,�G{������g���ʬ��R\vi}�U�BWG��K��k���m��! �@y���0��@{{�{b@\�(T�\�@A$9fܤ�f33%��IAӑ��6�Φ�E-|^�zRć���v,mծ�yk�4P�C���^������h
M���j�<"_��Q��O���̒�6��Μ�p�Z ��i���S�M�5������f�AZ��e  �?�:k��+6�ɫ��3-��5�{*i�PN�*�rUAH���PJE�`![��;螟���yʿ�P�-S�h��6@(U>��Ԃ��z��v?��o�W=�x ��3��p�+B�M�~
B~�����]����������h`��ޝ�Ғ��ۛ���0?/33�/��*B=�tuG�XA�z7m�7�%U2�;w�(��ܥ]�?�i��ԡ�z!m��Z�+m5����\�ꌛ�m����vݘ����I�ʞ�f��|$knݻ��#Pھp�Z.�w�#��&�����������o={UХ%*�R�Z��x�Dr1_�a+�t�"����.|M�@!�͡� ����(̖�>k�Ӏ����$P�LA;S����3dЛG�FWj����:�� ������,������\N�|�Ʃ���]#�����V���+S�Z��K^���7�ã�#�G�9bD�ȸ��aq1�q1�ёQ�!�~~�¨�8 �ً�*k�%U��j\qG�J��05�ef�sw0tl؈�ё��^S[+C��v�avF B�������Hg`��(t�pv@ؚ�A�q�Ǣ��m�޳f�*)%�UҊJ��!d0�-]/B�����C���?��df_<q-�uڬ� BW7t@P����4������������Nź9�;Z�ٛ�Z�C��z�:[�!,L�A�8� Z�~4Ǽ��������������'����5f�2�k�Kk�˪��jA���j��r��b<|�7��P�/ ���h���O��!Q���'��2oظ�)y��bz�{��A������E)�L{��U��|uҢSU�ӊ�ѫ����N<C�gJ�LQ=��S��������ml�|�]��&�>(���e�r��:����hW+Z���'��-44r���w�/8[P�u�R�ʝ7�X�,)A�"ɔ4��&o��h�6�H"T��5�4`�B���/@��VV+S,�x�ૠ�3�N
[��^K�uP�*��@H�1\�L%�ص5�DB}F��#��\�|�����.�v�f�^HP�
� �������k�?�-���
� ����� ,8h����=�v,Y��ʥiO�����ڠQ�lv~a�R�&��@���tɡۄ*�B�/z�&���x��5�cV�9�����������%��[U�rFό�g/<�������2Կ�Կ�տ%��'��-㵖���+w�_�(KRcGD��ZJȒ2������օ#I*I�23��d��p�̵JZW����Y98ɽ���2n�;w��у��p�InŶ�W9��4���*g�����b���c'L[�q��7/_���m:-���.mo !M����ShXrh�mh&t�T�^{/�v2�<�K�Z(5�k��=K�;[�eK��+e���FYX��{o߾�s�̭Ȉ�ÇŎ=ft�ȑ��G���642&*22<<,8��?X���p������5Z����k)�#�ְ�e� ��hS{K�`��ѡ����������Fv6�m�6F{3h&G[7w��;�<�lg�lg��?�5(z���}�yfmy@���i��d�?�?�a����z�5 �~f� E!(�����������1���������f涖��[@�%��l���Ct23q0lkh`9��|04O���`3c{+3{G[g/:�ᳪ�My�-y���������}'�z<y�����-���^H���;�������ᭋ'�=��؉S&L�7~�����2����-��_�T�m�m_��TB��+i[O��ӿ֐�� �h��FƋFf[#[�Ē���XC�3J��]`����)�	>mt����_�v���S�.�(KwWP�zz�!\��a��mw��ݵjKb@����ױ4�|Eo9(W���*TAtJ�A�E���l���׿b�����=��B�G��h�I6�C�Hy� ?���0�������ݽ�����vn�C��ޞ(}��!P��^<w65�ɩ���͙�J��g���MMM<�{�K�m��D��-K��}I�.3���ҷ��~������iy=Z�+�΋هi��n-A�˕��� � B��Y��B+��6K?��ƉU���w��v��yS+H�R����C�`	?P8�"�,)%�9����7��>U���Nf�Vo]�]�,1��Iⳛ�O읱lIrn��C��O��>�B��Դ��j2�K$����jhL���v���"U��z)���
�P)��n�4zD	�B����a��@T��M'C��%�M!M�#��X]/	��g_��{9g��GD��Ā��b�����F���zHPpP@ 4������ҵ�5��}�ַ���XK�X;�a�������'�u�q036����t|һ��Zhc<�/�%����ǭt�156��D��7�G�:�^���g����a�m�_�B�_Q׼a34Lj���Nή4h�����������������1��na�=��&��(�< @h:����`���`S�Af����z�x�~^�R\ͪldW��U�Ԫfrm3�����B�m$^�O��@���7@?]�Ey�� ����<}�O�1q�¸I󒲫Ҫ�wUQn��?���%y4��z6Aت����$�j�6������~������\�%�J;����r���+ 3L�@�p�����쬽]aX7�
��j��8�f D9C3� Y\~�7m�7v��"��әS�n`��� ]��.j}�ڠZP�a�D��<9�bR�M᫩|ey=����������c��.�@ d�8l[��$<|c%�֜������ib}]E� B{;@ �����.�=����/���N����� �+¬�M��BP����烢���T�ޡ_]H���/<�.lk�K���(VP�/8��r;��^ů�)%��ۯ�V�ğp����_ i�/5��m%E�,}�M���%٥�TRmmyF\\HzYyz1��UP,���W��	�3��2�L.�ƙÏ��OZ?Oۗv��y�̅�I�JK����:{ z���̒/�5A���T(�
�P��T<������7*ūζOD���P0�����@A节BIWB��.����&|�ly���T\�����p�P��M��h��P���+��E/]jp�Ј��߹��s����ؐ���P��PlH�OH�op68�/(�/��?���?@�S ,Ǒ��9�R'�q3�uF�06p�vB�����3qq�ss�����<�a����A#���(';w���3���8�{���Y�zu�Fy�������ϭ?���aүP��P V�-��8�{ﾐ�� 4�67�23�2��Mhk:�37� �4֏,�!T���<d �y 8��6!����ίma�uZ#��'�����x|���isN�5?&n����o�6����s�`��}4��<K����G%�G��2��ZZ2��Aq4 8��涏Y-��g�J[��N�J�����y���n�7�dd��
B�L������������h��6��f��F(����l�B���H�wd��-ۮ�Yp���&ePV���R�J�D�_��.[HApt�?�(W���7�oկ~%	���F�_5~��t���O�?+���9�N�H���\�\�g�[@9�k(}����c��_?w����`�V������!������������� H��޴a��5��M�|�҅�������F�Db��,��w��>��P7�� X(n�� 8�H�X���Z��U�y�����æo�y�nU�(HS}ԇ�����;	��a�7?(��?L a��>bD���'.^=+&vᨱ����1隥�ץ�d�W�Z�x��6;�����LʉcǓo�I~x��o�9u��e�]=[���o�I	t:�0����%��$��߶6��.���!��N����_P���W�<�Xث`��,��4*�����ȖjA�n���5x�������}��͐�h?_���b1����݂�p���:�z�zxx�[�ܥ����O7
,�W���2g���v��qp��x#\Q�@A#��fec9��������Z�^�!���������3o(�-��|=��C��?f��#ϳ*�*)�e�z<�;�,^=�����'�?ۏ�oU^���6��P[HT�O��V�Y�{�ޅZ[[������[qh:��z�����x�� G�!p����	h1&���C�-���@E���3fF̨yEU�!�i��4�jZh �z���ka��eu�Wo=6zRp�0l����	bC�9�Y9�X�;[�"�]]0�Ξ��Q��ħx�Lr�6=j���y�����j�3ք�و���*j��b����3f�֡36��6n֪᳖MX�f�%s�l�&P�|��嫼=�}1� 4���BwGKG���u����p�f�vvE��ƍ�t���q�6���$��_q�PxR�HBK�9C�bH5�Ц'P�~!=(2h�h�Z|��)
;]4�F1��"t�5�O^�a!:�k޲�|.[�g2���Y9��))w�o[}`����-�7�a ƀc����>��`�O�e�ߴ�P���AA���e�9�01�̩˗.�~�J������B����TUU�OHR�z��Y(T�օ�n�~��P�R�z-��"��*�����\�(��iZ�=ଂ�xGU����3TP��_H����݂��;�9����6f��ȸ��Qq!��E�M�6)&vJt���o�@$�B;��L���gl��5���I�Ӊп�V]Y�\W���yҎ'Og��I�u~�`YM(����f*�Ca��$&����V��`�T|^G
��b�;�m�Pu;G��Sw�/����|%4�����׈PQ*Bu'C���zB���_}�"0C�M<p�������1���Ƹ��!��������Ƹ�"�pDph8x�<{1��,;�<��<�Z�X�²:bY;�9�2���k�ǌ��q��qFc(�SP�'������?<:���D�Az�FxL5eL��aᑁ^�x	w�����!>��Â���V^.�A>>s�,�/l(,%�V3�x�����X�Z\c���/��_�?��O�]�ᝤ������׼n݆�#G�����A�����%�����������H !8e�YA�0�` ,ĺ���ݶ��l��C�`A�C�,�4nڪ�-O�k��F���T`!�H����)�k]�~�����������!&6��փ���X p��0�9{���<ʻ���tb���SOJ�g���R��5���ϛ��X�-�YM��-홍�l�,�Q����ǳ��J2�O-k��^}$�E��B8���np8
��sD�X[����:XZ"av66v�111���9{Gc��7�,?�̐yR�PL �t�����-m�I�A��!��8�z���������K����[���{��l��\�TR���(9l�P-�%����/_�KK3n�<���؄�z�t� �(�+T~S�P7��C�B��`�����S���(���J���ٳ��J6�����$�\��[�e�H�B��"�k�ꭤ탢�Wq�'��]��&}K��Е�uy���L�w�ԯ��7�������}���h{W/��7�����xzx�0X$
Z&�
a��X��);0c�]�p+�TRV�g�pYUbasCcɥ�Ǉ3[�{�����j4�����P9,P�x|�Bӡ~���������R)�����K�+f[��O����w���ҧ�.3��VC��&
v�4ݴ�N(�v�ۏ�$F��q�߸��y������������`omcefemag�;���no�	^T aV^If�삪��ڂ
��hi�����!��k����#c"�|�������A�#}�ܰ��@o`��9�����=4hL,�؏D{!��|]GFx{8�`q��nV&�c?v��������:.a��'�?���~���d�ҙ�d
�B�����XU]?r�4����\f&�HgG�+�
�P�̆�X�� A@Ehgfhg>������ ��$���pA~�p��3�7i �J��zk[Az!E!��j�y����҃����A����	eG�B����fv.�V�A���>~��dUS2*)9���jZr=��WHU��s�Bj[^V@�$(����$�o��/�'��I�N7��K^�G��EGE�(
���m�
��V���������f��ֶ�$�pqwu�9f��ӷ���Ja�%�{(�W�l%Y� ����*U�r��;�hG֮��� ?�D��<Z7��]���V[@To��������Q�˱k�$�y�J;?���Ǒ
9Ė���'%%���,^:�¥c7�/�� ��0�G�'������n���9���=f����,Y{����������6&�+�+�kqz�C(Rh�|Nw���(_�F��%͐B��^������]���������ƎB`K$��nb��h����Կ�n� h77w��ٮ��.�X?���[��K���ZZY���T�֎����<�haڱ���D��ϟ�B^m���<?������i�jOF�S�d�L�
����@�|�u|���gu�㴿ᶿ�h^�կؚ]���,�{��-t���-]�uU�?4I[�[��5��%����
'h��o�N�:r�O�P�w������C����044d�`sSSkK;[�����̅�y��y�� �%�}aE-������酙�p�Ơ� hz?_W��F(����۾q��G������rs��p�GE{��?6.<��gݼ;V�>�x����ܺ�,=W����A���75�uu������������������� �F��-�����������/_<�~�2P�l�mL��m,��Z���YC"xX����}���q��^�� �n�(�����K�A��c����)�8���LMD�a=���L�D�kɗ�ݟ<uђ�GO�2j�̑�f3u��)CGM�=-n�̘13&�^�f��GYU���;OKK���ħ夬:F	YRNU�KH��~J	���*'����(ѧ�(�"	AtKU����z�LF��2t䄑�M�6w��y��&��	��
�7)8zL��	����x���xbWNI�&�ډbQ( B���:��.��\I��(W��!�Y��t�e�^q:�>� 5�o�w�.�[{�T2�A�Q�A�U��sdz���O/,LON�}�Жu��]��ȱ}k�.s���� �hw8~C+�#�`_w��
�@�{��oV��Pg���^�|��㤽�v�;:9�����mjm�3Ym]�tM(U��P�Q=��
hM��3� �(z@�[�z	��ʻX���l�=tE7C�"x 줩��)h���=�������m��عy!�PweP��=u;� ������z����Z���E-����<n�L���Rq�I��\���B�Z��3� ��kw��\v�����U��c�����Q���=C�J��i)�տ0:����>��>�P����T��T����R����ߠ}�U���wAH�_m �AHmIm��Ed~��{/ܾ�8�ȥ;1c<�#�m��-��@��g�6�`��#++ aph8xQ�^��_\QP\RX�P����^��evq��cã¡u��������⼌�o��\��a��XwOW{wx��s0���3yL�̉qS���G��BJ�*T���c����� ����RY���&uW�/��t������_5:���"�o ��y�ɩ&����nH<�^&�W��l,�B��Y��Y��ٚ�/lL�=�wC��m�R�n��0,�f�����:�M��6N��NW�0���i�������V�'W5CB�FA]�O+���Z�#�M|��𙥫�L��@ሱ3���>l�4�`��Q#�E��>kѦ�/>z^��S�YҘ[ٚSޒ]֜WE(�&דKq��Vv]+���o 񚨢f���!ke)	l��!�T �������`��-G.O_�mӡ��^�|�ʶc�w�����Sw���w;��ܭ�M{�҅���V����,ѐ�"�\)(����J�<�@����НB��V�c���9v�a�d¶���K#M�t�Y��E���xKcJ*�k�+�AE�T�+*r��Z������ʍsU�%��w��x;�fquu�s����4����tttb����\}d�7���O�5�߰/��g��GTT����f>�x�k�΄�	OR���糸���ʪD2��r(�nL�D�Y7,�C���C�g_�}���#��S���=��Lw
Z��� �m�[?wk�5���Y�;�����)�,�	��h��iَg��>}�_���?'��?yvw���
�O$�8go�,���<�}���r�;ftl�=+�Ή=[7�XN!q�Զ���<��'UmY�WE�w�x�M�y��l�Vp�	�߳[��di�_�k?�_i�/��ڻ��:��ڬ&��������O�������:���N{)�X�j���K�������#7��<y#x�$lX�5���p�@C����Pׇ���> (��aAIeQY�r\�N���ZRu5�0Ojn6l�d� ?_?4��A�(g��P:_>}T����;qdT�?�	���V�� ���"�\���#V�}��W�f�fmd����8'������{i�(R�Ɩfe���?;��l��w����h��d��C
�s��CkKsp�*.̯�(}�p@�2��t�1s���9��m���Bݜ�&���{�B����͛ꏆíìb=�N�!D�~ZDȯ��� ��FReD?�X�J���-���B��7v��qP�.ۺ��դ���9�Y�UMŵ��BY��� �Om#����o�5�қ	�V2�@��
SLeI(9�#�� T���W��5���~�G����o9yž+;/>�}���ˏ�\I�=�������:q+�I!�VJ��Ug�TD���3E��"m�r�=P	�Bi�ST��l�.�P�⣤���5��TJ��]�wk��_��o�}TIS�"��"�����x��'��*��*j���:������)	1C#�с������������������O\}�?@�B�##���ȉ���ٻk��M3�� >NN.,.bqxT:�Dadd灊���*�)Eo�[=���n}~�P	=ȓvB�n�Qt1�t`j?��6��hf�恄}Qz�� !����l�7b�w/'T߼?5-��2�������k�\̘w�I� L��\�n��E.]�7z��sf͜��N�zbߪ�+2YK��9cKJļ�!sN�)��-?�Sis�/��V����ک=� ��Xż����
-�G�P��sԩ�I�J�v��ăI8ːs<�����ĭk����:�4z㥱�-=�P�}��l��k\Z���g�p��X{�������a/�ߚ�����]@@�= AE�W+k��U���|3�P !x���)aH�'8o��r�͟6a���K�L����/��R'�
��M���Ve�#bu���@�;
@��(���ZTΨo}�P@����E��'�?ۏ��c��O���)8
ز�L��G�m�MlL�N�'�޵s�¹������f������րC`����ȡa�/��r�Hd��;��b�������������
�Z@̫a70J(�8b9��O �4A�-P���t?���Cg���d�����L��0{�S殚<g��-�^KL|Z�4�<���������ka�[���&
���o"7�PZZ� D�L�zZSKDcK�\)�/�qe:-U���Q�:q�����^,|B`�0x��K�@����� C�q&��×;��}&����x���A����d(d4����x͔�bJ_�;>��kOS}��,b�.��۷�(>��;aSf����H�N$�)�f�R��R�K��˳�$][�a��+�>�߼m� wrځ�삢f���@A777�G������[��5?��C~x�� �������|HTlę󧞤>:u����<Jx���_\�����Hedd ��ˡ��!�~��!�U�%�P�
���Y� Au���*��B�~����"<|��B�B����p�@�c������`[?���H������] 
�	/��|t�ٳ7�iO'�go_��x���W-{��p��U۶oY�`Vx 2;�����6���`��N=�L~��}Վ\�B�.zI�B{�H��بMW�_���}�����&����v�y��߁�O��N��]���w��k��Z�[m�w�ɴ���R�T��;�VH~�qª��\\��:4�BSc#�!���E_�e������?��z��F��Մ�JV�����C�F�8Z����l��� �F@>P�;�� =]�=\��ζ('[Ӂ�����L��b΄?�@oo/���Gyz�p��aA@��I4f�U�����g�����n"!���'��$����C� �M��M?��ikmnmnde2��x���!�@���l��x��� c��؂������G���c&͞2{��5ۗ�۽d�=�.�J�H�,y�W�Y\�_ހ#0	̦V&����xR	D:��&Q������b_�*��
d��I$k+pbM����ԓP,9���݊��K��/<� �DR��Ǖ�k�<��������nP=,d��^�M�O,��(yK����deE���|K��E�?C��5#װ��,e]�#{��d�5�b��bΧ�N�E�������X�I�QitBG�D�Bӵ6U��K7�_���Jjz��
D ���D"ݜ��A���Xl@@ �����-W����~�A��Ó�B_Oo]0^ °=��?�y�W������a�ÔT !���C��] ~o�%�?V��!��;�25E�d�u�U=��_�䓦nO�����.�K�������MG T�/8����/p��C����5�M��'�tx��}o\�QѲ�t|� �v'~Ҕ)�qq�v�X�l銕�F��3�����K֬YH�H\�^v����;H��KjP�\�|6sց���{�f*�hѓ���S��L�T7iO�6t�Ø�i��r�N;�����u�N�km�m�B����N̬C�s���;��|v�T�=���w���q�k`$6,�� �[��;@�`v�֖��SS���Lwi�[�Y��"�[X^�R^��x�27��^辊@��p`5�|��x ������J�>��|	�tu��674p�1
�v�p6��jo�'p��T�B���X\V_�&�'3h:Yx�G����!�.��䩅�����5 ����Č�dj4 �����
|B����ښ���Iژ@
``o5�h�� �uvq��AX؜W�(n��4��V5@��D a}����OƵ��*q�i����ٸe��5[�-Z5}��	S���f.��`-���xP>+�I+��*���������zr5��c�q�wu�Ă�E"�Å'�5�ť,N�P���Q)�՚,�E�����Ie׵4扄ړ��A}v?�����kW�pgU�/���A=���I����	X���6�?��~#�>��>U��Aq����(�J{��>yR��!8�@iwBK�ɻh��;�ݜF��e)u�|��I�.M\u�~������6*���R��ML�7���
_y�޵�������&�'g�;�D��!��.2�>޾Xh�__��@�s���������A�����Fy���[��hfb���w�?~������Db��4����P��Pګ��s�.�d�НBuz��N���/�;�}2�
�DJ�k�o���2�!s���<w�C#��<��|L��tvw�O�+�@�������#Ay�䂶CFN^|`á�D�P�E�S�Oq�����n�Nxp:�`����/�񍩙�KW���:f܄�G�m޼uc��4��_�t 2&��|����q�6��-8�O!| �h��,�|�3~s�Z��h���(�����S/9w�\>�x����
{S���38��^'|Ҋ��|�6|���\�ܣ�F,h"��>;G̛����͇�mك
���G8��Z9��]�ݐp��3������eή�H77���pw��� �K�A
J�����7���2R�v�Q�ac���A���� o !4��!����@{sh8������N`���Q7���;���Q7Ѩ������������<�����_��Z\F������qM��V��gKxB�D%���/�i�~���{�u�	�j!�@�O��҄g��60dla����!P��p���@ ao!�!�����-�02�2�ͯ6������	B�@pX]�RXZ��Yx���c'/�=pbˎ��n]�l(AFO���gi�u  ��r|N>�����PZG�h�T[� �,��@����x
(�آ=Wn{��9nþ����?}�^�L����-� ��":f+<p	:j��w/%��|Z�T�<l�d�L3t��Ǩ�kN&3���7�_~�-jaܼ��֟�p'E�G|y���`���
h��B(U3emz�n^�[����$Z���մ�:�'R�6��=y婄�V��38P�$J�����*�T�)���-o�J�M�*�7y<P������������Po!H��.� ����#x��^������D��ۚ[G%&'d�647	�2�D~RO
,"B�4I�L� ߄)���V�F�;ڋ��S�-��b�Ð�1�Mڵ~cc�d�B�y{��|����Hdt�0_l������o߾ms�s�ָ��Y����O<U�D�	�}
�O�	q")��)D�����Ƥ��sWn��x�Z|���o�NJy���W����������2��Xb��dZM������SK���,`��X1r�ɦvmR���#�ס�����
ɒs�q�<l�{<�HZ��Cj;��o�aˏ�ui[�i��	Fm���jgxX�іr�3��(¦n����͇m��44��������E{x����@��;'84�� �-(�-��/��[RR�/-���J���1�|���|��|"B}�0nN���MA�"ĺ>�>A<� ��B��� ��@����=��;6�any��N�~�	��������!Od�+B`!�6QEw��Z;�Y������6�FC�X�A7AE����ξWAP��<`!8�33����3�Vbrvs�q�RДSC-����e-��V ��(���1��*#�(!����K�o:|�����6k��	3bGM�>1j�d=���� ,j �(m|^��)oɭl-�!ד�ixzu+����%���j������ǯ�5r���wjvޮ�$�^S��-h恨�'7��[�7�+r�K�+�r�x���񈝻���cw����������pO>�w-=l��%�ɿ�R��(��~����'-M-#�4�ɂ�;�d7���mZ�Z;uŉ>�_�rtM�d26_�'�h-Tb}Kc~Y��qc����?��6��~��cE�������pA�Z�YY���^����d
���蒨:@���~�����y��!�UZ�Jw����}��:BJ�$����$(�I���y�nݺ}ĺ�J���s�:|�ꥅ��7�6ggg��P�Y�=t�d~a���7�-Z�f���_|��K�'d<u]�}g��8�Z�Y)k}���~�va�z��9��գ�.�}�j����w����~����_j�/;���k�6vi���.m���E�.$��Z�F;t���e�R��|��"�Rv��z�v�匭7�G�=��~Q&~�0t6,v�M��	[�Ǘ��D�ėp�f���m�բZ�gT�ܹ�/�ql���Q��ё�!������!>�^Aؠ ��� (A� �aQh/��WAE�ST	�[\��������R�/w����a���b�ㆆF������K|�fj� �������vV�	.0ݲ�Vw;/�+�0*zLVN]u����xaS���m%�[��
���?���g�S����o�hx�k���(�if�ƌ64�A��l�Y%,M�M�Y��!
�-��.�6�B !�@�dos4� tq�t�t�K.jά �Q�����CX�H5a:60��nH���a؀P$��
�522nR���Kpz�*Zr*[�kI@�R<���Y���&�@�H�J2�,�(l�K�pwj%GKh�J`�Ͽ��q��2tۃBi�]~Cۥ5�A�&�ߗ��b`�s">;����(�V7w�Y�����bb{����'מxT��P�{{<����
��r֋	����r�,}�����C��AȔC�d/�%�wsv^LN�嗒_�?'M[q"1��-�̔v	U��KP*�D��H�\9�+J�4���r��Q��n�Hwol��3���tZ��'��o��S���.X/]�^�7��=���:$jx'PY"�U���h�E�.��w"h�X�'�-VA�O�
B}��,��"Dr�PM��f^�R��Ӯ\��,/��(e���)����=p�DmS�ӴgC�+*,����$�~£KW�>y.���WM���&}��ʃ,��	g�==}�鉛Oǧq?k	=�g4	�+h�KH���*F{����QAՔ��L�o	i5�V�U��-���f�PBn�V�R[�h�!+��d�	�=Zb��^�1��ѡ��I>����8����N�F�Ֆ�J��-B�Km��9����"�V��4���ŋ�_��Ժ�}"#�C��~A���~a~�a�aAa!���P"�A�����
���j��  ¢bJF*�tP�3;��`��h=��!X$+���p�6A¬A ~z�]�G:���;��n6(���&M�WZF��I�K���'�?������~��B�S�$�B���B]fD�aE�z�!7L��������������C3���"��6��5�k�C	A�E��6������@;��6�C�mL�mmX8���>)hzVJ���]��(X�H G=�1�;"ж��0$8����|�`� (�~!�n~�AQ��L_�f熝� ��2�eU �sk3J�r*��Մ�"@��Ê$"�����t�%�W	{t��ٛ�&��>pWTH�Nٔ7z��RO9�#�A���\���OԲ����S<̣�Ӂ��>7r�J�#�����F->������Jλ����n�L�������p+A��!_����1�h�Pga7U�Mu�/I�����V�>i�W��s��Li�I~����y{�P&Pw��{�2��'�e<�R,V_ō��CǏE��1: 8������z�E�������vwC��c�]\�4,����+=A\�n��08('�����H$*$$,$$�D����Dyy���g�� o?O�54,�b����N�`���+(�o��~�  ���('����[w����n���D�X��E����s�"2�r(��*�V��.��*��.=��Q�6�P?���`�],k�%W&e�dT��E�N�����F����˗�$��>{te����܌�ϒ�O�Y����6v�Ĵ��PrA�ݺ �lfR�/��W��/�]��申ي?d���ү�4��]��j��{{nF�?��쳖�=�W�N�]v�B�ە����1���~���C�D���G�N���W���=[񞫁g(?�'P՟���ͯPھP�>Q�>@iE�O�����/�i�;�$��Z<�U��E�w��y���C�}#@9���������-M���@�J*s*�׀�+2|I	�q"�p��&����	n Q@����
�ø�:�r��t  P��n�Fc�������F��4|�w[���7"]�ݑ�^� �E�6d�4d��kk���W��cn�����72�x2O!�(th�W�̯��Wm8<k�����ap������3#c3�!Ɔд2V&6�F?����޲7����,XB�40`0�|=�� |�����j���E[�CX�'�U2�!�-F���s�p�	�3e����Wn�r�̥�)����>ή�,o
�mn)��R��(mdU5DaERG�3��LyK��w�%=��s	�2{Cn��D���C�=�[�������7�~-&��j�%M꥛o�D�Z������畲2B{^��i�V:�����Vج�a�� <� ��r�A��%��UZP��5j�6���_ �.�����~���������ܪ����)l䧔P�j�%��b���y�u�J��L��+MȘ�6	O�gKE"�L��RY�ǩ)3��>z\pX\P��������Bc�#����>��N�CB�|}}��@�ᑑ�9pb���A!~~~�F�
�"266�w�F���zy{ ���(�酌��@��0�qq1�U#�`�����>r�04��O�<�?�;{�\� ����qq�z3%�qQ`�8|�D(�tB���,i{������Εw��E�E��b���BP���UV�\�Q�xm]T�����k/z�};��4�R*d�ߟ�pBfyAbNvysCYc;c��F+��B���o9z��i��m�/Z~��d�;@ G�m��_��T��7�N�[�������3www"$$$���@C���[�d��.�0s�3��}w���J����4�Hׯ�]���ߝ��U+��o��;=��Q��4�G�%'�������W_I��%:�n��dJo��E�������*�kY����h֊����,9��C�>X�wL�[��NSg�u7����>��al�G�䝸±[��^����3W�t=@�?�/0�'p�8��.�bDܒPs4
��\�=�yE�0�����,�&�jd0j���f�fz�B�ㄉ�PdJ24����:`�,�77(Z��7�11 ��f� �({{�� ?�O�eˡܼ��|j~!�'�?!�GҀ	���W��(!K%�R��BP�c�9%��;���{nێ���^�PN_G�����XOnRo�kj��	|5�@@!�����P��������0�a(�!�~LC �C<�&;��x��I���V�Af�]le�bfngni������?A<<�K������Ξ���X�n����}FY��Lι�2!<>?� ����a�հ���XN)^XFU�%UIDV�h�K����~9��H�1Z�R&d5���4��=�36��!�r��rzL6y�c��w�R�������:UA�2*����K��5�����3c��_V�?�UГb���U�Oe����6�I���C�������(�+�M�5������^�\~����
R��;�u�~c���q(L1�(�-ȸ�&W&�I�pQ(�p������=x�4�q(�������p`���10i����6����u+�̍M�[�n����u�ݼ�W�����ͮ=����������lm���?hffaff��~##]�a�vo1�0�<�m���ls��4��������g�����;~Ⰵ�x'N��󶰵Di���L�����'�%������R�A�G�����㝪��փ�4��_!�{z �\[4W�7#��6A�R�BBPCH�i�v���1e˔�7�DS�p��XY�����J
1�S� 6��J�I�<{G,f���ȟF%����M*ډ�֜ޞ3���s�s���<�Ȳ}�����7O��p���;B˰�P�
Z|.��kQ��A�����,9 �DU�D��)�re�B�,W�Ȕm2E�T�)Vt��+o�/Qv2���j�&|����oj (��[����j�8k͑�w��yz����cǻ�x�cNO/'p|�\���Gs^9 (�ܾ��O�W.iZk(,��$�l��-]�+8�A u!���6ӷ77r�0v�F#ݗ�-�A-��������j��w%�4�7��P@�hg�C��� ��nh�'�?�?m!�ZG!h $AQXQ��.�o�z�ة�6�rq�!�9Sc3#�7301�11��th#-Sá�������P ��������>���!����^c�,q���Z��ah ��W
�q%�4aE-@jA�������B @@bfi�kln��4f���K�N[�<��}̛�򽧯-\����Gێ���ȕ�/m�{n��3 �v�߸�Ҧ�9|����^xZFk�(���|a���E䏕L�a"�y��7��yJ���S���J����.3�<���tM�=s��GqP��l�,�v���R���v��trǥ��^f;W�v�����Q+y;y���/Rq����h�,̮c<��|����{aɩ��#�w���/�|���!��T�P/��>~n���*0u� ?���yR1�Oa�@ix�N�I�ͬ�Q(�1c�_�~���t��1{�m�/�����3kZ}]�������8\��&M���1]�~ݺ�H!�;rɒE���!!!3g�d��K5����ƍk�Z��'�

E�%K�m����\�|��d邝�����ܮ߰Z(�.Z�`�Eu57�?e�_���᳜�&�^�mܔ�Sgo`��;z!U���M�#�AлϿ�>}~"� ��'Sk8�!����S�_!lE JU|!_��m�iwn9�t��7U䏩����b��q��R�%Yuu�DB^eUIM]��ObaH�j�$���P��rļ��$����q����)����C�?��!j4zͭ�/�'s��{\�D��� �wh٥��ת"�4�J�ƭ�Bi�@�U*�*�\�Q4���F���f��K�j�|%��U�@x�����N��D��(�
���Ne�W�q�ԥ��޾v�م�F��������`�`m�l������
z7/x)~w�" ���/�0;�(�#�3����4��ݬ-[�L�6������������������>��d��b�����:.�oڸ�&��1a$[S}K}[w��Y�6�HϬ�- ��d������1��G~�#�בIX
Yj�U����8tiҤ��(�0}]+sks������܌� &��P��X��d��������!��`����������	m�dj�hfdo���sW;xN�L�J-!"�U��6�������s�[�����̭ll�]�\\�]�m����h3#��������n�?�K���_������ح�Gn�9�hϹ����ȵ��o��������swc�ݍ<?���W�go)'��%W��>f��_\Gou�}��W��e��'B�<'���g�2�	+@)�4�6�B�^&p��u�Rב�A�]|�PUBQ�	�A=���5�^;��jN�����/��lۨ�p�V��9h��A�n]S��r�?����,:�4�ޝ[/��8y���YK�K{�E��o�Mo�$�T���U��{oIY֭{�"�^*��"![�c
9TK&���rƅK�gϾ�|����Q��9s��楒�5����N���Ǎ�w����~Y��UOȜ8eLBr�EZ�r��'�d�ys"#_r8��+�=z
H[�~ս�����+�ܽF��׮[�:�9�G[�f���P���ܺ}M&m޲������m'����C_�aM���Ș���ʬ<\~)������b.�K�Ұ�����@n���|�'Q��n��
{��}  �ۓ����w<��G�������5T�d�����F�nr�kj�6wRU]����V�!�X�w|q'�S��3E�Y'l.$r:~��-�>BP�g��ݨ��=C���Tw$
ɻ���>}��+�<��DbE3�_r����ae����%�:t9���LRh�x�W%Rh���[oկ����ԜC�B](�t`؍L��-s��Z��A@��p�ᬲ�I��B�3�-Ҧ6��IaE�._E�5�]��O͝PS�o��o�ʖ�����O�.>n��swn��|#t��)>�Ya=C]�����%���A�������@��p��㴬���2�Kkr�j�*`s�%��3v�9=e�_?׀ ��@_/'�X��3PpT���@����G���چ��L�?k�ȹ��Μ8b�`�Ȩ �@O���!�Vý�],t������^��MB~i3��6B"���5H�/�B�s��6B�!� � �mk�ҫ�䌜��Vx���9Z�̜�,�mжVƖhms�ah��`x&�6h-[�P[4��ek�r��r�Ҷ5յC��[��Z����,u,�L�-���fL:�Er<���!��_Y_TU,,�ԃ ͬlu��t��w��fV��ր@-��Zz��h]cS;w�ѓg��zp���v�֗���؜ZN%����.'�J�"�2��	REVUQd�4a5M:q��jr���Kx�E�̢Gfr^fq�)o�9����e����g��A��ʈ���&����K��'�^V�h!I�㥽n��캗95u�f�j2=Q��/��s ��F`͆��Wp0�H�!l�~:�@x�ҙ�ۖ�����w�Ji�nDd��6�(jTpۚ�-�ҜܴWQ��A��ri<:���������e~'/�PV^S��Z�b^F֛���5kS��|e���9�IJ����)o�R�̹���(��6�LJ�es�;vnIMM��Y��{�&Z,��ڽ-1)�/`:�/:���:v�PZz��}�w%%��}���Q@�m�~}��B!9w�t\B�T!ڽowNAaie}A)���QU�!2�L	�&"4�*kH%E�5�:�T��뷞��ʦV
�]U[_RQ�B��j��_@[�BM�F����lb�Z�����1��+��I�,iw�G(��U@�wBx��g	u���['��W��,�J�C4�op���f���A�U�>v7����c���~1���^����B	�S�ʡ~����W��N���+l�rT%�|��������wA��^~s���CԬ�4��{��o��}E[���E�թ��5�����w�=_��_mm�[�B]��>��R�A����6��h�#n����&,8u1��W�o?=qF@�8s��Zô�����@����Ѧ��VV6  B��  arZ��B�WF�ʑ���ذi��1#��<��]���\�,M&��9q�p���`�,��:~����A�Ƈh 7�k��˄���N腓�n]5�����l�̅ᯒ�0̢rV9�'�?���y���GF��?�\O��&�;�9�:X{x:-Z<}��I��N.&N�:�(s����x���@AB�!�����/�^{�Ī����C���\-�\�� �����/�Z�VD}�Z�A���Uu0��ºY��YYk���!�	xS�򦎡��������I3�l>4o�s��n��^�W�%f'���ɊJ���",�pK��b
���o���0�IUPE�����������tU��+�� v_�c9�,Z�l�awԲZ@j�M �2���(��4bMzH��������ZAp�f���%���mzG6�*QG]�������~�|] �s���mn�x���2ڎ�$�'���)�2�
������@������S�OfP�b6�G�3�d�KP�ַUU�K�8yEyi��LHzUQU�}ۦĸץ��@���C�2V�Y������E+�?y񰲮lۮ_��?��N^�aŝ��Sғ,�{�ލ̜���fFD�g�e�ߴ��;�9;��z'�(gպO�=*./\�jɳ�0��SgN������/��\|���EK��%&��?>OѸ
�@H�S�5Մ�bLvay�\%m�lk���e4���2#3�ʍ�D���G�_� �\��!G_��X�>C8h�(����+o�(Z�������������V�h�A����#t�i������s�u�c2���E]�O7�U���Խ���z�@XL�:�����{��31�Z��Jh]X�p���}/漥�A��N�����"� �
�BxDi��"����(�DQ��)��-}��^����iL?UYI�H4q�}��/��O�ބ���\�W��Q�,|G} �7�ފ[!q$m�����B
��� 3e�ѳ��܍8w�a�ؙ~���,ᗛj𦣥m��gl���6��Y嵹������l�����W�y�@��n�lgj�����鄜�7'� 堏���p?g`! p s��
��D(O�&+��˦������u�y~��-�pj��?!����m0�O_G<��BM�z
�D'�{tW[����S��R��\|}������P��PSj 4G�B�A����v�t'g����������#���km>�����u�G���ZQv-��<����:\�dּ�0�z� B�R��1�������ȉ�W�zp��������De�<�I�X�PHL�f�c(���,��@/"��h�2��s�4%�!��eSʭT�x^+���|5��>8������Vs3+���is04U-C E'HE�-#�K��
������IAp�F���*n�qTd��.m�qeLE3��n���?@HQ���}8Q|�i��;g��;st�����i�nƒ�_��"9�Ψ���d�55�2�JVbZjF^�\O0]����5���	�*0�Լ�褨��6E�	/.��`���G.�i���g�#;����U��r��;o���=�+9=��8��Ƀ�_>��Nݸy=�/� k�����eŇ��y]X\|����ȈҊ��w'��Wb�w����[8<r��ݕ�V�%����n)��09":GFcKi<	���3�դ
�`Ni
�����ΞN<�PQU���������L�E
5W�`������p���C�X�w��9�6B���*��4���<�:��������T�썷����_���O��NAI��-ܐh�{�,��A����`��4(;�N���>P�-m�<o��u@�/(+k�=M�C��?�1բwI����[!nt�^��(��i�����>^�(�h�'s=I��Л	K�T0��K �Y�}L(eߏ�T~�0��'IuGo�o;�����,��L
���H�t�e~B�Mn�u�N�;'�ĕ#&���ofᬥc ��گ��a0��:�FF�&����B aJz� �酕%��2lN	5#W��:��yvn�>A������>���G��x�T6��TW�|�4@ Ҁ���fT��Q�����~�Bݪ%�Gۙ;ػ��r?��RT�-��	���l4�h O_�j �nkz0!R���w��M�W�����F�'T�&��i9X�l�(K4��ei<Q��D��T��eg��qy�JZT[�|�hs'K���PS=']'c}{cS������8��e����znI���^��������H�=�������1���HPC��]mCCkgא	�Vm:4k�>��N���/��
p�qe�Ղ�jvd.&���S�,��K)�� WEW!NYp8�XZC*�Xʿ�k�c5�2UH04E5U^E������"��(@4��Hk�����2$�����Jx�[ڄ�78�!��r���}����5��87m���y��Y���b���G�ʉ���Ņ�2����W�RW��I��-��ʹT!����J�Z���Hµ�ia��$f'nۻ�E��k�/�ݻ3)!��3 ��/^=��qvaڡ{�E����/�*,�}�*,� `v��͌��JL��K�SS��ro޹�����z�����r����Sv;�ViuINQ���2�2��?����_Z�{�>*�ŗ��\	�'��P�T煽�O�djaw__(���e��'$%��xEӛW���D	(V���@E8d�L��\���_>�U��9&��oj�^��/����j���'/ߊu6�\��x�5����X��e�[e/�rg��J�IW	RPB8U��3�A���Z/�%�+��}�p��#m�+��	:��P��A�Mj�oOk������(}	{ ��G/9��Hܴ�^ӎ=�R�=�X�Y%�ܦ�񜹿���r���U��uʮ��VK �G(���a�/*Yo��a� �6_[y���;��v��_�?������ޱ����Ia�5��o#�n�p��K���2i�������>Z[Wy�������M���h����_`Ѓ�O�f�W Ӌ�@2K�2�)y%��v�GO��������������hma8qL�?P޽z.���]���v��s��; Ep_�Ź�F���5�/�ѵ؇��X�%��������N�.��W�~B����w�d2�v��mm�a&h�)�G�e'ЈU7.�5bi���DY��Ԃ޻0�֮}�g����([#�������������5e��w����<)��S�*�2J��2,�;�@�jpD !�� �Ǣ��ii��@<~��Mg.�ol=��gU\>.�^�?p)f�櫩��:yt�YJ��=7���:�\Nju!M1q��"9a=[\�j"��#�DH�!|��
8����Ða�Z���#'�$��.nA D�]�	��ˮ���'����zp�Ǝ#g���i[/��QT}�,)�ɧ0�4��dUWV5�խ46���$)7)�0��V�[�R8�S9�s��w��Ӣ��SW�^�u��GO�B�2Rnߺ���T^U�����h ���G
�s������'��Iu���u5)�)��>������|��y-��c����6�+k��޾Z����k>n+�N\8�_����v�܉���~9BP�٢����܍s�y��u��b�L �k9y@��{�38���.�)0�28�o�B��gT���"�! i�.���QB�u��:n+����#��y�n��<h֚�/��gC<ǟ\ ��e��eX�wf�g�B�y�[̒NXy������P.Y=j�֜Q�#l�*��Jo{Gj�6�S�Zi- ͚���$$Շ1+�>Al���дu/�^���ADIw�q��o���d���˩4�m��y��Y���z�ϲKW�8�hƞ��7�eg��5�wB�2���uW�<�����}6�,�N�MQg�ec�l_���γ��<<a���h��Ο^��Æ���ŉ��aZAEZQ%HFImF�����j��\|�=\}�� ��NV���#������͍����с���@ !p����@7W#7+�q>����'�/�6a����+an9=��YZ��	���o�	B2��,���[�B���LL]��G�����3�Bi�ja4ԂV�:�f��f[S][3m[�a�L4�GY�LQ�(�a(�С���,�������-MamF9z̏JoH)&�k�T��U`�*k+k���J�kA�.Z*B}CCc�Ԍ�"���j�]K'��q��m<0c�>#���+SJiU��<��%'�\�����@��o��N-��|Ɏ'A3��ר�)M��?C(òX�G�}�)�D����`�R89��  A��t� ! ��-'�� B�H2P� ���`��r����a��/^ݾk��+�/�{��WL�r���]�oe+�)&2��BOPZ\��SP�j�Ց�UE���KjHBy=�-)���|Ѻ��v|N��K��"B3s��ß>~� ��8@�URU�U�y���j\%���z�]��(���Ҳ�c������zO��Y<~JFv�R���|�V�#�D��".�V��.�4VT_�y�S�_R ��x�4O
 $�U8½g�|��ce-b�R�%ԧ�d��zu��%������
�� T��y�.���(laR	~��M�c�������M�Bx��9NGf�-��lʕ�J��U'�g�K�s:�pry�H�l�p�q�ߌ��]�+_~�ʼ�kM��>�,C�Fnl%7�R��iMjF��Ѫ`�J��J6���1n��G�ŕv��0v���hӹ���)���3�߭��|%�e���"�������#��"h���	��O%���_P�A�K�xUS��Φ��;���
^�����[�x�Z"�q��l�s;�=X��t�ą�#�,]t�t�ttt� :Z��E��t����>�>~�O��g�疀�啧旧��cC�����C���l�lg�=3Cd�QcwsOG�x����Te<e6�rڨ��6!�>.�~Ϣ2�+���?!�	�?���$8`z��#-]csK[j�j������1ZO�TW�LO��P��D�
^�A����<w��x���0[�������P �J��o6T�B[�m�oib�2+"�:>�V��(�d�V��U�WVT��Y�mi�g�ob�6��Dbfa�635B����t���L,]��M]��д���f���L�`�5_��lV/��<pօ̆�ϲ[�����|J��d���˚rB#(���MS��.Q$��?C���~���Z�~��Z�5%�aC���y
�P2 !���@/_;_>!k�4}d�CO򩯋	|)�]O���-����rA��}���n�g�qLP
�q$
�VV^��٫g�^W7���ꒋ��fV���^oJm��U�^��q��b^ �^�D��?+�(RVY\RU�U���)ɺ����@�QC�C��5��o�+J��r�L��%Wo�{����:6K��a�/޸*{P�=~���e1������[O#�xx��/�T�xp�[����|!i.��ܢjLD\tbvr|z��x*>�(p{��5�+�AEXK �B���M�]\����@crf��u��m��|���$�7�~�W��xG�|_�Um�����TE���/jd(?����\ֹ��B�`孌��wlIU�&���@AZ��Ѣ�@(��}�w�g���Щ��7����TŁ��M�����y�㥑5߇�6�DNhهb���͂^���	6>�[~�t�3ܝҶygSp� ߍ�մ��C�ߡ;��i�"�;���<ɷH��j�Z|�3wӢ]g7���r�I�13m=�[9�[���������X��-�ͬ,��Ѧ�46B}���F��� �������nژ����|�\�<�=\�-�<��zC@Q�di�s�1q�5u�3C�Ј��F����,�PN�a����v�1��^��i��
6����_��	���?n�0����!ܡ�Kd\�v@_�glnjdn��7 1��A���Y�Y�ľ�MA�}@������)�X�2D����C� ���Z��!hSC3�`+��q9��e��e59e�`A���T�& B�"��Z����������mef`n�o����t�����[N��^�RƎ/��?��T�z�ް��K�,���X����ao��&���,h���$8h%q�)�����)��`|,]���&��I�t)��@T�ѕ�2p4�#PǕ�r
OAh"��!�ݿ6&�R��`)�
<�C�Δw��p�U�O����Wς׃�k�
y�ʄ}���i��������r\-��'��*^�NX�b��瑵$rY�add|~1��(l��X���~{)��S���z�γ��e�`!LEiU0���
��-�w��� @��Z@bYIe9�����Ĵ��rLznQRFnvqUN	|d�_U�S^u��3
_����eB"�D��>z�B5_Q��(,���+�`qDR�HN�KA(1C(*�Tde��o�S�w���M[�*�Z9�4+���#פ����u8ʦ�p5Sc��&d	od6�fN)W���wP�m,e/���a+{�wLi�QMW�)m
z����LiS3�۹�]LE���S[����IR@��JY������k{'l�Ȼ����f�ۙM ���f8�NS;]�&��:u���wb8��b�B�V��y�>�1�d��A�n9�9W �
����<�c�M�U7n��I<O_q#�\�����
Eq����z��4�4��GE�OP�cĚ�5��<f��/ǯ���)x��W������3ܺ����������[��� �����A�>K��K�.N�)N�+��Eխ6�s�Lspw
�	�	����h�Ad�5[Sx����%����?��6�l�ZxZ��8�N娫���������y���
+��qpD�D�i�������`a�N����O���O ,���u��	����@hb���F�z:��zڦ:�v& ��h8f���Vv�h3==�!���p���fhT��U���̗�Uor�*p�uy���:4jln ���r�pu�p��u����3�],��̬�\�,ܫg5��{Er)'2�<w�y�Z��{���x}%���\!	�w*2�SEj�K�q��KNU�P�=TAkC���/�@�#u4�K�0�X�j �L%�.9RGF��A�B8�B�z(�vDA���A�V�h,�t.�u}��N=Y��8������s������=�H�/�~=���ű�W�?"�ʭ�����x�����W���&�0�_�Wr��Fg�n=z�5TV�Z����Ƞz�4����������HmfaW* �,��| |�D,��P]�/(��K�n�H怽�뤬j�ʗ�b��x�+�#��)�\e��!�g���r�jt�(��	] u$�Em��E�뽇�xB�t`�r8��BG��V� �
�G@�(Tu���U5s��ؽ���rO������j�੻XҷT�{
�w��t@���#D}��������z$
8%��[�	/
s�,
��(i%�Z&.>�m��i��j���aD���rq�/�+E�UH�yM�|��rx�[L�Y ����u_x���r#�dT��_��� |��Ȕ�7f�;iǍ|��X|�ĭ�6^�������Bf74r�k���z���#g\�G���s�rr�����{����J��|~�-	�}���=��MV����Y�[���5&�^V������~�`B8��̨B[� {s ���G������ ¢������6°W�@�*���Yn��i �))�ON� �-4156660��7���f�?��`����9Z����������������������*B=P,4���k��i��F��̬a_h �\G��|au]1[^g��ehK+Cc;[ ���������W�� `�'<��h�7��p�0C�~��
�>M�r���l���5�G����´��3�\�2akr���ف�K3�/S��DN�����i�iBj�ׄ��Ejޫ�KpL%�)�D
����
� �h d�A�%��3�Xn3N��qF��%{�?A4V��]g"�0�_�|��4�\.x�I���m�p��z����sd\��ʒ`��Ԝ�������*2�W��m��^N�;PJ�>)��H[�$��Be+O�b
�t����иl8<&M��ʅʎfeG+O*��Y���{�\8>W���ژ|�''�E�ע�:1$O��#��AtQGc�wU׷�ߠ��� �"e-�Cf�HL6��)�$&(�Y>T��)<.K"dyɹ��>�%T���� �K�Wj�W\b��&p�Ԃ\eO/W�E@#��
�j[>a�z�Dl�0�>�!a�UC$)�BeB�R�Z~��}�5){e���K,�(�9����{ٍo�H��)>�F��E�������������|[H��U���1��\�������M+}GP|Ȭ�
fS��+����G3�I���*J1ELQ��:!��Cn� 6�Y��4}�H�Vm;����C��?s������<}���G9r����G<<^�=(^�=0h� arZNjVarvarn)�0���,S��.�d���,&;{���j/?���C|F�uu�����,�թ\-�<����g�[�:� 9�]�!�L�pB��'�?��n�!|�2(��k��:nU�	��[�f����P��Bm=-Bx�Qcm+3Cks� wM<}< ��6&F��C�5j�j�-���(c=c�@3�����~5��K����k���/Z�@h�6qt�{A9���������f�hgecijk������1i��M���S�<�<� ���4m�ٸivCǳt���M�/�Y���A��]��\��c�k�3��+i�3:�f,M��y�4А �����҄-�W���CH{ގ߶]xr?�����+�B��5H�V0j�����Cj�rI�C�"��,i`S�JU�u��ZflJYr^]�)l��U_�*�a6����2�=q'[��)���@�Q*��% <���T����*�@!��E�{�2_� ��͝��e�{��Y�����Hy$m�6��Q|�+_����'i,����=�����%Q�����ك!�R�&�Sq��*,V�n�M��5� �l5g��῁PS����T� B���_t�KUB8]��`D����xI]�\�'R3|!<�E����3u������b�wi�W})���rE�D�-TtÇ���{AD��=ߥ��`w�=��nns7��n�5�2[:�m]�wA�i��+�� l}K�h"5(X�,���]�ԅ!ѩ���S�����r<S��� Rw��Q��Ū��9{�;�._1n�����G��>j$�/0�W�`Pp@`��@@HP�( �a	i�IY	�����B !|5a&����%46��5B�����.0�����`e�̔A,�A�C�l��ce�`���3�:�u�Ѻ~��~� Bo7��v$�֦RҋE�`�x�D�����������qD4P��8z-��	�X�%oپw݆_����,t�u,��F: hC a��F�f&z�h}S+3c�������������6b!!ZkZel��3�64�7����MeL6Yb��^k���x�*3+kS�����;\�c���� ?/o'' �����������i��l9>}�!-�)h���y̨|zL!�M!/���R�K/㥖������4��F����VK��ㅃ*����BC�)�����H�*DN�I�\8�!_N��r �9d��A��6���&��}f��_z���̓zf]��U&�M�U)��zU�w�����GV�Л�]~���uG��"q�i�N�����VIRa�m�v���L��d�SJX���*.W�A����k{�l�f�R%P*`�T�!�\"R"��
�B�0�"o���6�t�/EX�UC#�~=p�i,&�B6w噤<��mw��ȲN|�����Y����C ��D��A��-����S�l֬��?��9����Q6� 5ä�eA`��ؚK)4������v������ZM�c5���G�9WM�]t�eC�A5jh������=漲��4-|䪘����@I䟀�Jy�P�����@��G�
U��v��n���k�OL�U��&�R	"T7�[
�L�
k��D�G�j��Q�Rj�4j�W�JUʦv6_4oѲ3���y���͛!�F��08<|d��@��`�Q�G�3T� B�@ �������S���p�������EU����)�B��!㦛X�23с���"��,�t���c��Ҵob�;��� iC��0�5�j����j�ByY��;f����Vo�˨L, ��æ? $Rx
�-�������'�?��m0�_Da�p!X�@���4a� ��[v�Ξ5����~��H���4�bb ��[2際�����i5��F�`M�5�F衴��Yڍ�r�_��ɨ d���+�B[S37Og7' �_�O�p����������5���������7�:;g�q=��f�Kbr�y�7���Vj3���UF˭b�⯴�[� (�I+�MU�&U�����C�o!!8�8���EABpT�(��ݽ�BB��3�Eda�-�Z���|�5cݡ�������Ԉ��l;�8}���e��E;�]y���J:�1�]!� Y��(zw�Eш�����n��l��0��7g���^l�w+:��)�qe���|�����rd0���?r句X�X�N���!�K����,��
zU�=f v@��ݪ�wY
�Y����5pKd
������A�E�hj_iM(cIp�p9H���7�@����![
�e�[�
8�#��Dsi8@� x�B��5
��?Y��a4�����֟)2�=%�`Z����;n�p��_�����:?�jj�����#-'$��J��>��	��/@A���?@(j�!���j�_ `��q�RG��*�%��
%8p�J~����*�A6((Q�
%j !�Cx����O�^�}'h�ȐQc}��4k� �|}���	B�[ƥe�e��e� 3Jj�I BK��3�p�p�7fke�lgjA{s��h�������T�N���E���	@��P��P��r150s��%k��fV&��
)�!$јD*��c����'�?�?m�!]Gb���T��Z�OÑ�Bc��@hl������Umllhd��o��,4ւc4l���CC�"�
����Er�����2\fi}n9|)!�}iôh�J ������������3R�#����������������쿴h�I�96��cshq���|zR-���^�ˮ��[�˰�J�ϭ�7b����(�c@� ����bK�~"���A�AQ$t�r �ä���!E��Q���Gn<�d�����v�:}�ّ��U)�����U��]����
��YM}4YY�Iu����'.>��h�ߤ=Ռ�ie�'#�mS��A`���>se=  ��E��h'F��1
t����X"
*���n���*yG�󑦀�J��k�ǘ-S�]$� ~+����b���\;w���Xj���J���n��fHU B�D���%����p̏ ���&�����(�i�N��]�� P�?d*m5��T6�@T� �!�h֚��Ǡ�&<E����30�̮�a���[(�WFku�Tk�J՞�d�����@������;&Fwt���r����3���~�+��Բ6P�EJBM�I��o���Rtk���w�\�9d�R�k���d���VPs���H:���=J�Ji���-8V��xՙ+�C���z�^��Ѿ�!.�n^��^���.~�HE ���7�06-+6�0:���g�CW���t���쥫~lie��j�����f��d2�\������3H��k��K�����#x���������^��T��T���68 x��-qYU	�ĤbZa���B
�M�S\�ϊ������@H�O���SY,ᦀ� s������)ZS��=������� 0hlh`bdh��g�=X���B��=�L�(���)k�F�~�����3J�9���BM����j�%����h+kk[+ ���;���.�N6�V�f&:����&^��g��u�ڒ�g̝���L,d��Dr1;��W�U�LMa]]iCCWN T���x%��)�j�l�9B�����$ׂ�	B����������P$��T���������OD��
�>�Ԓ�Y҇Eg���J*�g�
����Oi��<�������CVu�[���s�$I^����-&_�9n׹�r�|)��+�A�~�ql:�!��)>��=\q��]����!�!��xr8���E#�N�59]E]�G�����	���wF��휺���H�ߴ�gB��h��+E�l��s��MQx!�PC4�7�)4�;���d�'��D��*U�G(�&���m �c�P��Ty�΀����%*?j�����x�ᰕ���C�ZP��A� ��a��ܞ���
j �a��� �P ��ӗeL�9Of��`��j͉2^v{έ����/����莍66q��l�x�	%&�_�	��ՐH	٭��v��K$k+�� �=X>�M�[��G�	�#Hۑ:�H>KS���q�3D�W�#���rԽ���k��W��ށ�a�;���qL�l��v���ȫwCF����st����s�v�.��5����n}�<����|]��n<x�:=/*�$:�8.�$)�>AX\��OJN�89�Y�~��)�]l�}��=|]�r�N��킽]G�y�	��7~�?��A��!>n���>N6~N�������F���v�6V�{�V�� ,,���T�T�'�?��n����:���L���5��8Jqi媕�,̭@a������F�F��F�0i��FZ�h3S]s}++#`��0����������@��O������9Z��b�����Y�x�X��22�6���Y��aʱ����: ������	�������mci��A �F�RZ�:�&F s�;qs���m�W�Us�kXiv�$���S_��P[��+!ԗqdB�QIP���0���)ml`v�8�:�����X�����Y|$D&K B`�!sX��	U �� �|Q�:B$tq�@��P�?a ��^�H&hjO),�HN�_[P�4-u��3[N���,_���x���,3=�L�����&�����Nk�d4uS��D�'�Z�-tі���_f6B�F�vDռ�_���w����g��-K����g$J�T��OGj,�������3���4
R����o�� V;$� �۠uǣ7���Cy�QK�Tg�s�ư1�o�T}�(`E]^�-��F�t� ~0�"������^J�%���U�o����Jej�:��%�^*���	ʓ�v+�y+�]%�)o�}���bKHo*�5|���?C��<���)۹�.͂����5? D���4�,�f�R��Ru5�%ԶYO��;����a�
P@�-W=]z��AK.��gǛMOӟ��=��jYk|����_nUPۡ:�[��R�Emr�R!Uɤj�E�n�J@�T�p���L�p�'�_�՟C�>���ޣO���Oa7��Kc���{D���廸�P�A���[K�^���Շ���\��$`����v�F&���hScKKs[ksgG[/7gOW'W{�2�� �t�ErAdvML^}L^eLfIR^�f�(63�����Z�e��Q^�.�~�p�	w'[�q#���fM=:�k�� gk��n��H4͘|'���c������	��n�B���v����h�����MFR	>��0B*����)Lꇯ�B�s���� $��a�"��F��
�zz��������!<��� ��; ��������������)���i�rB��Q��ZVhkSc{3kC]s��Wx��~�\��M/'f��s�p ��V�/X����T��Fh`�0�}]�ZF���+�6T�����{����O�Z��8�����Vӓ1ԔjqJ�0�������k��ul1���B(#1ʉ0��A%Y2���e �p0�{�d�d����?���cJ��*:��b��Q��r��Ֆ������7Ο�~���7_�*Kɯ�}����Ǳ��D��(��z�'�Q�m����oW_�-��ˇv�MX�����Z���n��<��a�e�~�6AQU�#e���AZ�
Y�9�Ƃ;��m4ҕ]teP(H��o�~�J>K>B�6H�JmxK���P!�*�"�A85��r����p(���$��}�p��]�DI�J9�f"O����̕	˷xMY�5e儥{&-�;~���v��ܓFy_�
-8�8�ȫ�<��=������8q�򣡋\Ol���AO�(#7&�@��� ��Gs���X�@�l!ȏ2Y�V��j�0��+Qd��=F���1lJ�����'K��RB���Q�gQ!7��}�5)52j�����]*��D=C	%�H�)�$�F��I$mHې ��@4�v စ@(��2T}�.�$��B���aXݕ�v��G�;��wi'���ni��d��G/ܻ�0���P��1~�c�z�ƨ�ÐWx����6G;Z���S]t|��&N�t����9�Q��uϒJc2ʒ� �ɖ�8�]�l�_����w"0�=��8�`e�noy|���,7}㪅���v�>��)c�&��?�{�� _7K?Wӭ��?�˕�����7жu�|�P���o!��Ñ�d���?!���i�;���j<n����������Ff �5�Vg��`JK�=�Q^)��堝������j���'���>}��6���R�f쭭@l�Mm��-�-\}�{�Z��O���gV�s+�����JBq5��Y�t���������	�"x���ن�14tt��9qm�c�"�][�SZ[̊-fĕc�+*�15iuu98|�XJ���9�&PVQd�!�a
kX\�:f�,^��c���#A�OB����P2�@���P%�H �?V!IK;S"�+�ᱯ?����ϟ^�~q׽S��7ԤE��q�ڑ{��X*WΧK�X6��J�I��߲D�N>�/������a�{���_��с���W�������%� �%���$�;��-Uҭ��g�H4�rh���S��5�Q?P?��L]d��]�v�-d|,��^#�&��^̃��^N!|� A��$�sύ]}�Z1Z�c�jR�z�r�(�/~����j�TI�ȹ*5��L��-))JI��H��e���+J
SRs���E_^�G,�X�ն@�#����уW���LIa|!}�2DФ�QN�3!��=N$�f ��`��G�H�}�)���;�lU+�����@SA�N�:N;�����K�+B]��̺R�W�:�"5�q|��ͦs�y�r�s�-���]�ĸ�������7����m�h��t�[��w��|I+O�
Js��p���~������S�?�fh,T�*z MMW|x�^w9,���g)u%�Zn��w�;���q�A�߉�O\�����������������s���4�����������I��k��3�n���м�WW��KbaCBveFQ-�0+�TV���p�5NN����\V
���/�xt>�p|�6P@�m?* ���<�g���p?�Ջ&�6��-�Rښ峭m�<�C_'��kֲ+�y6��"����������W�<��c`ff1g��w��Ŝ;q�LO�\o(|E r��m,t�-P�f��F�V��bNO�B[q��u�2s��c���B[�����h��k���o�	�U��JRA%���T\M,��k� �!�`�K��ې!C��<&Μ����[8Ϸ�[]X�2�"���O�,��.�AR@��y�$Q�D�dʼ�Y�
,���%�p�Bd�����aQ(q ����B�g 7�0%b¨���Ϧ�Ee���}�`z��GW�ݻ�����4LF��g�l=s|�R%�K9���Ȭ�Ts��/w����o�>(���I;���V�Z%ն��׫ |3T��je��ɿc�_d��	�E���xGV¡��@H�p�j�d�{��_|���kQX���拉ZnR�f#�/>��M�>b��i[�����p0��SZx���j��]����l�IT�B^c3��,��z��^iJxU��3�����ܿy���KDv׍g3�ߢ�A��!LT��I�;L�5��K���}^t�j](�gMdt���(%�.��
!D��P51M*x-ЦV���U����n�"�O=>nッ/�������P�(�zX�e���ͷo�0�������-E�����cA����w��0���U�S��X�^`!���f !|Q�?�PS�j�ME*W�],��������z�;;τ��ssԂ������Z��"��s�2�s��q��;gn��w�{�D/BCc��C�ܙ����0�v�6����6qi���g�0���#���z&&�"��6��]@./o��X<}�2['o_Wo'�`�����n���������_�u�u�O��L{ !PT� !�Nc��'£� ��>6��L'��l޸t�� '/P}�J)���B*�SO���?!���i�W1$zy�G�j�T�H��D۳��}+�#��UWUٻ�3�X{��*�����	������9��:8�I�y���1 a��P���(m�,,-�-���Vh�M���Ҙ\J\�����-Zae�h`d��g����=�pl@EF���74�wv;u��C�: �X]��,�Iň.?/\{�Vj/��R@V��K(��7"����JjS5MXM�N�{ �HZGk�2e��F�H5�n�XB<[L�H�%�44:p����`�"$2�D>d�����C��2���-s�"Lٝ��c��ܻx�Ʃ�����zt׳�g�Co�?����_.�:��ւ��;t���y��%G����]�g�r>��CPBG��9;n�5Àu7���������ɴ�nO�9�2x��ŧ#���x7o��I���-���A��޾W���z!f��������m��
Nwt1gҚ�YĮc�n�8�pJC�ˬ�N3OD��Z��3uK�Ũ��Ne�ܟ�;���ka�e�l<t'j'(کM���T���bE<{��Zjč3[�_ڽ���Q�-_4@XZ+����i��RD�
�_N�,.�},�A�wМ��Ko�ν6�l)zʵ�����&P�FW�QAZ(�f{G�oP��I��P6�Ch���=���[.�1?A��P� �V�q K|��y����<V�J��V�U�����w�������'�7�Ō��7JoV�ܭ�U�CzGh���/<y�T�,�6���A�Y �����"�k��-�
!A�F��L��96� ���.�{���z]�
Xtt��S��v�
�i큛�.�o�w�g�,w�q��^&h+��910���ڛ��	�?��՘�a�#��;��H��״�I%�EXP�Qr�d�^K�O�g�j4�z9�x:���{�����ٰbтA9�jk
 D��j�4c�!(}\-�uP#|��oU%g$�X�r���������		���
��Q2��@���۟�� !l!�R���:pt��!��|ҤI�6�_�`N��7 �`�p!�M�� �6�v4Cy�Q�&9=�;�ʦ	���xZ�̴QF:C���@��L-�[m<�L����2*(�e��rxtt���܅�,l�sF���z���@d�Dk!(GO������+W ��I�ŌY�y��w56�\��/�-�|�s��J !܃�pҜ�酒Z���.��B��P�!���`I|8��B�L	�QȸJ)���F�����G��_�x��٬���|��0-=/)�ƹ+���ڿ�0�/���^�c�]����؄
���1�4բ=7�'�P�ʦ~/n���ydM�����E�bb�Ǻ;�o���r��WƓ�l��;g�C����C��jk��=g#rV�3i��c�bA���ڲ���SO�e����칇��4n���L����C�1�=f����J�Ev������Ȋ��箽�_'�6�fK���	;:xjuKow5�����㝿�Z6g�Ho�_W��1s�ֽ��Mu�n®��^֨W�}=k׭]7S~��P,�F�zcgXŁH¥4	ẕmW�(���?4�G���HMm$u��3T��=� m�+��n�N~�4��݈�so`����t�Ѭ�zs�-�^��wk����siR.eJ����֝�����/.��E���vX7t�m�ŏQ�����w��p��T@W�A*m�J�O!��,e����_2��4�7�G�A*q��erh�ƛO�����V��j�7�)V���⳵{������;��������^���Z��CAt���u����L�F��?zፇ��r$F���r6=*���(�M1�T���������ѓg;�;xz9���=\l��F]lL��c\mͽ�,5�@� ��L���=�к(S]�B8�.�+���������G�{}c��X~M=���"ј?!������!D��mׁ�(CC���u�����XGKo(<$2B� ���.(
m�(C��!�Ne�F]��Q�27ԷB��u�̆��X[�ϋHk��m@&� ����,^��511စ:C���DGK@h��2r������Yq��u�S���y�b�,4������_BfȪk�b}Y�ˍ1�]���p�(�U�f�C����I�2B���O ����B�XΑ+�* !W&�*,���{�:�᳗�����<��TTX��ȩ�%=� ��c�7���}�A���R����%c�s�^��uɿB%(��u���G��՗�_���9|g4wش�6�/���~���sv��	+�K������,�e0�Z|ٳ<�=�v߈��|��|������쾞\-�.�ŕ
A��n9��|܆�Sw>�ڼ�Rv�k~/'�|��B˷��}�v�۱�@������-R�$�h�5��}�Ÿ��ҍ��{���\yh��6�8x!6,���{9���\"z�~�WV�I(`~+�|�z%v��$c՟���j�N��)�ob)�-��%�dD���	��\ZǼ�O�u��� �	: �&��qT��GL���k������L�֟�a<'Co�C���4~g.����ϼH����;w��%�A'��K^�/HGMK��� 5�!j�i���3�o�/RI�B�̕�_B�Y(��!ɟ!�X�g~"Mu���/����������5��%�t��<-�T�?�ݶ�Э�����o�w�1������ffV��֖vV�����������.V�����S'��7n�E-�����^pL�v����↬���2zJ��cшI�����<�X�X�{	S�!��t "�����Qc�����Z�T��CY�,5=P-і����#�'��ռ�Tr��7��On��+� u$�΃G�zF�:::�������tP��C�s�ȬQ`�����6JO� �>��@g�;��H�ҤBc� +���S�^�`��'r�py���/\�@hh�����T����FH7(�!��������cȸ������|���\Ǡ1������I[����C�?O��6�-��eT�Y{���Jr׏�P<y��oBȒ*�29W	�BM$�R�5dFA�UR����'Qyy��j�:�JXIRI:!n<��
1Z��������~3y�MK��-j���8��m��}�"	���k�V?ĺ��l�c|N�3Q��t�}��9\��{��&���旋�m�]���\9f��"��������82w��WO�K&ʾ�֫]�tCk�<Χw�z�ճ\��g"��"��(�N\͍���zo�����N�2�l�B֭���4)�N����L�|p�ދ>��y/�w�5nƞ�g"W�����M��N�˦�oPAD5T'�P#|��ڈ�V~�G�⫬�7v���� �A���c�.��XM��{1�m6�y�n\靬6�h�(�y����-g���O�E�^��W�]�~�4����x�1if��V#Bu<�N�������Ϲ㰱Z{i5jYjZj�}�e��nr��Tҫ��� ��D�Z��Wۑwֱ�> al.N�	ۡ{o�{U=�@��-7���v��eɁ�8ŧq�vm:rc��G���3@���g��jkk�������������������bm	 ���9��a����9[#N?ō�{���t aZ	>���W�H��{��8�qլ/
�C*����n�h ��P���P'+Ws{w'ow��� W�ϒR�%5" aY-�e�� B���"����6��_��*a9�V��+�Z"u�(}m}P�����[xCN�����堙�������oj���5m���p��5������M#Rꢳ������p9 \�l����������������u��E&��YY�Z��Tss+K{g����m=:e�v#�)V��KI�D��U���ݻx�}��'�T�/�|N�h��3�P������N��?�D��7׳��!�p�%�p�C�=W�,���1*�&�*����� � A&� 鿈P34
 Ԍ�·�>E(�2��$v9�[F�e�E-�C�c��罗�Awc�6y|�F��5�ˤ#�����Or����u�\��{���U�o�r�j��Cqt�_C��(w*m����=#v���:S!��������'3��^h���n�Y�����aK5W	"���8m��*ĩ�A����3����
"�e�PHL���Hg��q?���*mG/�#Vs�J��/n�S�8���Pw��X�S�v�����Nܻ|%�^X܋���������N�]Ɠ54v�[���xYI���*o�+��k�5K��� 	�9�LE󿆮�CS6STp�?��|b�(�{M%zR.zB%z\��̒N��#��ݜs���ۃ�˴_�!��Zg�����0�YI�ӊ<��Y���Z��nqWAd�����OQ�Ps�P�rQ��Qc��Y�R@
���Z�`�<@�9�~5AEΙ�v�^�����~�q�o:�z�98;ά�y��� ��w���ſf�2�M�,Z����C��n?|&p�dO�Qn��.n^����ޞ�������^A~ށ�MG/;��!\G������	�o��xR{�iٵ������R��p+>���p�ę��v���GN��f�joa�ֳ0Զ5�w�0v�F�ؘ"��Uf�� �.tw0�4�E���������������[`�pO�1�^���Sʱ��Jnş!$3( B��Onl�B��0���5g�^w�����o�X�g��3�������������������x������	� X����15�17�������@hdh�:+"�&:�6f�`�K�V�
�,^�
@�63wtt��t��t폻�����������������i�Vl�7v�&m��&.�^�a���yL]{���+v?
��7��=��9:G�m5������^AQU�xUT�����P�`)TL��$���VK�0������c��x�D�;����H�fߎ�>t5""�>����̋��c�z������� 5~;�󢀑NjN��]On8���Y��@]L�o��y)��UE����g�=I�?�(����w~�j�'a�".E�I�&�b����wH�	*g�����.����a�υ��>Kx~�������o��}�܉��6nX�|��L@�K�r]�`���=|ݤ�/lb���&rb�˰�K5�����˧�_۷���-	��ܹ�V����<��⽋4���ҌW(�F���
� �`X�x��
)�4W@*����@p�ϛ�Pco�z�"�hj�є|�I�F��_p�翃|��C��]�`;/�vn��l�)a���Խ�v���,�g����׎3�<��9L-4{��%����%oP�P��P�KPӣP~��H�I�&5����{�{�o�.i�g*�m���-���b��1Y�1�p JSa�߳߾J�WuRu��8{�c玞���������Fxzy�����}�F�x���͟4�����e���\��<��t��.!�#Ӫ �9U��j6��	0��!>�fN�=c�� /� ogP��|�=?7w� O��~�<G�������Dա��	(�]����Y��9=<*?#�V�Wp+0L-�c �2�Q�'�?�?��!la=�URS�i�NPl��P^b(hgado��!::Zh�cognc�u���C=�HK�������<��G�����cӋj�9e�����\ 45�pqqA ��r�^��nN�zܾ���^�i��Y�꘏C�͌)$,�q�m�"Nb��M��i��]���1�����*�݃!�:�`v�������׳��l!������@(�2_��A��f�L���|�{	��VU����@�*���ܛ���7on��e����`J�q%XB^U}lFQ5�-i`VS`�	
��O�_g�^~��I|.HQ=���"pҎ�8���#'���]��^v[^�w0\�G��i��>�}������o9�y���RƊ��2r�����3X"����kk��Շ욷p6[*`�$��!U�}=�
�$�����&�|s����_�����7W͈X� a����� %^X�r����w
TIx>de��!�X����Y8@ �&^��^��fq(zf������c��%L�ԛ�rg:>����%�+N��3]�i:g>��ss���O�=��3L�����_�,�[��jN�����'R���h&d����������/-�pYp�~"���d�/�M����$� �9D���-���ȡ P�*����>P%okj<��&�e�����|�!����j��$��Jԭ�:p���KW=<|���p_�`oo��"a��7�p������N�v^�{%e쪫:K��N����3ˈyjA;9K��O�q�pp�r7>d��oOG7K;3CK#p�diDԌ�Z{9�j�Ax���H)����������������&8�����.��/Kϣ�r�!�J!��?!���u�7RAH+���p�w�>z��!<_E_WX���,��vƚh�"sG--A�51G��[��\�˭�Pz&zh�������ibamZaMF���V��(��3��tw%�G��=�� �.�..�'O߼�<k�e����"��/���}_�M�nP���Fd~j7�Fx�uQ	�������e����C��Y?���2�",��-���"���]����AfՁ狧�f�ņ���b͒uW�߿w۶m���_�~��cG��*ʈ�bC]\ԫ7��/^�x��1�Lep���+�����]�h�H�p|9��]�����~g��ݼ�;�Ǧ�հ[?�~�������B_��n�~2&��MbvDT���'�R#BC/?{v+3#����s�M�J,�<s�S����'��%)C�b���=��W���-��v|󥹓�ϊ�uY����䆼�+gּz}�'*�{tl���U︿AΦ:-��=����G��^��E�z4�zr�oP��ϋ���ל3_��|a�ł�_#xe�T	d4%�zN���X�.\z5~���}�B(�]���}�jz�ٴX�I��_�\ygɑ�Z���^��mg�U,���A?�9��L ti+P�!�`ʺ�.��O����K����c+{�H�������D&�`yՆM�Ϝ�x�ډS'��==|����M���;"�w���(_�>AÃ&������I�t����x1���U�V�+���W�R��n�K�L����k0���=����������̭�C��ӑ˴�yy:pL��8X��[Z�i[��9X�>b��y�g��K���gd�1J��M�-  ��IDAT� B<� $�H�	�����B"�� A ��Q+k�-Y4Z�n����564��j�7�DoL�&�z(}\�12
nM����h�����t������=m��P�/>t(J�X��c��ǜ�	Uq�������
3w�[{G+k'''_oO_o��24�?.��������j�`?r��m��-�p��}���o�ɑ���RFR#CO�����2��� �-"��IM BC��K4�e�u�F,S���mp,�@�l)�#C��"!����'p0���j�	B5S֤	��"�&��ԅ�rx��+�R�@�J�M��C�6�8�kD���g^>;��Tē3��{��jF\xj�S���qO�$E���1�2�_?�o�������{�T*�|�P�I�b�	��+U�L���W��[M�̖. ᬵ[���Hl��%4*mϩ��6�I�(޲�𳗱?�����~���ˇёOΜ98zl0_"`K��Kl)܎�+�;���\���SfQ~vi~y]E\����6=?x�������?�/?�iB�K�]���(c75s�:�M������g�����@ ~�?��U�����P.�˾��N��ؑ�0�j���דY�+:�Q!����
ʝRY~#ć��>hǓv�qq(��#��,�Q:���_"RRU0��O�����%��KɹDƳJI�m��-Y��!ng�Ul1<U
�'Х� oH��0���3�G~�&��"�By/[�)\���,����+�o߹p�_`���ۈ����N���D22�o���pO�Q~��GN��L�e��%g?(�)�����rj��5�JFZ��-`Ř��}]M-�Yhx|O��ës��h� �yAu�C�C7;P z:�x9Y���d`m2��X���|tȈ9�M��@�S��@ȯ����O�?���l��s�c�R��avI�╫�::s�\P���5=����:8?16�26�6B��16@�j�t����P�Z�g��C 445����{���
P&�פU�V�b
�k�+k�+�K*�.^���bam67׿@�A'[;kgW;���fm�wv�ƓVns&G��~@HI��$�S�p�XBf=)G. ЋH�r����YP�!�4goz������Ko�`�_�� �B�4�ܗ,ᒑ��&/K�b�D̗�ل�ҝ�.�s��(���`ԥ��R��$ze��fT+(�rj�_̭/J��"%�VA�'�Z:ml蕳�O� �p0�pw�B`Ic;�����CWv�Z��������[�Q����-�:p�d\bҫ�WQ�/c�^�D��F=
>z����K���E\��������#�^W��MjDlҝ[���<��4&�ILzXL���Sg.�pa��};.�綵��:����~� �`��4
�Cɍ ���NP╟)���J�<2_�Z�<h��;�G��b��A�/�7��[���6Wս��ߠ�P�'��t�@�K���˯��25�P��-Q�FS�rAU����V�k,�3���QP�C��y���τ,T���V !l!PS�͒� ��^�ᾲ����5�
 �\�X��5k/]�~����׮����:��������E!�`�`/�`������u��`ؑВ+���q����<lji�0���^$�Z5~�"Ww[GK'{s'[S'K����>���ބ?؃ڢ-��4�`(|E�������i�����ӧL[ �-bg�3�UaM��Ƒ�x
O!�������o 44��`)�
��e+��\��`b�6l���aں���憆���>�Z0~FZ&&� �aR-34��t���[ �6��ccb��Zؙ����9`��蒧�EI��9EeE�����JHye���\=ܑ�v���~�p]P����5��������yƂ%�] ���|c�i����2R�\�M�֤��e���D"�q�� ��e�B������KH%ȿB���_ �׊�(�����4~4	č`&*e�B U
�Ԛ��օ�?S�����y~䳢��/��E\/��U��I{^�Q��,/�IqrDޛ���Ē��Л��Ϝr����W�%"�H���T\�.�)jbH4�w#C��.���������n+�jW��8u�n~u��S����^�B06�	��7�޿r�֥�{�#��ȁB(nC�֤�J�LA3\�T�e�Ŕ�\n>5;����O�$�Pb��$��GV�������mz�Qkz���l��3�H`UjJ�&�
e'M����� ���C1T�ae����I���_g��>׹�&�sc�咧��uB�ЕBh�i�����}�v^��w	��e��"9T��=UX/�S�;�mr�Zʕ�A}���? T3�M?,l�tn�H�Y�nd5Tx�\��;I����Ȁ*2��9�/���[!L�P��	�r%J��]�f5 0��#B� `������3x�!�O �us�wwtst���5��e4e>e3��c�}��7�u)%��jBF9-�T�=|�ĹK݃�<���'|�|\�@��no��G��&�?}�ܩ�A�L7{��Y�FO;|�p�?w�Y����@SKS7{{?��)Ӗ�Y ²
�On�}�7�O�)���V`�58���ѦV6�FF����PC���К���kAM9hb2��en������ -S=#c+kGw��37�.{U�P��_�YX�[XV\ZY^���������7����M������XY ����-��,,̴t��쬭]�g-Y�����k�X{�7q��_?�z�`�.��ͧ�@�i�j?���? ��#�����<���"�#'�`?WW�!B�F����&�8�-�&P��'�/��[��&��Q&hT�<��+�U4�ݵ�������|U��yqDX��{�n��ސ�I}Z�^��$/�qaҋ����	E	n\Z0k��7b#cd"�H���\Q3[� U@������p3��|M<ς�~K5��f��2q����'�?��Rlz�����q?>�yb�38o��%�~z���3� ��Jdh�	
I���3]��=g��8y�����cf�7sY�v[b�L�{���u���[,?<�x(��4~b��s�}�i��.�5��e76�hC�� ��C5]���f���&�K�2��*j��>�LО��;5�pn����Y�KߠF�{)�j h�3���L���s�W=s\~�w��񛓊PCT�+�PV��d�f![@��IL1XȖK�1p��H���k~9�v�_�孂Ə����Mtq�_'if!�'_~�D�%W�߳��l! @��W�^{�����x���7((�����min^s���5�N6�����.ý�&������7~9�8}��{�^y��U�\X�U�K/�d��}]��B��G�y�kz"A�y9 �fN5c�H@��1!@�Q��>���n�~.� ^Vv�v��G�|S�]@�,`�T�;�������6���L��hbjfh�oaili����Y�[�[����F�����Q�&(#8V(P���Z��Y���LL ��f��NƮ^.#'�t�[�$�$&�*��*��<�������S]U�dժU�����aZC�C��蘘�XXX���i6P)����,L��-\�����+X{.4v��:W��*�SL���!�!㊘�R��I-cp ��$UUPE��ǔ�U�A�L������ q|9^�@B�"�
U`Ǆ���D�? DjD�:�D��2@
��աFA�/_�*�JD�2�Z.T�*5_�̗���+�><{!�Yx΋�/�
"E�/~uT�%Qw����<(�{T��qћ���[y��rc��9u`��)a7�%��j�(@�)6	D��6���+�b����dc){ٍ�0L���{�gW�U��q����9~:4!�R�+�^�q26�qj������ԨԔ��Ը��_��tn�\��+�ó~�M4yU��ەw1?
�!��SR)�}�ʀ�ۆ�N�+n,��f��i��qǣJ?_�=��ǌ��kY�di7A�[%o�+'y��3���xpP��DM��?ބ'��pd�\iU�{�$�=���
��9��Y�rآp��G�OWd�B7p�:sn�M�қ��?��uI���t�q�"*����`��R�Y0K*
2�J%O��3[�yx�vR�J�O� ������j*���	�$	�4��]t�[���*U
��U�_e_@m��TI�bhBP+�{@��V�I��j��֮��=���Hڴᗝ�����K^ށ�#�����q������KcC���������){�?z�ź��2u��{��K"Sʓ�k2K�3�ș2π�g,t�us�p�u�3iT���}����5��~��f:Xz9Y{;��o���oL���`��#|G��yۃZp����i#��;oX2k\������{��'�iل�@H ҉d*�L����߿�w����~B����!P$��vǞ#ں�C�����޽$����P��mmhfi`j���P?0(j6���w��w�Y=��������������������Ji����URubv]fAunAEaAEEi��S����]�t���= OGG��m���\��[�gfjlk7q���'�M[���}����y�0���jL	6��&�@(�ъi�B*���)#*A*)�J�`����\i��!�@Df� �m��?�)�E�@����R�S���`���f��Y"R�D*�H��T`g&���/>v�r��'�/ò^>�}�y7�����[1wA�b�ǅ��yX�89�(�c�;�g����o^L�~����"�D���ql��c0���{eo�q��1��8�\t���'��{�����V��������III����c�㢎�8~�҅��P�eJ����[Ȋ��K�QD�}�H�]����4"��۰�f�����8�N�TB�6%����r�bR��3���.���*k�1���T�@X���`��_���p�����7r3�/��'�Z�-ԝU0lnj�!�"Q���9]������g�֟�?��p\���j�	�v�_�Ll%(!��T�R�$|�Tu�sOR�`(�4���R1�͜��t��u��T�z�}xQ#���Dm�D��R���>��.'���T���D!�j�8��]��]�J{�������vC��6Q�o ,y[��n���$�NSs�7�qߡ��O�<u�vP�Dop��C����}�z��& BoG��ç#2 ��k/;�\�?qeDbqbNuzQmZ!=O��lܴ��^n�.��^NcB|A���d=:�kڸ�/��ri�e�W-�r��˨ W�сn������fL��P�, �(�g�	��u������)b�bDUu���  �9d*�L�����������b%��@X�c�]�xcb��k�t,6}����C,�t������ӄ&�r���6ֆvv�v���Yy���EY�i�������mofjgada1L�@m=�-`ER-��^P�[T[\RWQ^��n���4�_�t��=����(j�8@AB��� !���p���֞�Ѯs5b��r�/�1pK�J\��YO˨�f5�s�9�8E1^^Fᖑ���(��2Z�X�z��B�B>!N�@��	���
!2	b���X��.S�*�T!�J$�O.�(%,:����n�Nxy7%�^jԝ����73cne��ȉ��//�~~⃼�	����e��{��5�G=�{&�MX����r�2�D&���{��-@x�M��Pv��������Lj�͌�C�3w�~y��\��c{�޿��,:�Qt��בᑑ/Ξ?s���G���4E3(�~.��HP��Q�J?@u��ϳ�fo�4A��P�
�WC�o�lN\:��Edh����K��.��Vl���	b5E_�C(Si T�� ��;��<M��ʺ��k������FS�t����,ӝ����d⩜��Ѓ����&��&d����
�4��}޳�%�$�V��*�L&�7�h��DW� �d����Jm�X+�z�g֦W3}=o��UǞ㚡է�gӕ����K-[��N9�3�	���9� c�մ�WJq
���8��'#w_��Aɕ-Kv��s9q큰Yk/�l�V����z��\�����J1���ٛ�s�ĝ��/�z���g��m`C8d(ܝw BpL t��@ �w<�e&-��4��z�m+�ɯK����
k~@��/N7<��T��'�M����U!:}x7�(8��(��>6�3����^h<�l�����CJ�P�N�����bf�p����LR61��UT�)�dU���lۀ����'�?�?m���k7i�Y��ڷ��*��2z��%f�(sC���P�_\jAx2�����������~G;��>c�pC��>����0=m�)��Z�����Y�Y��(gd��sJ�e��JrE�C��!U�-[ini�g`���;dx"�y�@h�� �q����� �fn� �Ȣ<I���UF�ߔS�i	eT8��bS	IYC(���j~@��a�B��(�� ��w���R%MlU��x��7xO-A�̨xr_.�D"O$�Hd,��ԉ��y}7�ՍĘ;I�wA��$�=L������$39$�嵴ć�	�W��X�p̣���T*x��L,��y2��L)���}��MS�1T}®�v]x\@o-��m��[�B���!Y�|���G�ſ~��Ẓkяo�~|����QO���I�qa�h2xD��@�����������s+��ƫ r+�(1��5�DW�Y���g�y�$�*h��G��I+���U��wEΟ!T��P�R)5��H��9w�6�CȒ��E�(*(dQ$z�+��e&S0F�*Lfdi��?�Db������S/[N���h6!�~�`��e��qo��߸�^�\-�+D�F����j�WP��5��)>֩�'9�6�=+�v#��o�_�-;����B\��uW�z�?z/K�o�Ƭ=w/�3v}(:�t�k�R)]f���5��=�nZ����XƜ-O3�?ec?�����S||~�Ϙ=��9�⩳�����L��{�~�uy��3�.c�}&���Yhֺ�!���@g����������s�H ���ʉ����+fD����b�j��	��E�=l��=\l����c����[��;��ގ|���u�r/'K !_'�PX
AxM5WKWkg��&��+;�e��������G1ɹ��2VA%�#����6�,�N �?��۟����C��x��k�̌M̵7o_��� 3������Z�]A��(�L�u�������6�pE�e��%�G��h��W�����4tZg���=�U�4�%`UF?�O-�gV���u��L`66PDU�Q��Y�������!|������@����	�{�������]��;��JK��������S
���%@,��q�����������>���Yg��z�k͚�Ia���sˌ�����f����U��%�\N�e��Qq%�Ԫ&G�:���,�M_}*��[��t�W�Y��ʳHbA}K~-���=ԛ̇#�E~kP���<Ջ�g�(�PާB.9�9�>Đ�t7��Q�����h��6�1�E	Lx��έ�2kY�Z6��A��S��u��kw��޿�б��]<r|����'L�1}�9�gM�4nܒE-����i�+�Ϝ>��M[�,߽wÑ�;�?(�,D�'�%�Ώ$~'ȯ^�T1�j�ݍ���$���Cj�_Ͻ�<�h��p�y'G/�x�~:]��;|i�����}c�{,��s~��ث���^�j����"r�+e���g��k�+�JLlBB���svEW4ᛑ��֜;���|����^|�轌Y[n�>��a��p"�A� ���5X��B4Cs��m\N�[�c��9���2�̂��&a�uA����QrѾU���/ɶ�MǼ3�n��v���鬚�^\k��>�C�'�z�}�q^?jÕ�!���:~?����H�������V($���b1N�^���w�a��Q�<$O����:����!ųO<���8/ٳ�Vκk����Ť�d��W6Sﯿ\��Cv<,V�g΁�6dӅ�+�Mr6��*�!�ț�n�8&B� u|d�ᰱS�EȬ�'�<�j���돛Y���ZYz�ꚢ�	UTe�	��4T���A�fzZX}O'7�I{��~��aF�v����%�}|Alrq\JI\re|��uP�XC-s}g'KGK0���`m�oi�kga��d��hqP��~Ü|�A��f��BgK,�p��цy�/��p�8G++[;�[��Eg���i��bfQ)�����&W�9(>�
"�������D�z��g__K7g=u�(���-�\������XC5�o�F
�:h/{U�rT��'��BQA[IQ.Bm]������+��Y��"��D\TnCZ7,?��Y�v���j��-����luLTd"��BXQRQ��������a�5��;}��]' �E�O�,&�N%�z-4t[0zΑ�Ҷ+/K�Fo|Gy���w��,�H�}�m�����������*VgCRN����������9�?� �(By��%�4�FI�� ��v�-�&"��N�]��u�%@�t�#�d�6*�q�O��zq���k6lUQ3�`�UTl�M�ki;Xێ23�ܰi��Ȕ�o�o�r��̓'N8s�Ut�A�qV'�]#�|*�t ���G�Z����X}�G�v��-����֋���i��ӎD�Q��t�����]ݵ���n�D9�b��U���d�X:�������Q��^D��mh�n�(e},f}&u!��}�)�]r�u���L#�Y�9{���￝E��y1x�٧�s�\|�PFo��W�۫Q�zԁ9�"�)�ge�8�;WZeЂ?]88/��9�L�OeTt]}�t�t�n�}�i��]|�$�� ���b&�Q�<k��,�i���G�\J�.j�F�h&��ɑ0�O��P$��"p��q �oCv_���s}˕��G�<{-����m?w��2��m7���6<x�)��y����咳�>��cȄ�/��*��;�H�L��IG�OX}*��	!� EL��gwd��,"r�r�ȉ<�l�I�),Zuz��?Q���!Z������jk��j�Z&�:��G�{��f�ɋw_��ꄽ����G%��SK��).n��͵sr60ַ�2tu���� �iAOS��!!�D����,��M,�4L�����-t�u0���,�٘9XZ�Y_��<$�8*� �0���_�(��WTQp�z��ӗ�߾}�-���g��E�WQ�_^S����h�&�PI]2�����U�TTU1��e��������E��*���0��,M��2:[X�"��4��r_�>�W�ȩ��U	"r)SV9mӲ]���	Z��q�s;'UM��"hOS[[KW�9hCM-#CSG��Sf��qd��ͦ�s��g�ˬ�*��y����}��Mg�~ۘC@��D��l�Ob�2kZcK�)Ҽ����OŔ�rzkY#����CMF��_�����F���8Yw��}h"���³zp��jOQcO�;��#x�w<�+�����@�~*$�'�=~���E��QWnE�[��(���/������*�1;���p�Thb
-*��u��GqaI���Z�@.��Jpޞ����G$���\p�7���Hh����7���$�<�4u��D���?�w��MXq�*F3ꫪ9�%G���?��ك�ܷ��ɓW��yCd�׈��v�Ԇ�H]+J	�{�K�)"�O�u=q��%Mh]�G�p����t� �9՜"J��:QO5������ȑ9""W@��jx|@��A�������	 ����*��)�Kԋ��vW�G6�S'��m�D�|q���������4�V�~��M�Q+f����>!TRJBCX��Ƨ��*[%u�&0����6A4���Q�DuB~��W#�
�O��χ�E��}��;��bz���)�|���ң�_������y��ZZa��֙(	�p��"�gn�
����{����.d�ٰ��*DH�{H��u�����"I9�[b��i�71�c�l^�����'V�?dn��9,�����������������kd�g�ձ21�51�51�86��������!��b>z���W�Ǧ�'��H�'$�]��L�g��fmg��j=b��ر#�M���P.�a�V6&:X��*�Hc�����X�(�[��>����ֳ�lbJ=%��U��^\N+�l�����&~�������*B ��r�╚��Jj������F�=me�s���|`5eUMUmup�Vk�ad�id�fb�����h`4d�E����UW��R��W��7P�i� 4�!��WB�et1�)`��L���ߒ�^$�X�V��R�� ����/cj"���kh�.��4�tL�L��&�X������L�f:�x�\QH6u�i����L_�7�]j������+����������xk��æ��s�n��a�R]�1�}�QV[@���3�fA�?E��&�r�-�E�D�T$T��'6�v�3m=�8���:���S���fo�u-�z������箿�C����x��ҟE�����/O�?�h�C'�W>�y�{�aƎ�^���+y�2�ꝨS�B�=K� Y��I�x��l�ˌ�15ߎ</��p�Eq���\s�qA����h�|��K��U7��]1sp֎7a�--_�b�(��r��ӝ��8tm��[��r���]�N\}�.�
L��]��N��W�y�/��W�'^d�O��`|"t!�n�Φ"�#B�EJ������:a!Y�cw��)�_A��ί�OLI�\��4�""O�p���|<�M)�%��;k��4�e=m��-(�)�	Y�������_��o`o���-TQ+E��^�/��w�Iy�M�S�=��X\��ԋ�wg⾔��Җ��z��1_H�����P�N��CG>k���	;k�ZO�l�!���%[���3ڑJ^K��� ����혭��vd��Ak^�q���ۼC�bi�N3\z�E��D��B
�<M��~�{?bϝ��Ǝ�!9�v_]�����:�9ل�W�e~�T�f-ٹd��՛.]����mذqN�^�.���^�l�l��m��,-Ll-��- �a#�y�-Z��𹧇.���&�,�����&fT$�W'���ܦ������a�h�9�q���1cGXZX����E�U����.ր��( "�j��7�Zh��Y꩸�錰3t3�q�0�1���������솤�AU�J����/`��"�]~�_E��������	IY��6�Q��bԌ-�Mm�u�4��0��m-E]me-Mt>
mЛ:趱����������Oj���+髩�k�buU!;j�(jz;�y���ʫ�ί�ʭ�)�����m��I���n����@����G[[k[+�����������\���45wr��4u���m7q�	"�D�&�B�iʨ������k����g��/��k�?�ʨ�Z/E�W_x�u;��]&s��?]'��\�T��kȫ&��s ���p��F0�ÿ���7��rB���l��	������O�	��mx�L���bt�h�s���2%Y5���W_��ݒm�����Oݷ߿�������S�˳^Ňl<�m��]�o/%W\|r���#�^\�(L*�.
��:{���]�='-I��7\x��lpY;��G���������׏�ք>�L�[r!��}��b1r1�Z&AR)Ȳq�.$f��� �ߐ��=�/�ܱwՎ�_��y}���{O��}2��I�F��{8{�k�����_{����Ԧk�^��V	�W�p��������o��T�>�j�5�^RS)U���ZA9��:&�������O�����^���K����h���<�	O5�,q������1d����<��Tޏ�T��g�i�L��T	�HI=��PR�K���Վv� �"e��.)a�g��������YI�>x1��g%D�bqsE���GX��*�ҳ�\�(Ջ�R�A��Y������k���U�o���y�f����ND{[6�x�C��'/ˣ4���YE�Wl,�w�8틷���$���zN���#�f��?~e���1F�����$ߥ�����/�
��ur����l<<zʲ;O��D���Ǳ����ݴ����{���.^�n�.�nN�����h��`g�dk����3r�������|X*>2�2&��]��Y!af��m�������{�x�!�ۙ�Z��������������q�s=0���7�a�6N���F�ֆZ�vj���}͆�Y:�ںz��y�R�^��G�*d���S����.?�� B��j ¼2b����>�J�:Z���&&z���F:���*�3=]UuT�jJj��GEp�1V��@�HO�P��Pm2
"�׋�i*�i+�誨���4���&�<$��Idz\~]dN����i[������sD��]CK� ��"�'��������������������~��)K6훴�c��Ӄ�*�8a�1�Ax}q�����Ș�=��[,Z����u��e��+�҉]��ً��t�f���$)����<I>F��+"�+���
�3���ӗ���I
�=e�/�dĬc����nZ�f��3r��2^�j�j�s��S�r_Q��Y�	����~��_mF����n��~u1�"���K�N���񮓗�m>Y)F��xq�uX0G�T �bd���y�#'xe7�d�Ys=p�Ce��a����Ǽ�J?�}��r��#�3�]�k�R�kz�����"��R^\XGKK���]�kg��9�eI5�:#���,6�+Dn�Ҟ��Xw%���Bа��m9B$���l��4j^"D-X#� �4a�w���C!�_��O��F��J��\%�*�_�����kC�7R�7���(@��zaB6I��(�@���JQ 2�,ȃXB"yx� ���fX�k�.����	�Ht!�5���g�x�j;R#�^��DnE�ߐr��Ԋ�RJk�� B.<�t
ZY� ��sqs;����7���b�)}H9�c1�;������^��/���i��VVE�|��.
��_����H��[ګ��<�L6.AQuC-�[G��R�Z
EڙGa��"��ߓj3��F.�G�Q%�l<=����W���G���~�썓^�w��0��#��<Gx�{y�{�t��*[�c/gggG���u���/�㢓�#R�ާVE�VĤ����L\R��B�����SQ]���j��W@�������	�B��lM��^�v�n�`>`����0� �1#<`\hi�cm�"�7�p���3�d�����3�����tBdZ�0���S�[����X��Q
*jK�f�Yn�0���FC�����n����U��QU�RS�TUQSUj�)������zJ BC]E}-Em��:*
��2)�bT� d�b�'X�,~S�<6�iDjB>!*�D^&'�?/돨�\�f�����ho�l��"4�15���pq .ڰg򢝲D8�^x��.�H�@~M}�[�ǫ�K�NY~c���������,^\E��'YN\y���rWh���/�g�������N��Ut�+@�D��r�@>�'����x\��Kv=��	殻I�hR��D|���^̹�72j����s��|{�򋓗��be�_�?|q+:3�����]��u������nJ���y5u｜)�@�|-�|+��g![����y`��Gs'��C�+6\IM!#n3�>Jm�:��	Xv8�*.f���R�^9^�:#��]�O.�"�;�i�l��IqI�ґ���QV�#it$��o�ƛ#��o�}�I��#���{5e�c��݉��J�'�� ��br��*^��71�#R^e���������OR�Ͼ��^�"�"��*�]�Ȩ�DR���.N7RAmi�����8���c�&��@YE(_@ʺ1�8����sXQ����\���|%�X�g#��gn��׵"�]R0��k쇟5� ��H>�CH5���]�w�E���=a�-�ȳ|ޟa������� ��D��Z���#>�5#��J�J �s���)�n^Ǘ�ȯ"$	;p>�����KH���Z�9�����/lQ;���$�w	la���1����3��'j��U�<��^��j�"�B����Hs��]{Μ������'N_���3��_D������	���{�22"� <��L)�I-���P�sY����GaT��u휬ܼ��-e󘚛�j���j)h������|
m[S}=]���L�h(��Sr���y��=��7�ѻ�Ȭ��lRb=���]L-(���H��5�U��O�M��"�]~��_�#�M��.��6s��9�G����*a�4Uu�5��Ե�Te@.B�u4��uTt *�D���YP.Be��`�3������}��W�U��G5c���m����o?}����>V����9�\��&�� XP^A
.4�53���pv��p���&��A����_���L&�Im|��H.mM�����wjeGX./��C�ۉ�iF�1:#<&o5wO�����8����5��S���D(��� �o>y'���/c�Y����ĭ�^�P�o���q���t���5x^_��	��WƼN{y������^ƿ������7/<�{��v[Gq]㋨��O_>z����	�g�yZz�rʾӱ�v$���e���oK�>˴���Qf������|��j����bk��V�M���8��jR����	�<7��-���w��JQ7��;�^� !�eV���|Zuf]�Ø�?.��mŃ���J���%���E<$��mၗ�M�$$���|^��JZD���+/�&Y��)�#U��U�<���UP;j���˶Y������G$�ݾ���QKw�>}��sv_��\������ͧK�=p����׋>��{>:����#Nt4�F(�����D"�XT!�s�w˼�^�]��`�Ʒ������6���hļ�E��f�轴Y[��"w��s��t�e��;.ƞxR�1�8|�{)M��<���]��u���bt
�Y�]���X�:�������
1�R(��"�PH����t~AI�U̶>JsW����k���y5bt
�ª�D[QE�.��B`�+X�"��+��%8~�ӌ����B����T��qu|���ڴd�VH�g.�:r��װQ������0l�0p���7��������ٻwQ����G&G%�Ĥ�Ħ���eҪb���{x�jc����i`��k�6,��O�2�j骁a	�� P���������9�X�m�t�t썵U0�X̀�^S'M�=D� \zZ!3��������:S~yMdbFbZ���^�-h�4C���VCY�VQP�p0�Eh��頳�h��wU����:�e�D8i��7^�>�HN�M�%��.Y���M7g�}��t���V����LL��ѻN�.v�Phkgmckem������������w�����Yu��e����WI��	��q�·i������%��2[��"u��l<v7~���;/�����㵇��M-�`�J��bc��＼+��,8�\�r��W3�]�r�M��f'[L���xzܒ?���,��1}ˑ��7,�s�u�N��X�����X� �̭��2���{�<>p�D��c�myp�f޳�Fq+r�Z������g�;���`Ժ�a���۰���H2��PHL6��³[�9�Զ�bʎρ�"F�9x3jʚS�=�j�"D	���*C^�y�5���TK?�$��1�U�߼��(.�u�����W�^{�XFo'� �/�NX}|�ՈIk�<p#�z(���s�柸^����-'�o:c��*R��V����W�z	���W=�)h�D�)��*��#����*��9i멛�eq��l�|ޗ4J��M�㫗�g2r�ɇ	�\OԊ�-�z����ZnW��*�c����x��J؄K*Ē2IS��9��ep�e�7��''�x� �xS��{[�6}OV�z?r�^���c�L����c�H!ɣ!�_����)���ߪ��
��Ɉ���=�D�3Cݧ?
+��؜���=���"����&cԂ,�\��6�hS "O
"�b�q>,�q��|9�t�&��%��H���
6X���ݎ����Y]�̮:fG���a�{.�r��W=}���g����.^Nn�.n��y"���*�]\݆���Mh�����ؼ�����y�I�Q�Eq)eq��IU��-0���IM[S�P[�PK�Pma'�����������LF��=+Sg[kg+c�<������`̴�}=�W,]��t78>,��Q��",��-���?��F���Y��n��x����Ag�:Zں�Zj�:�(h��/"�RW��T���.�U�XU#uu}5%E��2F��j򜃶^+��Hy���Ϭ��������K��N��|V�udfn.tt�w�p��P^_
��[�"�4�tv�4c��C��2s�a슊�ejś�jt��Lt4��bLQ]t	)��_N��`�Ϊ���ǅ7�w�8t'����=��l;��aDFS�[C�\XBb�k��<�����I�!��\9�7���$|@]�KYm���bV����h`u�xQo2�^Bk+ 5'�r^'�\y�{�f���ѧ.&���q�z�ν��oW�J�0X�zTw���;�'�_t�~ޙ{��e�U7q��K*�揠z�Ga?�l�B�t�g�g$� J-璛�z	BnE��)����y�.����(���I%�o�$��`�3kO^�~����+�Z����qiUJ+R��yW�������*Ηk��/=O��a��Hu�⣌;��y��`%�s%�#��8�$~Ѯ��κ6~�v�ZT��W�٬�Y{.���u}�A�EH+�,>��i:e��������#���Њ�z6�zx�e��K�w�%�!��QO��8QK���L�R*i)�����Y�;�<9��8��ߪd����h�s7�yھD� �+��F��-/3�7��U���6$���i4��u�w���J.����5�`�n����i����HC'�0V`7n�"�bH�t�2�](�VH�!Vs��!(��P���EU,	��$�E�@�xV��S��ct5л@�,A��ջ���~��S�n�y�y��8ڹ9�::�9�::�9��[���θ��z ��S����=��̀\��.D�XK*�N*�K�
��|ڼ�c&M3��2�1��5l�L��L�����aռ]��̇9ی��>>`ތ��gN�>>0�wT��a#ݝ=l\�LLtA��J�]�-�}��U�Դ"�L���z���?�=�����"�{�(\��Q4a�l�a>&f�::ZZ*(j���iBU	 z�U�D��h��h��q��T=UEUE���������퇯��*�yLnLNUv#�B�Í)n���ڈ��~kFN�cmk���mljdekq,�m�fo����������K���k�Y�����Y^�òj��Csk��<|x>.��"��2�[V�k����֝y?s�IǠ�~���/�5|���K�=
ϭ�fU�J���F~	�[րRN◓���r2�H*IL ����ȕ.$��~@�򇨡	���D�g�"�f�"��X��D���P;���O��o��^�������/��Dͬ���<	A�^���c����Ӎ�v�]���r����݃��0���x��M�u��Ǝ��R.�R-�/&�i\aK[{gg'��a�;g�����&)���(��lA:�"��Ϸ�3���B��B֝s��Gm�L�_�M�u�����?xr�U��w���<;�$�IBN2���vՋ*��T��*Z[����RT�/#�=E�_�i�?A)E �C��p�Ʊ��Y��-g�>�i�BJxy��H�7�ܞ��2qۅ�I����`}R,@��DU�L�x�jn��G�v\��}�q�UJ�p�Z4 ��*^7:���B�Y!�(w�J:�%�η��3�s�,�-�������#7b)�K�?I�մ#ۯ�8O=�P�Y�{��BJ��B�C��p��Ϻ���x��@(��B�k�Y/G.xB�r�n����xb]���k"$2�QdiE������BP  ���D{V����-@5��Zf�*V/��Gd��2���������}���˷Ehg�aifgajainaceakmngcأ�)d]*l���]\<n�y��ehXDrhdjhL��ج�	9�yQ)(q���O��Dh��b�� ^�g7;w٬L#��G���v��������5��g��_��Q�����q�������������������������p��/cޥT�K!�DH�*!��J*k!�����_D���(��W�&,�����������������穩��5������#:���B�� BH��jm��f�u��NH�󸼧Q1������ƉK.�{���NzCwଅV6��Zj�:���z�f��֖VV����j���6⥅��˘)3Wm;<�a+ϙ枳��I ·����Q�U�eay�1�e�e��rB<�.��UJJ��1;�8����d�(<��Mjա���
r�
������Bԅ���J9!Z/���&���`"�"��TSU��j�t<��/�%p�^�3e'��+�Vh'
{���v�5J�(��e��ߘ�"N��7���h�WK�y_�|:��{���s1��X�Y��G���	?4����tA7�-������Z.���Ƴ�eN�_�m+t��:��-�xT*�A��yEt��-j��c�Y��Z@b�R�L��zVg	A@}��'O_y����)b ���ᚾp�RX������l�T(��U.h*�I�Y�R���f{-��~-���.$2x�Y�X�:�M]~K�9��-g����r�}>�;���X��� ��o\�nGF-;��ģu�^��us������8�,���"��؃�8����B���'�{��~��?V��~�
N�U!�*u����D�a�<���>�p��Fd�8��O2��1M����~��[���S�c7q�i��}�Ɖ���ѐ!5 k@����;�uM��Lsئu��r�ȵH~���%�j̾�O�Ͻ.6����g��B~���h!0Z���_]ԲњRYe):=(��!MTKG�aH ��U�6`ȂU��j��j�<��Cf���	?,Y��ą�n=?r��������������!k��C�� �F��&�ff���. ��w�x�.,2\�>D�!aNT
Jrn�)s��&Y;�8zx�x�;y�8:;��[�ٚx8[�;��p��v�����������9�Qýǎ?fd����n���c���������swsSW�w^Ǘ��/O�%���KH�%�D�`)�D�	�-������C��'�\����g���5�������Xl��
"D��C@ݨ�����1���u1fX'k=#]K}s]3m#mu}}#K+��+��n����Y|ᣈ�7	ŉ�<S��s4,g��?q�&�Q�F��j��mEE��@��٭F�(����A��g��vl(��փߤW>M(|��(6)477��$���YCI��%��������
F!�+<�2˟�gx-��<DXJ��0ߐ!�����.&Q
j��<�XY�����k(�v���"�&K{e�76}ll�����Q��������j�_�U�7��'� �VC|o�DH]��u"��/�y ��!�!���������;�	i�G�z-kEJ�\'Rۃ�@��:� 4^Ok�F&��b�Y4<��.�l<�[�Bk� ��ٶ����l�OOa�#�Q�ݍ�t&z'	��;��v9L�@!�o?|�븊z!ZS�"�q�����kʹ�@����V�h�'�*z��A`v��!��DV��RFk����=8N_9�o�K'Ǥ74�Ur���I��2��<fW}2nž�>�u�ͥ�!�$���#w�E�W�y�E<�>�Kl�ɢ,�u����r��rq��'쐷��J��K��P<�o��j*`��1���OZw�����Y{�����V��tv��N$4�����3w�����ì�"���C��,����O���'o�p�UVC����e���-Yu�VY��6�����6�{`�QֲZ�-�T�(��I���40d��ti=����Z�h�J��I.�&����+p��9u��^$����%����2�ڝgN]yz��݇��8���02����WWWG�z�ѫO�TSS_G��u��������{O^����@���(iy%�g�;a���������������#�������b����w/޻|b�������H/��ޣ}}�G��N=a��@_OH�#]��F:G<�E*N/Lx�f�w��^{�R�\��KJ/"������D�D���ļ��P��"�/'dTN��@SWk������ZV�1i�/OGU���f��/����V�a�v&�N�&&&6F��z����Xeu}3�).���+x�X�.��ELQzQӑ�����_su��{k6�����E3+k+g�I�@�����"|�\�_]B�(��+m� R�+����%����NI�Om{�P�b��1s�pX�z���rvQcs�Nӕ4iE��G�(� D2��ʩd4��xRNE2�}���koKN>�8�4���R�ܛ�����P���מ�9�x�5�ċ���+a	���o	��՜{G8Vs�=AF��p���*9g�+O�+=��r\��Xҕ8���S!�3�u"���75�^�^��~�p0���;҉Pҥ��w����%���$i�^���E�4��Ŭe�a;8R~%1�H�2���h�2;h�N�V�!��&���h�ӥ �!ep�9➳W�8�8}�v�Q3f���V.���*��$��)��k�K"����RK���)��á-��xk�������	�d8p�ͺCw����A �2;�L��}v#��m����k��kٟkX��̏%�d��+�����Z���B��?<f��O��yH�` /�&��jxm� 2܎_ɫas��jNG)UJn�\#���UҢr�d�@Q����şKH͂�ނT�{
kZ+�D�"�S^J� �H~���Q
���a��]��%�oE�q=��Վ~vF��z��k����7�̂?D�^KﬥwCj/#IAr��������%�W�y�ij9�kvC׊�wǯ8�9q���
� �b�����:{{˞� B[{/C+e5eEE%%ey�#Cs+'G7w�a��?}�&ad�������K&N�ei�`iggko������6�������T��ޭũQ9qoA�~^���v���>^���|����q��v�n�b�?����KE���G�o3�������q��1���ܺ�BR�����2~�-���g�'�}��|ܔ��5�u�u�^?�����E;����_�����h(�3Q�D���ٰjꦵ��^>����P��@�
�o��5��6�S�5P�0���7w_t�m:ZN�����QH4��s�'e8~A9	D�51P��/"4����p���W���"|W�o��}�iL|9��|��O=�)xS�Kj*e����%h�����Ʉ}�_��.��VT/)%7�(M�dq%YXIAg{� ����
���.$�Khٵ��`���)&~w�F����}S���A�#@�#l�c��A�&<B7�1���#@�C ;���{�є�C`���C�m�ُ�f=����d�s����'>6��
��Xs�c�ia��5�k�3
xk��k��y�mTV?�Γ���:���"��@#�J�� `х��K�bS+�M��qh|9B�D�kb�yBQKa)>.%;�W�@��q���X<2�����Q�$
�L�P�\*e:�=ڂn��it��B�7�h�_�:���R�؉;�RU��&���u��'�n%�hȶ��JZ:;� aґ��O ��l�v��d��
������ƛ�*H�K#���������Ct�#5���_�����qQ�Ch�U��ĭ_jE4NwF^mn1��V�|� t��jo=�KԌ�6��5�x.����^]ˬ��3�M�z&�-ap%d:>)�%Ba�g�G�
MH��VSDbJd�2M��ag=����N�#9��=z�]|!�AD�Yۯ�l��vֶ�����_/�~.���|ǩ�{�n;pn��c�.#�"T����Wf���򝇻�������NF�K�HȈHʊLΎM��Dhn�`ackmkcoo���d�ձ�1sw0t�l]I&������\������������a����a^��N&.�XK�����Ë���U���k�����zz���ꃘ,T�)9u��K�Ж2優�ʲ�o�E�����"̯@EXXF�̫�<m���������cb_ܾs�o��������**2*��&�;��>���>FKEOI����i+�E�Qu2p�}#8�uZ�����]����%����$��h"4!���)PV���������7p*$�9+8_`�>�ILqD�VX��������X�yS���m[�E6��V�����.����C�e��>yͶ�w
��%$iq���")��B"� ���Z%�",����OS6Fiy]��ya��=6Imt��hE�7R���������(Ţ��V�R.#T9�r ,CUCT�ީ�6.Dq�+Հ`�ɑ����&�iO�R�:&R30P��5>32	32Eqd��O�����|�.�PHu���k'��hK���*���H4�F*��R��� �*!�K�BK+�(gH�@fZ^������-`;���!��b��l!XpH�rݒ),�JaA�����"�F�T=���H��4"y�޳��cV]�w�Z�/FO�Hf#46�~��hbUu��p�p�Ȏ��܍��:���II����v�n	���YdN�̂����R2M�*�l�����j
�@�u�����WTF������ҏ��V*�������4�"E�lBM�w�4#dZWw�ݏ�[>֑�5�����g	%��:fQ�������t&�}��+Pȏ��Ҙb�%?E(s�\��PXbnB8���M"r��{o�˟��Dt��9��G��I���@1��č�˷�r���]ǜ��m��u,�U5��T�D(��WQSM�5455�U��1)��"�'����i�O�6����\e"�wqr����67r�1�1�g݂)���hc�mabhiin�`k�lk�`�do�`���б6Q7��؛�]>�m�Ya�l_������s��+��3��3� |RA�OU�|�>�[���_�����6�/ς`A #�d��٪ZZ�X��#<<M����-5��5�0Zʊ2*몫�����TM�ia�yL	r�xi`0������2�P_{0b�@���fgT=O,�ʮO�m=����q��r^|Z�%��M��5T@xJJJ*JJ�v�@��*��6�V>c�.[���=N#�N]q�mF��ؕ�V�~W��&�n9lœ�Zxh� ߕVْVٔQ)��8i����o����˄|Ok���d��[EaVQ���2��N��U|4���XcL��h�ŀ$̸�	�S2T&g`�c1>ᘑ�1>�(�"1�Q��q(��(c0c1	�q��q��20��	�SĨƪ�D% F�/\yL���d퉩:�24�R����5�e��F$kaFfaF�h�)0���<b���Hi���A}���6J��Yj�]VH��Ff��O������~�����#�e�{X�n9�>�htAC�C�wQE=����֏���:ag��[>iT����V�n�c���|��f@b��'6B%$��H�|��7���ds��	z��5�n�#���<1oٞ��N\��""��������)��
0�?U�% ���ڂq�YRO���-M�߉��/��k��.Y�.�g��Nk-�axEA':o0��"�-�a�:PI���&����)�~���$�Cg*��6�_�¯B�@�6���_Xm_КOn��+ �������l����.�
�����"�$��Wjh"*��'�d	��)L��A�����K�*!HD���e����\f"<u?1`�A�;�y�J��(��"�w��ꝧ���"�;��}�������������>NU�1�jX]=3c3O���~�D�gD&�D&���e��[:a�\3G3+kk[;''t�R[+������Dc����`�`�okifmmic�������\��T��H��"��*�b�]�\L�\��MLܼF���0*�A�U��U5�����/���"�]�R�M�r
JQ�r��O�������ia�kl�������@擋PKY�o"�'Bu��:FG����U��*��ʪXU5CM���P"4t�s#$D�^�6����v��S�ə��ZNq�kn"����������#CKM]]IE[C���������9K�MY����bC�) �М�cwb���\{Q:bҁG��YM�9�w�����q8ו�kK+oJ*��0����cK�=��S@����N.�'3�B|c�'��c�w�я5�C ����:lb�ڴ�ii���00�1�P&'`�$b�&�LO��b���'�b�� � 4*�WU��9v�1!J��U���N�֝�71^;0VyT��_�V@�023<B;(3��ZcbM�E:����OB��26�40?R�H9�K�l"T�{-�{�+����Hd}�A 2?�xZ�ߨ��U3��)���=@�~$�?Ur*��[b3R��/�}@[c
P*q|�*��J^�m�I�.i�(�oɫir�R9�5Ҝڦ!r�s�֬����5��RӉ;��E�Oi��TfW�`���w Ţϥ�ϵ�Hm+:�Q��=蛐*�@�J���Uԇp�<�� �l������T�zqܞ
^?N�A֧�:���C9��Ioh��bVW��(�J�|)�w�4!ɷJ�t�P� 
�s1�k1�{)�{)c}�����
�ɣ��QZ��@.��(��І�6�[��ЂP�r�6�jB���$_�4�?�g���H�C-E��D�Å�6!���ۄ�9_�.���}��!���W�\� �/�����M��/�e��?A����n�a�Q�]=|uuM��t����u�� -�gT�%l164�5�D������rJ��[8u��������������������!�DK�PU.B%GS-+#G[Kt�[ȎV�6��V6�Vf����J�zJ B'#57S=s#[+gO��7���UG�פ��*B|na�W��o�.)�M�D 5�$p�,eu��ZXC5]��
���lm��"�R�z5u�0
�50���:Ft���/"�3T�44¨����?���-L�"466652664LPL���Z:pMjk�h��6nʜ�K�O���e�R��Ob�_�⃖��[{�e��͇ۚ���>��~�~<j�䃚V3S�;S+��+��q���p^nM�`e����J���į ˺�S8
���
�~�csB{t�����Gb�G`��+�Wx���Fi�[�)!��ުL(�x�<���׀ڜ7�����֚�Fs�k�)O5&>��@+�~�}l�}���F��3�ɸ�����ݲ���b�3˩��'<���7��d����tF����a>��昫�W�'^��r�s����җ� P^�[�B��̺���ޓ�{���<*��$����SϋN>+<� �����zRp�q��Gy?ȑs�q��'����('�{Zt�y���y���zWq�m��'�{�e~��u��7��BJ��+=Zv6������!%���N�(8�4������3����w7K��{Y��g��A��{�W�W��a��`���u�q�Wo�]��~����j�ݬ�q!ƹ��7qKn����7�L��s����+/��W��>~��٫��m?[��Ϻ���l�q�f���g�לIZu*f���gBW�����U�]r&l�ո�{/?�Xx���S�k/E��>����Wb�]����~����'����=ʑй���92�P��}�g�}6��kx���w�%g^�w��z}��;A;n��ze��Svޞ�����wf�;c��Y{�ʙ��60o��)Kw�<|�!��{��&@V��BfI��)BFGu}W�4��/��,� ����]AЂ��^e'��,F������BrB��ӳx��%��>ve���.��.n����F涶�6�V���M�-��,�L���P���V�Q��Q��!ڏD8i�p�������\���<l--���A�F�0�����5*B[;k[t�aG'kW'gsO]%S%+}[����������	��������w)���ɨ��$aEu-�@����� �E������sK���<��W1~�,5-������������l&U�������������������ʆ:�Xc �EB!:Ě�
|����4��L@�so��L�x�X�>�&&��?���#q��rA|j�%+��,t��4T��,�KCt�Q+sK9�F&`G�����nq�]"|U�,���s���Jۑ�Fm;��0��75�I����������R�u'ߥ+�]�D<���,B-�(�����(��*A11�7ꩦ_��ha&(Dq�k����O��>�|����Dpә��S1-'�$��E���'�����d�ɢs)�i�+���)���[)⻩�)"�a��Y�PΓd�ä�۱����ϳ:�f�?�m{��|'A� Q�4��Yj��ޝh��̦[�;I�G�W�ܰ|nj������ڏ6٠�W���V��xn4��h���u���R;����7���f��ո�r,���1[嘏�b96��2��$`��?���a�6��n��N�o�������}Vj����]g8n�I�f��;̦��z�n�;��f�q�y�i�a�Y�\gs�qt��'�f�B��O8�9�<����3�8κ�8�ì�s�[��o�[�y�lg޶]��u}��?"��'�N�4rk�ϖp�K��9-|� �jʵ��b&n���|)h՛����z�;'l�����F/~>j��y���w�}�m�1�����\x�e�1�y�=�_4��8�����3��>����6���Z}�o�%�W�n�6n���M7�7�����o��wG�����Ϻޫ/[y�w�u�-�=���_ܗ������~[n�ʘ�7�vܚ�ǝ�;�N��pƾG���>�2������MX=i�v"E��v��[P2��*��
RBcK���`�艫�M߼b���7�*�=���5���0�o�	K��Ԭ�wv���{N\^�a������3;[[Gwww'[kK;+G{;WgGG'��471��aDt���(�0"��N�R�ʦ�Dhb�hj&�3:l����)V�DG�HS�LK���h�'!:��#:�����������������V��bm��`��fn�lajgm���w�ỷ)U��9��r~��TQ���w��]~)��W%�ur�W�2��<|cg�i�X]_���N	D��h�j��k�buLusCmSs3�����DU����\��Zj B��������=����K����/|�R�ɹ����r���='_[gs{[';3K3{{[����dk8�X�L�����h"��t��ٛ�G-�:Lz����K�y����ᥧ�����Tc����`�g��Sq�T�8�R�7{���<�7Ǩ �m���h����%���E�#�4l;�P}L���;��o0���Ύ,C�8H=a�a�:�w|�7|�|�'B�g	���>V������4u�I;���6 'l������~,��p\�A*xH��s���L�V!��&�o���Z�wQ��"���9����zz{���֍#����6>����2��>P���c}/e#(,��3<,a!�L����2��3�VYH����>r`�%�/%�Oe�y��|�<�|ޗB.��	�G�@����G�g#�,xC/� ��oŜAJ�h�# +C���o�&�~PM�VMC�d�
|x����,eoI~4�X�s�<K9��w�ˇE�X�����\��^�C
�H��A
�2D߁b��R!Z�+"$O��Ń|/����� ;���Ic��A�����`A�)�6
����0�a�֒���FV��Mb��3{��5�~<��s���μ6|��t(p��s�.�[����n#��<=\����rwssqpsq�ps��5����YD��C�¢R@��q��2��)�@FA��Y�U�,,���F�����9;8Z�����Mu���Ԭ4m�ulM�-L��&V��6V�a3G[S'[cg;SKmK#+U��������������0��ϣ��+A�I٤�<JnaCQICye].�s�!������'��O��"�_�avQ�SX�W�OK+��,�>m��������6FO�5� ���POK]_[�HW�XO��@����d��8$Bme������"V��P[_U]�H�"H�r�����9 d�����Npx��?�.Y}x��e#�,l��mlm�ml g{؆�����������?E�2�|憣A���I���g_{��3�ul;��z�"���|��_.B�/"�w�a	�%����Ցƽ���2������xr���"6zS�����������'K�Q=G\��ӝ�a�HP+��9@�@���P��C�Dn��u���J̩�R�҆qC����O�rYT����ـ������Kj��z��e
����^I�J�j����8�W��B�w����n<�9�s5�+����&֫��� <����'�Q�س��]��7_~�	?�fv˻���V+��]��-�t�s:ql�*V'�#��8 �B�}��O �T���:zdV/:<�|�h6:�j5�(@� m�#���L��J�O(�5��Y- ��~L~���%0���nX����})g}pL�n�b��B?,�y�=�k�]DVO�K%�[�{�+�|���7Jq�8AN�S��+e�¯ep�#�<x?U�.� <��E����R>r�~��{�Q�m!��+K��1�e=����0����w��^��o�܂Dn;:������w���3W/�z�u�o�q BO���܇{�{�=ܝa	R�5|İ�#�����.n���W��G��E(K���RQ�r+��Zfi�fk����=�/��w��������������������:����TD�k��h���ȫ�4M��5M+u+}5;#MWk��Ç����0l��׉�!����26�������[����˿�p0�	x<3=�4hܴQ�������0�Jh"��!���,\M��U��R�ꪣ��(�``i��(�����RE����8l���ԋ��De�N.K+��lH�a&g3��W���W��L3��443���tt�!�U���tDە9��L��`�I���'�U?�+y�Q�^�OO��G�R�S	�GQE ���x���?����+��]�#�N<�<�~@���K��I��G�
�hB�}�ym��E�I�uj�� $5HI� ��Bil��[�p!Om��[�n�L8m�g.*[Be��a.���i� ԋ|�$���T�oB�(�%t��� !��Ǣp9�Dp!U&B
GԈ�PR��؃m(��q&;���ޛ��s���4�v�g�Bpl�w�h=�s%�D�@s$�E��1(�Vy[D9�44q�B��C������>�!d�ɎF9u���ᵞ�+C������Ѧ���p��%d�E֣��.�C����'T) �D����x��ҕ|����[��_��	O!3[�6��Nbv6���m7�@�M^�C�?������P����h��_�>���CE�7o��Kev�M Q��!�|F.B�US9�	z'��e��k���Q{��!�?~��٫W�<ݾ��H��0���<����<��D���R�Z$����pv�VR�D�hÚ�h�����jk��E��p��^.������/"�@�ֆ BkC-7;����͞���;�^H������ƄlrF>���R�E����ssqK�Y�z�hi�3	*`~V�j�(�)a�1e��"�a;HQW]���,�ŝ����ڕP�Q���3"`��ٔS��De����Ge�r��
(��Xx��9k�B#K3-}mk�!<M�;��O��d����u�&<O(�,$�H�z�V�Y�U_J��'%W����L� ���U� ������]iT�!Y �z�~��c��$��WTF���U�F? D���ˢ�����:&����YM�S�ȩ'	dl%շ���)TR��Ao�dP:��N&��A� ��6�^vf�enXtzX�^"��j�<Y�dՊ�5"��z؇'��\x.z���mF��c���ILQ�;�ت;b�N���y砮"��$�h�H�n�h�B�D�4R� ��Dփ�J��<�����Gerd���ŕ�WSHc�it�8eTz _�)���ⶠ�dH &W����P�"_'�����!߿�Pp�!dG����d���#��s�l���'?>�`{���vpQ"�^F��ȷ�&��I��5��*��#wSG��O���� �!z� s��j������HQ2��� \�Բ: ��h.&�9Mu��<z�ҍ{ ޣ\��ܜ!z6l�0�Az���!�9��}&t;94&=<.�G"DE��3e�ҹV��WU�6627547�32�50�bM�zFz�f�����)���������������������v�4Ա2д�CE�no=}��+78�]��؊����l�6�W6������DXY/!�)DkG�2S���NY�v�����
(!O]YACEQ6+�"�?�
eD�Ճ��*5��:%������PU�t(:�Vc&��m5����G1!y��s"3Kc�*c3pqYeI9%)9y�.5�����2�2wqu�ݟ@quD������������7p���,�"ԱzS�.��Q,:7op:���9u��"JB+��#W`e����b��",%�J) \XBb��y�¶DW����몣�k����6����t&B�tSX|2[�����Q����FGh#K+���x����D$7)�jS-M�ߙ!EG�d�ԲZ��<h��Ur��n�����D�tշt�H%x/�D������bF����ڦ�:��A�A�����u�ǥ����K���,�M�m����(���P6�9$��N�E�1�����e�p��\<L� U����=Q������BO$招x��!���D�S�P*5	�"�T(nK�%�6��ڛ[�~e��������"C���oǇ��[d��d��dG�q'O��ᵢ�R�B��U��?��&)�?������G�CA�$2�*Y_�I񙽷��C���Ǻɡ����Q>8:,�܈���� �t�ёc�j�:�;�.*�����z:���s'�^����ν�\݇99��Zٻ:����.��11��'�DOO{;gg'�[���'~�0� *�(F&B�2yƒ����YY8YY:�X8��M͍��M��-M��\�,�� OW��^.ý]G�@
�����d���@��a��jg��hflka�l�Z��gqOb�_�V��o���a.)-;61}�ҕ����X�|��d�&�� ������4��bu�u͌�d�et��5LuT���4e.TSB'�a��	��k)�x��umf�{�86�mzfHZfxFATFqlfi\vQRnAJnΔ93��_������Fw7'g'7'Gp������5�����g��ێL]�D�m�8�H.�I�7i��<*�ܚ���_E���g�߬5O��Y��2��Fn����~�^���	U߇�>�j>a�ߨ���'��#@�R�C��bXi~ʯo�/�U4G��E�wĖ�q��x\[Be{Ru[Ju{
�5�؞B�����5����Db/�@莭�N��&�;+����E�tKm�G�3<�E�m.�M��m�0$G�͏ʗ$7��7�Eu\ȵUɯ"��%׷���0�G�@�a���#��¦fqs���Y��E"n	�A0(�&�>��d�d��eHy���;HD�&)\��"w��ֶ!$-�C�{����d�PZ2x�����. �:�@�/ȷ4u�A
�>�D�܄"_��o�o�5sd[�}�o��&?���[(E]ȀGB���m���ː��2��O�_~8T����-g}9p'y��=8jw=�2�Ć���վ�.�@�C���ˀ/*\��,(��	�"�"��ҽ'/w�;���ל�F��f��>ޞ��{���֑�����8;�����˛�>{�.4<�JC�a�������3mֲ��V`a9(BS+csk{3S'Kcw'��������8v��1>r�@��rqs��'Bt�z#mWÑNv�ܜ�����l�ǜ��,��e\�(?DX��[������"�]~���j��V��Yy%)y>����u����0����X5p$<-ee-�ŗ�d�/"�U0��kb��&�*&�Z�n�:֦�֦�Fޣ�Lَ��u�i̳�̷�!���3r#�b3���r�Rr�&L�j�l�c�+�����������l�fV��NN#�Lذ���Ż@�Z��~�0��Uz��̪�\��<�������x=�����d��k�ٵ|�9��9��8J	���@M����TX��Fg�9�W*>�*>�
#������SYB�u
[Y�^2�ˣ�کk�i{mSp�et� �	v<��`�cÉO �ɏM'?�������r�St9��t�i��i��.*���W��E[X�Vp��V��{��E�����z���D�}�S�n��]O��猪T�&u"�f���Ne'�Ki�����0�"��Z�)�Y,h�J:�[���{::z;e��u7�t���D��(r� �6!J��'�-m|����[�T���#�������-�b���L- ��M�<9�����|�_��tːAeO�y��V({3RY�G����iK�@���H��ܤ�߶�9(6c�Fi� ��������������T���*i=�y�1��Y�����p{j�h��6z�5"�IVg�$K��{���Z���t��.�L��r?���׻�srutt6�7��Ն�;{�K��W����5�������}�e��� <&#">G~�0>�8>�0%�l�U�g-qp�C�v6�66�v�����hKQc+M'ww��]G�t1�c�pWw7';K��&N����&.VF蔄�F�vֆ��&��F���n�N�
�$�"�c����_ʿ�p��De~Qerz���s0jj����,���ao`c�i��n��������Q^)*k2��,�����Pc���2�Y�X��aM�t��Tl]=A��/<��e�MKK����ϛ��媥�����������N���,�	�BG�E�29z���-��䋊�Ql�ܺ�Q�O�p`�י�i%���
j"K�+��Ռt"/!3w���B8�dTҋمdz��-�k�������{OyT��O��O4����+	RׁЩ���ny�DC���s��|�k5��Ѳ�F�#Ƅ+D*�+�W	
S�^uB�Ƅ0�4&�E��	�ǿ�zk:>�"����t�����>��r��`_���e��7:����z����p�S��-�߶y���I&BtLQ��,q5a2�Ck4*�Fv?��D��b>[��Jy� ʍ%mr���!�[yr��� ��N��"��w�g�v��fP9p���������K�m���V����wK!���Z����A��M-@҂�H��M&ȿ�p�py���;{��G�D�m��X�D���S�.lnt�l1�����꿉p��� �����ԅ����t��T��@�r��3{kX����g�C�C-�c-�Hmz��AA)o��քCU1:p�f�/��(h����Z���r�ԥ�σ��9���a�謯��n:���Zʚ���������320411355��C�l��Ԉ�L��Q�1i	��@FAռ�k��Xdb�`e�hmeogm8���[X�����|���yیf��lbgkdmklacbe��&��6�n���#]�x���7}��%���G3�t9v�ٻ4||>�R�+��w����C������bw]5CS��;�S�/?�o�hK[��������������������Ctd5P�Ƀ���c���N�Kc��1:��!VG�����on�e2��i����r�Ӳަf���E�Ƥ��Fg.����"TP�u
����>������Ίfg���q���Kw;�-Ҵ|�\�K���:�VT�<��Yzɫ���B�ä��d+���Y�Ϯ�ԉn}�T^/�����مr��ͬ#Ԥp>x����?���4*M�'KeT�����k�
�Em������F骣H�l��ʰ���ځ��~q��1�(�1�
c�ƅ*�`& ��Io �I�
��1S^c&�(L�T��:1Z;0Z������둄bn[9�5�D�R(�k�3��'����pՉ/������O��>��r�VA)�DX%��.���"l`��XR�Y[��K�;m( -q� �H'^K�ֹb$�����:�Z�U,��S��Oa�����]|)R
S~|I�L2B�����3��=m�}]�Ki��+iA�7	9�@���m�9-����P��h� MR�i�/�������vaS��/f��H?!�VG���MX��m�������C�"J8\!�����M��"��m��koj�a�:Dp@xi����*A-�65��ȫyE-�\q�+D�2��爐!��4��¯?���@�	��)�|>�4�a�V�C=��Jo��H��|����m��m=�vՁ[_�n:�
�Gp�%�����^'rK韎�yׅ37��~2f��#ג
I�D~7��J�!�oe�V�Vl:�u�՛��ڴ��c����UUUVUSTV�()�S�(*aT��JT���\��4L�A�ӢⲢd]�c�3���ܢ�Θ��51��u٣�O؂=��!�\0��4=%�ل�Ξ�f������ B+Kc[��V� Bc���]���&��N	���d�TȬfvn��܎L�I*�˺OȫF��w���?�Pn��⪂�JT��X+��v��],/z:c���6�D��(�a� �7�4��C��ib�u0fz�{W6�	r"��YbL�c=uC=]=}C��PK p@���HM��Dh�2����딬���Д�����Ҹ����"��s�����f9�JC�,**�ZZF��6�n~����:�-��"<M-�P�8�8��]E}_�]AΥ7��4�/&%��uBav�dܢ�ɕ�/�^��Oi̥ҙu���(���;�{J����J#s�F�`��M��-�%Aj�i�:Ca�9���=�~Us\�J X�{H�rb�"����e
X03�L��L�W�%j1>�a��n	�ZΓ��E�Q��)�c<��N�}�DU�b��cC���Z���h-gt����l�?DX���!C0�_@�@�	_��d�nY+��alA�bGo'���O�uqE��%���>t��`{[w+<������!mk�7c��6w�7�d��Ca[7*Hy���nV�6��\zQ�,�M��M����糛�D-�b8��������&�T�$"^�����Ç=}=4&TA�l�p��$��m}�_�@��xb�!�V(�Q�$6�.�B����oVA~�������Ri
X�[�A�T� �m��D���^���R��/rm�6V0>@�#�q���{�?X�����c�Y����a3�-��B��q)a����D$��X�^{�U����+F���&`��G^6�|ͯ��:���uT�m.]p��ms���w��w��k���+��`T�Q*JJZ�X,
kT6�ZjtBVtr����¤�⤬����E�6L�5_SW6e����:H�����o[S��{��''�0��y��lpQk#K+ct�mKcc3#;3##mu#eO[3rE~3��ZY�f�<7'gk�}'oF���h�YC"�]5���{�U������y�q��8!�����u��T77U������^�i�XCu��F���(�+�jjjkhi�i�BR�b^�V�r�Ȯ���p�j��hi��jC"���P����m��Wi��S�ަ䄥E���f�2�P�����@#�����������5;O�]���_$�$�=L,�~�U���ޤ�Vq���
ɱ8�Ƴ��KϬ� `A`���!)��K~-����K�dS)�tNi7����<�������y�ČV�x:&�����'�Z.ϧ�3i՝_�F�ݗ?TuMs�[�1/1c_+�U�M����2&��L|���̔����ɱ
����뎋��y��\%�)g1q\i	�5_О-pZvZa�1��/զ�a&�*Lz��Ng1>B����]!x!R�h�5���= B*�"d�� B>��RI3(�I�^\�&�#��߆��[<��cu��E����UT����=���4�� �u[6�Z`�����ӧ��n��%�Օ��?/]�!56�io���k6�_�iÜ��Zq��q�������ٓ1A�F����������j�����\����,��:0r��ѷ�]�wz�7����<w�lOoWo_w���Ș�]�w�
y]Km�t�
[��O�$|��9,�:[ʪ�W�_�|効�8u�Lm�/^<۰qݖ-[֭[�x��Zb�D������liA�7���M.BAS+�'�ϼ(����W��oR�4���9O�η\�c4r�)�f�O�"p3�-��ڶ�����B����K�$����:����<N�,�s�9p��j)B�C��59O��4����ص�ߘ:���_���Ek�Y�m��u���@��j��j�
*�%������爇�_���I� b�r�R�����ũ9��_Ehlhhhd�575��0�������xabH�;s�y;�[XY�Y�����aM�:fzZ�
-ՙ�~�	��Һ����f�C�9z�;uD��K��V��E���S�U��^�W��#�Y�V�j��&.۳w���Asgz�(c4Q�3+A4�PG;�jkB.��5mE���N��{aӒin.V�Z�x��
���jk��k��hc5�F�̾�<�i|��]r^xJQdJi\:��B�}b��Y��꺚hը������QT��'��͌��}Ʈ�vD�6f��aL���ݨb�)E�E{n?H ^y[���}�=����ݘ̺�lt��	�����U��d�7fPyɔ�Xb2���{�G*��*�U�f���T�4���gt������T-�U�I�Q.��ЋD�4ǝR�xGe�=��G���Q�c��A�1� ���Ԃ�"0�1c#�c���,�=L�F�Z�!Nܝ�H J~�U�]՜�^eJ���h��q��Rt�ƙ�}c9�JDakR9:{���/"
"�,�M���� qsO,<{�<FI���W�+p��������G�c[���D{�d0����Ϛ77p����iSoݿKe2�Gf�8e�3���k�oE����O[�%g��o���\����ى.o߼5|ذ��Ԙ�hS#JmC�@��J���kjj��Չ�����y����7ޫ�4�]x��)�Ƃq[�N�w�߻��!|
�QB��СCcǎ=�|pp��˗I�R�����������?E��@,����Q�z�S�5|���VB�h�%4���4�4�:�o�w��=&�ɠ~��b��[u;.�,�R�GElǮ�s�E��Ke#2g��;/
�<�|㱥���Y���i����� D������A]�(�*���zzXC����)&Q6oz~BVQJv	�SR�d����a����z�X��D������x��@;]�,?��ֺ~���F`Ac��1��Pms��a���`j0��:h�������<����������ۡ�eI� ��\Z~������X~᳷aE����o�kG���b;0�X��V�����NKGK�}�QW�h()�Z�8�F�R3�R2��Xhb,5Х-VUGE6g�����&$B!�DM��f8��y��I���S
�"�N-&f�Ыȼ�ɳfY�Z�i���P.¡DoOMW�������q�����=Ʈ԰�2�8�<M�z�3a֣7��k�)����6~���U�Ͼ�$vfִf�4�x�Ll̫�W	�iu�|�@D��滵����c�<V��<!B50Eu\�r@�R�+�'
/nB���ND�	IJSR��a!�{B4f^ј~O1�B�+T������p������p 3AFP�?L}\���wK�dg���#~K���\�_҄L?�7�Ƅ����)O�Q���<>U#0]/ V����M!��Hcs���R��?J[ ��@&B�� BpvΎ�'M��`>]}�*<���'��:{��
�\���y�����!G�+���B@|�����Y�:�T2��8\6le�;z�X�<u*O(���G߉T*�$B���o�;ZZ��e�����E(�8�Qv��M_��֚��VVW�����m���bS�l�����L�6���s�]���YL�o>55�ȑ#;�n����
����,����[�Z�� Bq[[SGW"id��i��#��o�m7�;p� B�q�"�m��
�W�}�E���V��o���W?5�>?jγt*���>r���*�Fx����i���>���@"���I���#�SN�Y�qϥ����zx����^Ffֺ�XmmM]YcE--5�4L�X]==�atr^lza\F1�B ��n���Z�8���X`��̌��-�ܬ��1f�+5����0[������9`afdabha�g�ձ6ҷ3ѷ5в�Sr2P�0�ng���b��~�ҽWQ��"���H�y��"�]�K�U�/�"p���
p���b���"+WUm=]C��������������
���~�Zj���������������,MT��P_ʪF5�z:?������ӌ�ϒ�����Ss��r�g̝"D[�j�B��O��Q�5��:X�f��3`�����̚�)ՓW���vh=�`柏k�$�OZ~g��1�O_|V�I��&�g[s	��
K�o�����X�:�܏d���m�:�)��H�Xu�p���x��T��d�q�U��M�:�dr� �b5r��\J�VC�3�R��B�׾��B�)�_���`A9��\�4>@]�2)�pv�ָ]�;#�%�Ou�%��3��F�d0��g�)O
S��8!Uy\�f@6vl�E���O��D���j�!V�{�5�6?H���"��oD.o=ub��#F�������X|���g��w���A����%9q|�e�,asG[Y�D(��Bx���&�!#���zF��B�� �X��px<x�ۓ�e���VZ%M��=���\ڕ���w��g���n���	��A��"�������y�p隕�Ұ�H[G�Kkk��M"��nݺ}�V�������6�?��������͗J����D(!���&�F��D�h] B���^$��m�ͽ;.����ND.2j����#�jF̹X-BN=kp�z��	a~B���q��-�$,�wV�!#�K�_��肕;�o�3i�#s{cs[p�X]#c}C-�����.`��H�65���=��脜��ed"�N��y��M[��?5:鮕:��������������&����k؛�Z�YY�-a��2cf�4Գ�ײ�S���)BoWW����%�F���!�~�/��08"D��_�]�t��ERV���1�Vv�F�z���F���к������������������������������ F��XU�D����Xp�?�0$5?457"�8:���Ⴅ�\�͌tt�lЎ����TN{6�掮�#��[�ǌe��ǯӶ	|�Z�,�\�:P�|���^����#7�R1Y1o�S��SW]̩�ʩ�ȫiɫi?�`xZc�����G#q$��ȓ�x�u�WJc�+=U��Tm�k��1���ǧ�M�V	z.�ws������zA)��D��Sz2[>D�~z+D���.x�:�Z)-�/"D]�5)�j~��o����t�纎ODq{�Y��T����Gx��a����J߃Ƨ)����k06�s���/�ܶ*����G�����w�b
�"d	E��IV~Z���Hp�ϳ��c�����b����	�ӧO������D��?|I�����6�ۼ	���ww����_E�.e��KW�X�aݝ��A�
�*iY�`D V��&�3�r��� �ǃ��$j��x\%���M����ԉ��\�+�`,ح����#hXE[#<.��F��4p��]�qc�Mb�Hk`j|����׮N�<i�'O�422ڹs��իׯ_�_E������'li����a�\�U�2�[6�j3��[EG�|�F�5�����f{O�]�V�F"
[����������^�FQo�
��ם�6�\{�vj��ۃ�Ȱ����Iٶ�ʊ��6�8:k�*+{w[;Ws+3s+k�:0���	 ��ke���5FƤ��#�L��!����򈤬-{����������������������Y�P��P��@,h����U�1ѓ�P��*Bw3]o{��nnVvnn����'P�����~�>�[���?�� �G2
���ٹyk`�U��zf�ʺ�}T0�*�5Ԕ�����Bu-3u-5t)���":��:m�P�PY�HD�c3�����Yo��C3�'��Pĥ�$������.Z�����������������oX��`�M��L=|A�����F�:�]~�����K�UE�^zV����x(a��7��Ϻ��9j�n�`N�|�����G�Sk��dJ�����,:R�?������oǿV��\y�+�I�PN�C�(ǿ�8_Q���#,�n��5PI�'���)_ҙ�ڝ"��Bf��0��Bm�L`(Z/*���P%Ey\��X�q1��;����+�E�|~)�)�֚�G̦�Q�H#0By|����RP��D��h��'S����R<�/��e.DEX)�N�o���t?�;$B*�"DG���'���^��w��M[������ق�ttt*++=z4v�X��J$����r�-SfL77�� ���xb�`��"ljoU�Ѿt���{w���������-�b�
+j�\������O<x0::���>���ёQ���V�S'O���V�f��2���������;z����ǎ�6��,��4�	��WgLk�%F�Dk��nݾmŪ�N.�'N��4y�ĉ	&ܻw�������ݝ]���&H��*¦�����H��D���oa�/U�2��a���DZ�Q�ĕ�_&5�?Ո����E�ch���bv_9�zX����4iVu_9���"ͫdW�ML�WJN^x���s�O]Y�e�����.��g���/�h�z;��������o"��KGG܆P��֎&唥�U K�o�w�q>�{���F�vwu��ZXk�k9�����ka�u�l����6���dX��!Z�8�{Ya�;X���L��"2<�24�
D����{��忔��0���8(¢���J9����Y%�F`M���MA��ڪ��Aet�P%U�j*�Zj�"T�6���5t��t����Uԕ�e���i*�kk�3ԣ"��np�Q���i/�3�����f��fE'$f���f��[���FXk{'{@6Q��|�v�5�1�Z��88x����b���{G�_�g�\5yٞ�K���1��T�U7�[t`Ӊ'�(�����v��W+ɫ��	�� ,��V@%��X9Q*��rO�����b@�bP�Ҥ��SިNW��61NmR��0��r|4��f�%���)�mC����;N�Q-j�����]���):S�+N|�v"�	
��(�*��BF��l2�z�)��J%�B!�X�O��l�.��^W�Z=0Fy|���(@1(3�%�}���Ʒ��bfO%@R>��lz�!V	��k[�Gm��đW�Ҹ|�PQ�/� �$�"�@!|g�޽�֭���f�
		�b�uu�as�����勄l.,���9x���E���BH~`#ȅ ���Q�R�̈́)k��T��,9> ������������C#����p���7��T*^tN۽|�r��o����:~��ŋ᧐�@�t��勻�/(-�7J~Xx���M�:Y���8wo/x3��6�x_C<r����Z��H� ��_>8��-ȃ��dgo����PGj���{���2��e^ο�YR���������pt�A�TS���j� ������Z�	��d�d��vTr�p�.yW�2^k9����V�����q�t �F!�$$ѻ��Mdzۡc�v�;{���-;1����H����������	pwusw�pw�tw�����5�j�P/�|���Ԣ�������%�vظx����0W[3Ss=3S]3c-K#����f���l�L���0"�`ab'��Z:� B-O+���Nc}|�����O��)NȪ�'~~B>��?]~��U�M�࿌��������I�����fzMEE%uE�� BH�*J
�JJ�jj��4��3V�3QGEh��f��l���UC��GG��BE�k��a��:j��Y��IO"�C���%e�OȊJ�O�(Kϫ�-�((/[�t	�����gco��rll-l-!��ُ�"��l��k����E�K�I��9��8fX6>����,ΩD哲���:^^ȯ���{46�����)�bn��k��L�	75��0TiR0 a�ڤ(X*O
W��0)m�9!X����=Q�s���� ��ӸB�"�kG\V�՛�3�)f�kL�k��`��j��ao��o��ZݏI8%��"	+_�9��[K��<P���L��L�T��	������h.����E`���΅���D��L 6��\'�%!:v�@ �T&�f�
!����@ ڿw���k`%2"r�̙J��¢�����a�X�PPUapٯ߅�Ø<H�����҂D����➁�@��:eU���.�"GXBj��(����_{�����i�@�A		IH�������Z�����Hq'H�B �uww�x�k��u�l�@i�~�=���|��������0;�\3��3p��k��{���f��j����Դ[ *�ݬ9s���MFF�ܹs/^�p�B!��NfHW �=z �h��
����*ԷDXB.�ת4�u�?�x�{��ܫ���& BzK�D����
d��e�E���-�y��p�n~$B]9���b���UJL��Z���L���m��k��
��	�-v���0;8FGo���\���4��&�ݩ�X!�U���]�x�����[��K�^�:u���u��@w��֥k�.�]{ �z��ne�Ex�N1�0���C��DS��1`���?�9�_����;����7j�$8�I�����-��i٢M��m���[��l�&:]M.���]+Թ����'.�o��>�&~��hB��"��aBEH��H}��bҭ?���Wʬ!Q�N�(<�Q�:,�Q˦>�|>l�A�4n�Ӵه ����F�6iմy`Ӗ8AM|[7iֺI��M? �n�Ӻ�t-��O :��aߑSZw�z��rj�v!�N-��Q@�h�R��ɜ��w๐�mb�;���Â�ڴ���7r��S�|�Ӛ�cf��0Dx�=!�~)����8�F��P��
�
8)%����R��T�#K�d�s�����c9I��WVk#�mh9p����&}8�:�p���h��ƣ����"�p��fc���>�z���s�Mזh_0l���G
�Ker��|��"�eЗG>w�g�Y�Q�?q���KMF\j6�R�a�M�]
u�$�Z�vSF��Ns��վ4w�~�}:�p�MT}�S@���>C���Y��Z>�\�2V��$�gRu�\��"�hQ_�o�P�uh�\�6a�����z���[����`�Ӫ��B,q��M����+�*(�Z��J����B7���Y�tɄ/'���j�֯�|��� J@���CǏ^MN�v391��d��?:��5% #�O;:\.\{U55�.�g��h�'T:��a����SF���0<2
ӗ�W�G����-�G}��W�p�00<q��G�����og��ٷL�q�A�@g1w�����oܼ��~jP��N�V�۝�$��QoA�j^r�RO�j�"�Qr4�����ޖ�2��F����ka�u �e��mv��_gj�B�U����f��
ԋйa�/��nڱ����+:w�	��a�=��8��x%�z2:4����ߡ�V%��[H�E3o<��/�کW���������h�sa�66m�D��
aTh�W�w����~��>�|�.~�w$$E	EB�K�l�/�/)z���!�7�P�	�S�鼬"
^�0� 2s)�CG}���Z@-l�ҧY��5��Ys��o��5�l�������ЯQS��w��o�,����E��>���y�߰OfEt���-�|�2;���!q�J�m�q��o��}t�0:6:�StL|����_&¾#�~7c�7Sׂ�#G^��]��^��M+Td���|sb63�H��ѩ�^��m�K�E(�#~�)���5�SuF����]�o�%-���ڍ&#Q{\��F'��� ����dlj�q�ǥ5{��������)g�'�J�n����X	.,�*����W��+��}t�g&����lą��/���y���y����U�"�u%��B�{�/�f���t=��|t��أ�<V"�X*9�j��T�B��}�Y�4~Y�>3�H��!.B��i��%B�W����ǎܿ�ٳg6����s�rbwHJ8w�}Xx�&M�����=~5[�"������P.Y�|���%L��R>q��P���bO>�:k��PM.Z�	���i��yu]-`��@uP�A��
m׶CtԑcG���+|��çO@�={�c=x��e��C���<�D����샷8w�.f��˅g᳡���8d0����S��>r$X����	o% _[�M»��`��8��އ�]�#�g���z���@�چ"4�tq��� ��.�E�,��]_�Q*-����|�杻��_��S�n���w��� v��ua�n��^} ��\L��q+��vVqZ�VF)�a./sK�3����f΍��i�:,��7m�,2�Udp@t�Ўa���Ѯ�Q��Ș���h+a��f��=��v�<���������q�6��mFCҘ|�@X@*y�~I���i(��WS�h���W�8�3Iws(=��hٱe�� _�6-[�n��.�m��|ݢI3�&����h��뇝,lҢY�_�P��4�	�E�i��J����~>���>�fIT��P��U�Vº[��*a��Eda	E@�#~?�Ȩ��6Am�C;w���)'2:��1�����v�?t꼵��� "j?")���κx��^�J+V��(�KUw��L�:��)`���R��"�Se��5v�֬R��LכD�S�6�_��d���[��bXR�ך���|�����F&�u�o��o6��dl�|�̀QWێ85�d�����tMC�t�T�E�0��۫�e�C�R�D4�D�b؅VC��NL\qJQ�p�*�1�U��j8��Y&w��W>�q�W���xT�W�M?N��u�y:��M�V�5R�s��B]��Tȴe^��es�Ay�>3���%�z�Kk���m��G������5RU�XM���y�.C�㐷6*����*�zk�_����@�����Z������eC���a��t�w_�wiP���_(��.�������wD(��_��\l^�y�������φwɍve�s� �Cf�ԏU��:u�N]��֊��v�B�_Cp B�Cc��Pi+Mj�C P*�uk��\�y�������"�оCt��n؃.q1 B̅]{t�ߏp��a}z#�N���Fm2�w�i9��<:(��!�"�f.[��wS'~?�C||Tl�N];Eu��ٳw���=���+�c���=bc�t�ҿk�ݻ��u�v�<�g��C@��3�=��_l8l^��7�ک[xǞ���v.�|�.;�P�OV��2CJe�BQQ)����sB�D^���]�YHe�ͧd��sJ��y��W���Ӹ��-��5j��,�ۢQK�&��M�[6kު�o��?м��f��4�k��Jߪ����-��~�Ʒq`�&-�ө�G_~:m��A�,�Y$M�JS���qQV^��T��o�m׾]K����x-��'*�}��p�]X��6!ᡑqq�z��p�37=30|8���S�e�K���t��Y�I����,s1�\*4S$F�LG�8�)<��a0�L����I�v�n��'�H�r��Ы-�_i9����@��$�`�d�QɍǤ4s������܈x5�b�೭?�}_�=�k*�
���bY�3r���|F�ӄފ�հ�V�.�*r<˷93�+UI�{���5p���&#RPE8&�g��K�0��qj��O��S���;E(2���6�_��{���z��#B��b���"�r�!�����ׅx��C�+4T�_�m8忇w��qi^V��3ٜ2�V�Խ�B\l^�y�m��Ђ8�K��������+B�u�jp�LW+4`"4Vawx.�(Ѐ��`
.B(��Q�����v����&����+drÚ5[�=��1o��ݻt��.�]hP����:uDb�!�5������'��Nf1�F�Φ���3r(�� �ʚ�f�W?M��'�ݺAu���v��׶]Pllx縈�a��;u��kH�>�{���	�����C���EG��k��A@#$�H�#���$%fpp���t��$<���R���3B�D�HC���T@a��/��@��/�?t���{���u��9�]H�MZ�5F"���yӖ�}A�-�[�
��G=�a]̄�� hײ1a�F�-�F�	�o4p�����?vaR�(�Tx��y���]��/敔
I�"��ˉP6nָy�f�!��< �u+���Z������l�9�s��s�n�i��!cfG��z�ԋP�Z��]�I'k���Y4c>�Zȵ���T���42��q_n�EH3����4���V�.�p;x��!7�^~h=�2"������ɭƤ4w���t߱�#�FɈ�ѵ_V����?��ʕ�pTV�S�6���X���g��'������K�i���Y{RD1�)�[��\j�gqw�|��!g�N����M���3\��7��7[y�*7���e�����
�S���"��2����=�n�E��xDhwX��*���cQ���������jˀ
��E�����i�	Ї�?�����P)"�;�*\���m��R� &�C���ոq�7E�6�g�_l?_�a~��#�����	�����L�p��9;�����@��@��(���P��U�t����C(Z;W��*��n]�r˶���^"�ֵO���fM��h�z���0	t��+&:��}��\�u#%+%-�}�NIZ.-��U@��Dt��{&Ϙݥo��]��v��e:��16�Wϸ~�;��ߧs��={��sX�^���`dH�^^���gX�P�����A=a�+.:,4,,��χ.��Y��#�*Q�дT���UAE(��I4ʓ�O	y#Ex�⵼R&��^�ӓn����n>m�̉_�P���}�l��o3��o	\�Յ��|�������߾o|��Vߢ	��o�����X�4��GN�ۮ�.f���w"�t�g���>h�.ĺ�m������6�M>����^.Z��s�;�u��KwXx���Ej�.�Dw���K7ߡa�˶��%Mi��t�c�W3�e����-?�9�u��!�/G�85�b䘄ȏ�F~|��''��ONGr���s@���EN8�yB�/�'\���R���n#��z��Ȅ��e�n��a>K*P��&�Vv,O8��ψ[>����%|8�B�Q��F��PX�4?���K�.~��S�>M~�j�F�/�f��RQ�c/�|���q�ϸ3��������M�U��N���j���j���T;�V����r��~6�ڿ7��sj��e46��fr8m�"|-�rt;��N9���3^�W�;k*\�eNp!�@xN+�'\`;0geMEUmUUmy=U0��͆j�x]�y���o��7TTU�w��mv���ry�]6/�2 �CY���x��᪴;�F�Re TjBe���㷛�o@�|�;�g�;׻�Z'O[�6>dZ^��2�OD�'b���	���m~�2>�/� �U��%�j
�n��6��mJQ�R]ݥ���)�aW��%Љ����v�_�a��=�O��#�S����F�4�Чq#4l�胦���ݯE���� a\l�o$����޾S��Q��EJ�CW�x ��`���N��1>�S��Nq1�:�w��o`ϑ�M�l����o\�tڷ�F���9���n]��ݻ B`X�������%�O|��a�蹷���[NL�41�Mh���H��F��+�&)It�����t�@,W��x��&�l��!���"<�p9���YH.�����@n5���r;�e@����:u޹{�D.����k���B�M[�l�ܷi�&�|�5j�߬}��#&	=�ک]"���5A���h�ƿm�_pDh���w��J��j.3���Q��)��JJťT��Q��	_|Ԩi�f�MQ_6�oQ�ᗉzzk�T�a�Ew���w���N����ؙ�c�%�3.�𒊕IE��)��Ͱg�\E�<q�]��@\ARUP46�VO�XG}��.�	:ahm,�c������4��Z�fT��8�n:<,w���L��jwS�n���*s�]n���q�yV�������H_2��P"S��jg����>ó|F��}�g�i�a'}��&�fu���Y������L��=pΕ�O�6w��q)>C-x�g�i�	��:�����J�?�T���
���k˄���J��+�`A��.�8�=Ֆ�̏ru�}�L��U��`��Z�5��� �Մ�}w��� ~�!��h��6�բs�e.sE����^U����8��6�ӎ.̇�[��D���ʬ�@�yǨ�)jk+��{UoPWS���~=�B�S��Kަ����rX�f��`0� Ċb�ڌ^,`���{�j��M�ĉQf1�:�C���v���B��R��T�*��2�B�딉����<�uU8Bu�@U���q��XV��Ұ3��g۫�߯;'xзѣ~����\Q����M#������ݎ1��q9O���]�~�٦�7�GΉ>uʊ	wx�����_8~f�N�v�Jؗl<8e�y˷}1yf�ν""cAu��n:��a=i�ᇾM����Z�7�=q*�f���w��C��9�x�SL��BO��C��4�M���q�1q�P��Eu�;|h�a��vm��\;{j�ѡ��wҳ���ַ��~�F�;jP��]�;�3�g��S��T!)k�ן�o�&4<z妽W��o���Z
���x=�+�(Ԙ�����D^������C�fQ�h������|$B��񝻜M8�d2�?�!�E�����4m�D�ʯ�_��X���ۇ��G�9��.g��8�="(,�]2�ײMpPx�Pt_��E�N/栋���R$T����|����!m�4oҢes��.@��A-�;����p���_�����i!�ǟN�&���h'3FO�|1_}�P{�_��`��_��ڞ0s�)����uR�:����6��1T�5v��lĴV2��tg�YAwUR\G9��tT0�e4��nt���|[%��V���gq��N0�J含�E���Y�z��5w��[s(�f������v֧ߞ��g�%i�֗Bs�RG3?�:ݷ�Nߝk:�P��?���k�>��d<Xs�Ϡ9>�~�{�J7��Z��U|=.B�����,(P�`���.Ԕ�s�uA�A�6��B��-�t�6Yl�2(]�J���&��h���j1��&��`�j�j�^e0j�v��e���0���Έ^�f#��!���2��1`�e����Yo4i�z�^����Ǩי�:+Bk7��0����@��0�Nk��z�Ao�o�|�b����j4��L����N���pՕ�?�R�T)�H��T�j���k�w���#B�����ᙞ3��Rn���7~Ŭ��I̲QӶ��q�cw���g���7h֞��Τ��O��v}Ѯ�O��#��s��&o���$]���Y�o	$����O�=�4g�7�6�4��_N����t~��Hv?B�%)�w� �m�!�#������",��]r'�z���K�0��N9�pҔ�ۆG��ƠD�D����>�G\d��D�NA�J�n��=b:������ �:�ݿk��/�g_?_����D_��%�Ch���6�M�dd�
�z*����B���*5$�������"<r&D�+a�sJ�5��zD���ǧi|�nl.G&����\�dA��6����·���� -��Be��?.�M��m�ɵA^ҙ�=;���r�U�Vmڴi�nf�
rH�<���$)�(�"��I!mC��l֪U��(®�};}ٸ�t6%��gg�W
$	�����n�뫕Ӯ�Lw���&����/�����PG1���4�y�7+�Eh�],�av��(F;�d/5� ��Z���6�H3 �F'�ڬ�БU���mFm��B���U����-�p/���A�]͆$}8����S?����D���=�]ȵ��֧|s�F���v���&��-�]h16�~�l?��O���`w��LT����BN�+@uBM�@]&P;�*�@mǇ ��)���V����]�zL�w�6��&��U&��^m�V��ej�C��`f�UF��d��B�`Dew�tVt=>H�Q�*�]ep"�ejC��Tb�k�Z,ߥ��dj�X�)�"����z��(��1��>������%(�b��W�s�gx��C��� �6���{�Q�J_�ԕ+4e/Y`���)�n�+6X��1���Z'Wm�h*��g\�{[#b�"��J)p����%���k�G��eֶ˲{n��UǑK:�\6g�A��auO\r��-���צ�9'-w+kܷ��>�$���j���P��L�|�o��˟�����GN�ӽ�H?�o#�=���"ff䢻/e���|[L�K���"�����зg����m��2����^<�/�w�ԫ�����=�t�ܿ[' Z@�� ���6�F=�o��MR��
��۷Sl�����U����p�qQ����s�v���i��$*B"o�?�#-��7 D�e����̛��w_|�q+�F�� �yD�����ޥ��^6/�r���Gw�X6�밠���|�����۵k׺M���A�Cp&f�A�Yd!jc]*���J����]۰v-Z�l��5��G�b�~��E����g��1~6~Z��߶����L��"��������i?g�dJv�|�W���z���)#��Y6#Y����4�����iLL�`�,������f�Te��R4�����Y'�:;G�D�DN��)���:�T����%�?�&��Bw��/�?�70�wpR�a�͇���6����w����G<S-�|�ayr�b�ܧ��֟{2p���1�[�9��~�s����EC1�c�� B]���?p!�
�P���G�%gHj��/=�Q�Q���g�#�����ax�6<��	�O ��!�� o|�E}��iȆ�L�|K��>���oz�7=E���Y4�c����{�,6'�l�����Y��x�� �����/���w|�}��o�*�R<�3��1G��	W��1�������g����������H�<�螀�X ���a��z7�v��90���+"��1eo��%���f|�ż�m{Ϳ\`&�^����W��~�ǵgH�|���qu�n�Yv�Qk
8n���o��Ki�������_��<���q��E�Dg�[|���t���oԬ	j%�.&:�[�^g�%�J���)��S�UH�%��(����#�	d��C'��aT,�&�C��Q�A]����=fP�a}�|4�_txP���}{tzw�ثKL�.q�;�����:�QC�5���VN��)�qǀ�PA��u ��A�d��ŵ�xv�����K���#o��"h/��Z��甲 ��zF��&-�|�h�n����ҿy��P6�i���ת�`S��f�Z7m��6�yd�&[�ĵ��ԦQtp���L-Z�5�mըQ�V�͂�6oٮ}� ����"a6U�G��E��R��L��iB2�;���"����i��$8���@�v�C��c�5����.B(%?�:���y7�e�L=~WY�y2p���Ŏ]���U��r���n*Q(�~��V�������L���4S&���P�)t�`���!Kkck�#�u4v��$T(@���+z|��n��ka}�9��|@���O���pȜS���{s��T.dXm�\�����#�:٨�v�{ڍ�5vgԘ՟-9t�6+_�$���2����/C�EQE���W�@TO��v���dz��|��o���Y�OK6�b�<�^z���s�Ʋ3��������R��!/9C��/]�@^y�t�%��՗)�.Q�)|lf����S`�	:��8��	
F颓�E�HO�,8Q8�hޜ�ٳg�IF�P��CE��(�(�G�y`fx��Y��8�=m�O�eN�{��L(�'�3iG���Ҿ�|s��러��њ�cW���40nչ��&���6\�g?ߔ��g�Ư����7���g�R�O���h危K��^�8b�z�c��1r�`ļ����'�ͅa=s�a$ Cf�<�ܠ�gL?�.��	�Hbq����N>�������|�����U��k���:{��O��eY�Id�sv�j���vqˉ|Q�[R澐e�����7U]G��X�T�{��7s+Vl�	"�j��O&/��3D�*8�?�e@p���﷕�o�V-[����j��A�;�t�ޭ���+i����J�i9Ũ0Dd��.T2D�'����Ј��؎�c���t��	h���A��-:����*:�u|�vݻD��ֱo�xD�8��v�����jܼ[H�m[���!*v�ʭwy���`�|���l!��6�7�P�G�^�EX��� �����,ߠ�M[�����5i���b�j����C�&A�����n�$,�>��>Q��UZ�l����׷e�f~͛7GGP;���Ew�����,����yTaUVDQ�(�E���#:D��i�!�NT�v�a�#�����o�D�gаџM��taD�/.�nR5�>�����>�F�1iŉtnݾd~���]���-�w��KN5jJ��Q�.�K����z+M�g(#���0l����z��R[&���t�چJ1����Jai��t�������տ��������kc���?I�W> �+y�*���g�a�~��t�O����2�w�>�Bn�����m�����5P:�P�:�fek�-T�����-68���{�:<旸��:������O6��xc�GB>��v�f�����õm>Z���U@��Um?]6aU�竽��bm��k�)|4�G�ڌ�P�& ���f�Џ�x�d�x�����lC���7E~���W��d�6ė;:|�s���1~�G�y`fx�W�"'nm����	�'l	�|{�ĝ1_�7��߀����՞�vEN���6���q"���͎�ɻ:�k�)zL;t��`�)����������{b��r�Ϗǀ�?�8���Ѐ��zdдc���Ǉ�81l��a3O7�,0|V�G�N5�ʘy�c�]�t��E;ohn��=��=��P��n��y��Wl>�u���՚�7<�{���fl<�����S(�u�L^z�J��Pw��_��ˤk�=�.��Gᕻ��_����d}����~X5j��N}B�G�	i�.<8��ې��!A�Bۄ��i�&�? \ؠ"��ɧ旰
ȼB�,X�Sx`A]���ع�'O���+�S|ǎX���Q!�C���@7����޵kd��{����+�_�x�0�^]��zE�%ķ[;�����e���yߩ���id�]�D�X^������$DH�u��ع�P�e�
h�\2�K��{���M���4iҴq��?h���A��>M}[~��(8�I���pB���7��	���!��l����@Q�%To1]��{w�6xb�aSr9�b�!�!)`H
i�b����,�I1���4-**�u�ж���;�u��ۡ[GDL�Pp!�ݠ�����}?���݆ �Q�k�_�;g���G3VH�=�R�n�䵷�ed݋�A��^p�)�@��Q�.��0�̕L���T�:�܀�� ��E@��S@�|�E������Ia+�HZ��м�Gfo=6c���3�pg���ޘ�z_n&�R���'2��C�����i�K�bg��{�_���xX�R�@`rK�n����]m�+l��se4XP��ˀ�D�#0X�%۪'�Q�n.��}�D� G�0[� Kp���G�b>���
ksUaE��*_ZY �(yʚ|U-��U���,aU��&KP˩�.[t/Or/_��H��X�����T��T��9@�<(�g4�s��9��e~ɴ��[�
aq{0��	�26 f�������^Rt��r���6ԸW�Bpln���������[�� �|��gCp�h����sӴn�����0�/��?9�W|�+���
�$����\fz&5>�b�#���@�@�y��@�y.־��^�n��-4���c-_i�(L߭���dz��L�x~5O����O�^�mpk﹯�i�}�n�7�3Y��r���^/�Ū�6��r�D���xr2�;��e݆�:|�L�mݗ4e��)�7~�Ռ��=�b;Eth�!�]ǘ����ȶ�D�G��[��ҹ[�>/'&gf��K�����!.dJ�X2�@C�(�ֽG>�zʀcz���)&�ca�@$��@��Q�zDu��G��@�ޱ�z����	,��0�u�N�-����ҾMlDDhx���<[G�ۙ�2!�g��̈́��m����+��-��RN]Ni�٧�_�&�|��5��m�o�Z5mآip�oHP�vmڶ�G�j�2"�YT@��&Q~��h���f��jC�VmZ���:���m���l���,�&���!]RL����H�t>����G�ۅ��׻�^�c{�E����>4�Cxl|\�����<{ܗ �Ia]�ￔ�͢ݟLߒB6�QmE�����]���6|���a?��vE��!��8�R����&������`����J3O�w��&��.2��m��������[`ts�n����׊LUbc9�P`����
����n��Mq������j�d�j�2tz�����_m��ʲ��"D�E�]>�)��2�LlQ�6��|��?�*�����]���������W�+̠���r(U��J��^ĖjM^�jx�:lX#PU���}��T�6?�[�O����'����Ǧ�G�=��Vk��X�U�j��-j�{�<h���@cAh��X�a�j�Հ�T�6T*�A&G[��>�h��W�*���r���.v1�.��%����Rb���__Aj�/�?�����E�{Bu�@	_�����_S��V�[bi�]��c�����>HQ�b�]�s ��+k@�֖��
U�\Y&Vb�W+���f��L��p�BR����J��IQ��5�,���!Y���}	"d�_,݋Ba���.U�5wiZ����k&��|ۆ�O��r`��?��[٭��N]����t��Э�Ft�٩cT�؎]���1&�CT��}z:d��Իť��D�IldA��|��}���c'|9j�G������1�C`P�`Ds����@��z��ҳo�}������߫30�W���V@x��ց�ǅ���v�j�M҄
�F���JC��x-�̼[H�%���\ ��fz}��I��a-ۢ��4nҬU���M�����Z�iԶ]H8�uXxpXx`hD`����Ȁ����B[6n�4�i��&MZ�����;���Vm�e火��ݑ�Ч�r�|���&*��HT	�&*��(T�̙�;u�ݷO���]�c�a�®��g	Dw��~����t҂^þm�i�\�k%�3Yt[6��V��J���mQ����T�TV��݇����O�}�D�V��r:��(�-7ޣ� n�z����&���U�A�"�\(VY�:��QS���Ҹ��:��!jX�����������0S�Fؕ��:��Z`v	�6��
�_o�h�B�Y���Uv���~�L�RM9�b�ss�:���X��D�*d_��o4 ��3��	� 6Xe��;��b�w�ʻ�e*��5��N�H���u�I�����C�׈E�+ʟ�V��
�J�Q��:��(5[V����N��a��lZ�E����EC�.sCdN��n�8M2�^^�S�UNYu��ZY���)��s��Z�Թ$r�����,���w�n�NJ�u����)��|�X����2��h�1�q3���Z�e�Y⍿9���@tJ�����*'�Cؿ�U�4H4�^��j�T�y'��R��U��c��}X���,=֖G� ����l��ZZq��k��sI���e��K�t�ڳ_��{v�׫��>����گG�=����9>�cLTT�X��v�ڥ瀁#��1���|���%��P�D�X���?~������?�]�o؈��z�.*
�M������=z��ߵW��=�E�;��@�8t��������Jϰ�Q!��6amۆ�K���عo��c�(R*�Jb�"�Wi(���"�!q0�1��rY@���������#|Z���i��4��_4ФUL���M�b���i����)(�s� �x �?.�elK�ئ�c?lDĎ6����е�&�hV˜�����4Y>MR@����D��8�|:!,�}h[t��L:����!"4�CXdtxTl�����������{��:o��	�/�?vzT�W�������"ѽBѣ\��,V]6�^��9����d�#�q���i������J��A��2K�;"D.TX�
�CL���i46��2�{���
 �`)\�}�jR�Ct��.6���آ���$܂B�A�A"�7�^ol�1��P[%�ֈ�`���-���T��?C��h��|��o��ZxF� 5�G�b�Yj0+���Zԋ�or�P*-*�A�P��R������GYu�e�� 6͝ph���/��ũ_��;��oO�������,8sp��/�����K.X�����E��Xp�y�Cs0fzI�ÃwJ���g�M;�{���3Nl�~b�ԟW�ݱ~��k'DJ���T*�Y�2ج��ܢ���R�X $�B,V��b>�ZRZ����S$��\�J��Z��j��r�w�E�E���͛�����Ea`��-�Ft��C����pO[����p���T�+ҕ�l�Q�����A�'�_޴������0uv��c�""c"#⢢b"ã#�G��Dg�۴	i�n �1:�K��.��t2�Of�J�������Aa�,���˵��fβC	ɛ?���5#>�2�o�z"{���1b�G��X�e��3��4{Ѧ�?-,۶h���g�4ꛎ=F�uԾ���]�G�lӭ��5[�w�	l�
�Z
���"$�/�P����(�;��vV)/�$�(�-�%eso�������M�>[����!C�����?��VQ_�ENh�Y��O���DL���u�Ć�����?�o?>8���>?����{�?9g����-΢s�<�.��)��
i
t��&)��~%���:�����ݺ�v�ԥg�ν�)v��w�!���i��NÇu5f�ߎ��x��K��?���"��D��D��k�}��_��+\S￪9�l\U�qUt4�w,�q"�2b��0\�=���!E��XBjcI-^�u���"<"����J���4!�Bt��P�� B��u_���D�w�M6��"���������Y�Z|�Y�#� Xq�"^V���m5_W!��g�n�y��f�/%�h�-P»`odx�ZЂ�_�*B�UE��`��r�U-jp�E����|�Z �p>����	�~�X�Yآ����h|�u��7~�nR�I��}����k'b����������~��{��Sw���G��?-�mӚ{�R��鈍3�o��qf���N���S��?�m��~���{vN+F�M�3s��b53+������B_��rD<.(t�y�����r#M&Vj�����a���;V	����c8|��!<jN��f�e:��p�ܕ��ز��i���0�¸�.�񝻢[2u�B���ֹK�.���iץϝ�b&O"$3$$�����$	%"sG7g��v�ǵ�2�i��"��8�e�8�N�u�غ�7q�U�4�ˤ�.��:N���u�ς�>��mx�BzNn�srp���}'��7�̀o���ض�����!q�:��x�G�'e��*����s��v.�"�	�r����|��9!B"o���&�ȣp`F��wI�;$1�Fi%���7vu5�˨������c�~?F�5l^�����ǌX�=tQԐ���G�ې��s;�=`v���qC�t��ר��G��>��cg�[u0�X�IQ���� �%�t��N�bҭ�Wnl���i���i�g��2c�SG?m��?�v��I�M�1hҬ!��������7+n��;T�wK�j�����b��o���y��羚w擩�?���W�OLZxx҂�'-��ۅ?O�qu>��QT1e��|-BoQ��"TrQc:"�P�^xt�G��+�-����P�0��!�uX�"b��\�ӳ�ҡ�@F�D�������
��� :���l|P� ��*T%x>	�_|B��z����̀:/��x���A~�%�ej�Lc�)SgO����ɑ�	6|D:����=v~�z���GfF�����v�~js��ߵ�7��p���ly|F�S����:;? �pfaK��"_��b�q��KG��X�|ߢ{��:��������\�M�Z����eq���� �T�P,Q*�r�\)��2�\�S*j�J*�
E B>G@**=v��R���Jar����2��x��P��[���D<�aң;�zg��M B��x����{n�}`��=�Vo]�~�ڍ;�o�y��0�qĆ]6�ټ�7�mׯG=w�RrV>����b��� ��$���o.�I���bE�m���ө���{��r��K��.2~=���,��e����_���e�~�S���?���w���M��4�t��ۂ��y'2�D�Rǯ���Q�x����ˣ(i\��`�m�9<�D�!��Ӱ����ʧ�6�%̌b��nz�0�X|�X��/8�F>t�`�ɔ�./�sn�Γ�~>�p���./=tm���Go�:���=������ol8~}����O%�z>�ȕ;�������tQC���!2�8��S�ϒ��9,��o��=�'�k�>a}|�����>�'b�O��#E�n5��v�t����L[>ӒϰL'P�r�����

��*(�
��"�P�IA��$PrV�yA�b4�_˯(��:���Ӣ�잃=(�*�2��RV�H`�e��q*�����%PU��M$���p��U
�cM�s�퉾��RW�%V��(S�����W�Im�5��i��Z�(��Z������)�,���:w.���?�����$�gb�c����@j{���
�s��������\e���O{�������(��LOщ6�ޓX ���NǗrl.��������O|6N�����Β����������0���و�_4���W��l�P���\��6i^��D�\��8�֒���b���Q@�
D�J��U���������&��Vw��2�ڲ�k�bN-l�w~P�����l�U���H�\�H�3 Z�V�R��ȅJ�L.K�"�D*J�1�P�P�e����R�7��N����*S���N��3��y˂ >]�ĞE�!�0������.X-a��*�w����:o��ӗL�~��?.��Ӓ�Ӗ~?s��VS筝�pÜ�[�ھ���+�y�%��RA�Ct8@"��I��/��Il]1K�M�'g���Q����ݢ%\-.ޠ �o��sI���K�\->}���Uĩkň��37��R��o�����.��.�Q/����lf	W_@Ӕ2Md�����xv����(�b��}��+B�D�Hꏝ���0��O/��ҊiE��~b6��-��빻ϥn:ze��sK��\���$�>zi���5'��:�X{���S��O&n:uy��k��_ߗx�؍;�3�S��4A>K�1�UG؅G�1d�LyK��Rg��\�Y�k��m'�o<2}��Y[��ڞ0c�ř;g�2��kw_[���-g6�~�襂|����Á_  ?E2[O��i<Ch��t4��*CD�6�:�D�V�Y2�^d�&H�<���@�F�� 0U�kB-3ó\�\��^�.��E�u�U��AS�8�J����u��.�
(�S,���bC-�q�27O����'0<Q��n��~6Kz�QG�"uUn��+�p���Jiy(5ݓ������_{�����2O�e/���u�[W��_pYZ�1�3<�9�4�}�����V��"��R��.����	�u�l3M`*+��2�Tۚ��-�i*"��r�ݥ�5y��/��&�8M�8Mw}��Z�1��OA	��@�	3C�Nk}zJ����O����/[n�s����#��v�1/6y~�ͅ����o-�K]��,HY:����C�J��U�#�VF"q.�JX������?��q���X� 3�2�Z�7�%B�T&#b�ŀ�'Tʔ&�BB"��n��K�����"|�m�%�%xE����B/�-�xE(P������.��I>~1��ԃgS��}�|�	w�\�<z9�Db��9�.g�Ƞ2�%LEY�O�S�ET��ס�C�$������������K�C��F��BJ�Qt9�0�Fp�Fޅ伄���7��n^L.��R�x�t5���m
����[d��lv>UU�0�f!�e�����U�Dr�B���KB�DވD�šqĹ$�-Aw��
3J�%|\�)y�k����.f�>sk��k�_�t���É[�\5n<ve�����W���J�}!����G��O�*��EK-�gPe��|�<(�0RX0���b�ҩҳwȻϤl?q}��k;N��:s{����g��9�����	��."��I?q�$�D��҂As�G�T�|u�@K��]�DG�)2Vz�Ű��@4"7�)�LhV�b�Y 5�:�R�V�.ě����JFt���0��(0��֊���֖A5v5�{!�LVY�Z]�P�V��t�E!Ǆ��K��B��#��r����GB�K��!���A.d	L�Vk�69C��r>/�Ҋ$��|����czT�v���(��E��:�˭�r�eE�ªB�}��xT(���t��d�ޥ[�)O�f�D�G WYe"ީ)�BC�6��fY]ԯ��r�ө�3i��	��'wHY1t�_��Lj{jjL₮��ğ�{fN̩9���"9�C��1>'��M������K:&.��
�݊� x.yU��U����J4LZ���
D�Y3����B��Vc�UB2�.����wZ�^��!�J�E*�r�!V�������PN���t�@9;���5C=b�ًHi�o�/A�¨_8:F�~�^8�w@D��u�z�`�dʭt��.Ix$!���;'�枼Zp�r���yǯ��N�(>�L:���܋)��"aY�Q���ߞ����A�V�5�юi>K�E���ޡ��.���n]N#�O.��R\�U����ih�3�$X)I�v�ee"�0�v�6��mFj����2-d���4 J��Z(�8ʫ>}�������W�|�����x��b&�0�,�*�	��W2��oQN�(:|5o���]'S����P���W��[����_�|"	�r��3i{/eL*<v�|�.�J.7�D�N�g�U`;�C��� C�C�e1�]�<��w�z���R\J��Bگ�n�v>�>���;/�=|9�w.�����$)�#��P)[�͑�<D_�/T�5@�D_*1���R]b��ѡ�ML	Txf��@e��B�Q��H82)J
�\�T�Y=r����
�!ԅPn��k5�ӱ�1Pɨ��I2�����h�Tm5CW.dh�G}��ۈ�Kw\U��go��q���c�F�h���>�/_�7Mhss4y��,P[���s�����OK��_N���L��N_�۾���|AY������+a�>o98�פ_Γ�y�m'n��>n贸!��>�#�}�ֻy&��[���4����Y�Q��5�oi%���:p�)����`>�
A�Ns:�z+���P��zмM�Lj��c�SSc&�1)�.ח�=;7��<�q���q���p���~���̈�c.,�xqy���Q�VF%�ꐸ:�ʚ�kk#0�57�F�\��:��
a"p}uXҪ���pa�5v�J)( �hM��
"��P���P�d2)R�T$��9<�����G����*�] ����*�C���z<E* T꽼�Ѓxk"��!QqdJ3�Q�2y������ǅ��\hϦH��;y%�tR���Ŝ×r�])>~�q��B*�z$>�["�.g�9QE��U�	�X�1�ME,#����T���|~�څ[��SJ.ݦ\�KOH%]LC����^��JM�\N)@�WS�Wo�p@��ә@j6��
"4�2MT�P��3_�+u��<}����?�"$�:R�G"�Ê�(�����@�wHB(Ԓ�W�����3h'�J���?t-��P��<�����q�m`��7w�M�}.ؕp���w��w(���]����bQJ�,�*�KW���y�L���$�.ɡ��hR �*K-���Y��̭�O��;���\���i��9����x;�V�".����T��P�œe�$�|i�@V R�"]�XO����ï��0l%�@���ٗ,��*��'���T�Q���L�,���ʍ<��+CH4+q@�|��L�
��\h{>dҊ^���4f���f�O3V�O�|q���?V��,�'/��?co"��M΁d�������wYA��ck�n��^���ic��ت^	�#~�f�n���/�s�t���K��J��_�!���HaYW��2��kdхB��[ԓi�CW��vg��2uݱl����Cw��������dF�W�Ou�v����z�Pׂ�=��_��@"1��o�LZnW/��߾�����B��	�u��������1 ��l�w�b�$�}?�����1Ȃ�#.�iwy]����Wׇ^�\�zcC���mo�k{sm��:HZ���ݵ���k�SW�痶<�0$���j�@��Y�V[�Co53��P��(�*�R!U�%r�\(���P�ˀ����R�D(�5p���kH����c�
�5l��x�6�ޛ�`�8`[�E���T�P��fC�<J�QgX{)<��V��s���N]/�Nԑ���Rt�zѥ��w�iy��af	?������Z�a�eHL5:%�2�X��a
iƴ<IV�21��z�}'o�Podr��eAmJK��`$9�ܸ��U�����R���T���l���vr:#-�SLW���\��c	L���Uky�}(�>��/ �F���"�W���B&OQ�g����(Y�B��(\-$�2O�)=~���ͼ�׳~OL��B��n�3�/"�t;x�΁+�\�:x=珤��)'�I����dq*Yz�*�C�e�$Y4q&�|vq=C*�`�nf6-�[(��N=	5�IBU  4#IDAT��n:{��T�#gS��O�9v�֥���ELX���(���戁\�$�'-(�"�&�"4��W��&�P�1Ez)#�̤�'��3�˼��¹_R��d.��ק� N �"^&�qБR%�G�v��h\].q���e��消���]���j�=�!��'(n���t��=o�m�l��W�n|�\�e��%;K2�e\C��O{L\�t슑�.H�ϴ��|��m�N����b������z����yw��)f�܅��w���y�n�_��eqJ�c�����%՚Z���7B���䠛���vw�f�W�W�� 2�5�u�_D��VxD�w
e�J�v�7}~�uhz �qG�^^ni�����ő��g�D��g����,�,�,��+cP��5H��և\�������M��l	��%$isH҆����!@��6�� ����m�K^�&yM�����txj�K�ՋK�$���i���-F�Qu�Z�Uh52�\�D(�������@"�P�y%T�(��Q���a0��7ߛz��Wh��S`J�� ՙdz3��÷�����k�J�L��y \��Ɨ�R���*��� %�䟻�s�Z.�j�٫�g�c��R�p� 1�t�.==��Y��,f�8�dv�W�3��BKIbjIL=Ti�L�a.���iƬE6Iy�rޢu���p:1�V� 5�JR�rR3�0LIg߂�]L�%g����L F�<@�P�RX**G�!�m[��-���sp !B"oD!��_�� Ub5�=���C��)��&sSH�j-!��̝���r��fLJ����C��q_�p�Z��+��&�~�xR����7�N�f���.��r�z	+�¿E�ӄ@]�I��E X0��v*�husS��!	��v'�u�Fh�S���#8�Τ�8_υ��bx4�*ȡ	���J�9����/J�J�j_/���
���щ=���85�Ό����$�<yxܩ�[�Z��Z^��
�;�>�X/Bvk=�D肊p�7+{|�*fĢ)���n���k�~<�bH��S��sm�y;��C��+r^�Y��3����ĭ
��]�3�J-L���~�i��K<S-_a�(���Ū'���gm=;r֥|���Uy�K�ê�ܺJ��(MWe���P�t�)v��I�o�dUnu�{����pXfuS�5R�c�#7��@�tӤ��jtH]�f<5j=Wpst�P"�S SV����gfԾ�8G��z~]��QǗFz9��î�[n���o[����btP���؋+c/��xim̥�Qַ��>����K�C.mmsy[ȕm��nm��	q}s peS ���ե�-/ni~ys0"��W����u�eo�F���-f�٨1�UH�:�J-Q(�r�H���|��#��h9$�Tk��7E����)=���Z�.��*~�E!_��r��{1*կgÞ�9�n~�R#Sh���y �|*X-R-K�*��2�)�WS�.^�H���p5;�J���9��\I.L�K��K�*dd��}�J���b���d���T��j2CKa�,#��+�h
(*�c	C�U$��ÿu�u7WP@Rd�ngrӳx L���g�`$-�w+��a�<h<��e���H(��W��J�D��Y�V�ç/��x�H���[Q*�8�ȅ2=��ɓ���&/�ʹ[�L/��*�&�_��?w;�dj��i�o��r2	q�Fp6�m�ݸ���~>�NBjFBZ��Y3r�n�����`�T�A�fP�YTv��G��@�9R�d�W��-��s�[�g/����
��x��4�3�ny&^J�v;DF�@�cs�a![Rđ���r�@����!��$Z�L��ƥ��"���~�3���!gO|4wf��-W��+��ߊPi��gtp�,\���0jʆV���5���� B���'��_��揙[3�v���YA�W���<�~��w�vď�IJ���:�2t�jw��>�|D�kD6�����0dF�᳿Xp@R�N�<h�w砉��O��ْ=a�f�~CB1��*ϒ�Ⱥc:�eԲ<IY��NV�2a���Tn���+�Z\]9CR�W=���4����"�����EX%1UH�z�A;gbߟg��2' '�ظ}BϬ�?�2���H/��vX����>;�����VG��9>/����+cί�=��㹵�g�u8�>��ư�ڝ��6a[����^����FT^���9��f a����~g���������Y�si�C3v�� +���"���e�]h�Z��Z�Am��U�\��-���L�T�@�X��zb.��El<���� _��Jd ]�@�� ��0�- |Ά���!��CȤ9�*R�pG*�����ЅPM
dj�DA�
�;��/M��O��y=%�zJε�\��7r��)y��%�y��B&�/��(��
��b:���'1��2KLfI��l5�h#1�4�+���_,��EKM/��c�r�!�W�`$;��er���
89��<�'�D �٬BV.���8"�@��k,[Y�Ǐ��|��@���;�Rp�:Ć����2&W@asKl�Y�d��$RzAaJn�����,�fV6���}++�vv.p7;��) �d���;9����;��w��3�K�(�l
=�� �hl ��@��
F	���Kti"Q�휒[�EiE�w
���|�H�I��q%%�VNIf1=��Ԁсl*�a.K�����2P nA�.Tza�T4�
t0�: t�.�X8<e~^����ܷ�0?E(ԉ�<��3��k�G�z �� �:��z��J3G�dj�LZ����s�/�,��[w��}Ԕc�Zw�q+f�H�9��,�;z׎���R�o��E��[tY�Út��O���e���u��m��l�S��|�n��~�N,��@����A�7�j�mzl7�Z��O�s��\�_��7���}��j�=�̈���u����0<`h��o�>x	W�B�����������ce�k���!�LU�,] ��S�f�r愾[fE��j�ęm݀S[:�wxm􁕑����'� K>�Y<�g�����ǜ�ǖE�Z{Xs|-u|m�uQ'7t8�)�Ԗg6G��qu]8pa}�s۞��8�)������o
<����u��׷۱���}�z�Ơ(�����;��.�Q^fu9,N��n��\����:�D��J�'�x�[��Hi�K4��d����E#��$H��J�41�`�_W�Ȭ�\2)��J ���#�E"�P�<�'����C�`|�G(��$R@,~�T"dR �+)ht�[�`���c0D�&3�B�/--(��(��e_�.���*��1�R'�#�!@À?��K<�d [�b� �'��%t�����Py0��%4�ԋ�!&T�^�k �K ����Yt����UXN�����f��ZB�c��Y�\�n�^RRB@�D�n��iXDJb_��y������W�bΙ�ϙg�Lmme��J}��A!���]3�tA/&���3%:�9�܋L��D��:=��R@�4,�d�L66L�W���	�.��'�,�.�N�jT0Y�ǝy5C̰��*G�0�?e�����H^�WP�J������ �X�iDog�N8�k$c��1*�-	�]Xk;�VM��[�[Ml�j�~�p���H���Ň���f\2�xR�$�o�:|[�s���!73NC}�E�M�e���h��Q'�[!���$��W���T���M��wӵ�Y��Kc�v�t$$6�����;�Q�Q"1�3���R�5Ƣw��ۘ�;ٯ�b�g?�
(y�;b�L�Z/S֏wyB�Ǝ�DǛ�=C�Y�o��� |\��k��
�JF]�Y�߄�K���lď�8�n�����+Wb>�3����O�-Fo/g*G��XAME�o���㥬H̯� ���f��VZ�(n<F�T�L�|�py(�#���w:xtnfF��Q
DnK��4�)tVWi[$5$(t<���{K�p?�f�p��b�/Hy��uQ^�����*X�	6<i����Y�C�a(:�s�O��j�z//�Ԭx^cQ��6���
8��B��?��B�Ρ T���5�̋p��D.5�<o%���`���VāI�ՊQazE�(�N g�<�:�cO���gE�0�A�J9���1��~~�衽N�*Ш��7�k�i�A�[�Q���LY�H_�J3�K�����n 0��b{� �0Kn��L�����p>��wG����(Mf�BT��-�p�;��o�bf�*΢�� �~��W�>02����;�/�O�h��e�-I�n6�Y_xŒ�"�\S�qng�g�`Hs��V�Ʃq_�+peh�ڡ���Ui$V*��`6n2K��V��%�9x�b��Z�Y�vr��-\q-����8?�g���>��x�ᳶSH��."(�Ѿ�Q5���צs�6J�A#�����1���1S�YYt�5G��Xn�O��j��+(���́3Y֋x=���R�򵱅%�[��!�ޟ����i���y8�O������Ƿ��~�v?�6t�s�}x۱ g�9�
��h���/�X,�4�~�!�<7�}�7�J9jWsEdA7�����R}����^����6h:�+\�F�ʄLL:����A��g#w��Hm��7!*�ǀ��@d�I�AC����l����2�^���sr����
'm#��&%-��ڌ���-V��e���֎y��|܄ϣ���ܬh_��Z���h�:M*;��u%#��trWZy�#��z�t��L� -hd� d��jg�T�<;ᛙÌ��W�H>�[��5�Y7�%�=������b1�+�7���)�Ӭ���o���R��3_Y@(o�Ɯ�Ǫy����U� j��z�L`�y!qoa:�r΂�����7(���J�e���j�Ю�������+�:xl3�n+}��]�V)*�X"������$W3 TX�KÌ�R�J=봊W��!�\�H��I���!i��?�����-�g���+�&Sl7L��C`7��QIA�gǛ:��=�廗�.�<%b���r�6a����srpn܏� ��).>e��d��=���^�g��0ѫ#�P)���%�����X����d]�^�P,�bS�Y�bl1�Sa4ґr��|�.3��n�\97�MX�d���u��+��[b����w�d��C�1tM��Q�|���%m'}f-�xT�*J-���3w��8p�i�<�4���o�@'��<�p�xVe�=E���b��/-s�W�5�\�y�2U�a���ZiY�sr=ࣝO��}�����/$�7���_K�O,�i�&߶��C������gS#-�X�硾�������D�S^�dA�#TF���[f����HC/��OI�_�q�@�Qg�c��S:���*dJh������qrӷ��f�,�/�[��d*o�N�?$2n�y��"��#�SbҀ�{�\u��X��f%1m��*m��ᵆ������P�qB��^kM
�M߬��.��{�%�U>z��h��y,SS��	�٧���B/S��zo�}t{v��J'���|x�}X����C��}mn�d�ӏ���ɞ��]CV��}f�6�OP�}C㽺=�~x���RRB�)��)ܔ�u�<�[TQ�f,��,�@�X2f��Y������V	�^̾����_�"N-	�#,��"
ТM�¾\���(D2�_=�Q�-� uv����,��ρ���Y���81~f�1A_PҾ7x�yS	p�N;�TDY��~l?��sO�h�dg&?T��\��m�΋�N"�r��x��N0r[|�\�<�4��i���ħw�x��>��E�a�$)���J{JF�T`�-���R���nb̛ ��aV�$D�s%�m�l�r�}�\�9dF��4,�.�b7�� �O !�p{!�-���.�NE �ذ$(�|,C�$���1�2���������0�h��@�Y�؍e���Ab�j5ц�Z0���ªŴ2�K��O�ۏ/�SN��jV��^��PTB^Ħp5����o�#M�2k�??)�+��������?�����6���,��ty��"%���of�W��wTg+�u�Ԥ��_B��4[-���?^U$�	Uqҽ�T��3�=���{���n}���Kc�X�aZ�yb��@��29tv�N�P��u�Ů�����i��~���TZ�87u��ʛS�T�F}�b_َD��Π��ɎɎ�*ۂ �4�e��>£,"�34���8���3�1�@�tU;`�!;�	\���M���~"�2��b%���9�g뗈���F\�U��@�1�z|rH�%��#[��F^�!гɭ��4���q�R7������ ������w��%^�w?��*�o��4H� ���D��4�o��0�������L��q��v���E��i��N�5�N�T��.��|ۮ��q?�s���7�M�fMB��5�5�U��Pà������������, ��r� ?q5Ϭr�`���R�g��=|���U°cc�OȊ�(��U��`�v^��sR��¸�ˠ�_h�t�0��@��~�/0r��H+��ٳZ[�n�X,GTM�����-��tgոx�uŢ������
�Z�����k�PM��ք����yp`�wLA
���(��h����q��U\��c�L ooh펺(o\x�wce�����j�2�?:�_A�&N؂�X��Q���E���+���(��F
i�>Է�����-�;��U�G�x���fmż�"^Y������䛎2���r��˱B��-̱���m0r	��U Oe_c���o:T�6�#��M�����:d�G�x�cT�?�S�㐠� Z`���C ���?u�6�4yχ��ƶT��l��`t�Y	��B�ӡ9�`��v�۷B޾܁���!D�܄���kH%�����@�̰Ϧ���\Q��z��vXHPY��s��ܖ	3��2�ֆ��`�I�Ʉ5�h ���K~bs�]<��	M"*j��ݯ������?�q��	�����k��-&����;���ȷ h�$4>qTF|����n�����C̰X�P������w�̩�ڪ�:&u�]w���^ؤu��,�B�b�j�V̘���#a�m��w�tY������l ��|�h�Ѿ��%�d��� �<��M�NEry`���I�VX�"@��)�"��ǻ�[�5Q�yY� ꨌbgǕ&�S�*����U���cH�Ԡ4� k���L�+��������|R�g��0����mO��*�����F��Xݒ|S��1�/�&[�d�2xCibaR�
l&�����X��dv��[я�(� �2Z����a��wlU�@��㸙�감�ߗ$g�K6�����t*/�ie:>+���@�>-���e�� ۮ�墩Ŷ3/}?B�#3�\�H�T��?hJM����i6�Д9��j-k��c߉3��3<�?���ʞ��(
4M-Ǟ	�=��bF�fN�Ty��%cI�0��1%�Ž���e���W���m��ki�����N��I_шKKP�
��8��`��_��Oqi�xnQ�M��a�AVTj�I�O�s� �f��"x���j�dXV��aG���,��Q�n����繴�dwx5���zCeT��LB�LS�1�;�E���J�҈�2���ɝ'p	Ĕ�5� �4J�����|������b�6�9�#7炌z����x���y�k��*�>{��c.W�C�]�ͧ�a�}A�����P��Lyq����A�U�l�Vѯ)%�H�P�����	u�dȁ3�ʜ?z'B,�9�t�W��^��R����Y�ڛ������L�ʀ3�����y�/��0�!�9�g`�W�A� ��v[|�d>1���G��#9���w73v��<m����y���څ@3�(���e��MEi%ޟ(�p�A�>�8�@�>�ѱ�E�N����3噃�!�Q�z�D�`�py��tS?�p�̸�t��Hs��k�B�mP#���BF���k� ������]�<�HG�������W۰���(�4�v�|�]��9?p��cu���D�|A�X�����<�Ȅ �n"t��Ɓ�mc���͒DYɑO���EK�7��EqՏ���ZQ����v��w�[�k�CI�n�䍑��Ӗ�#�*�?ݼΟ?~҅1@�e����Y�U��ߞԦ
������P��3�-n��K�)g���*o��<J�4b($�Dl����,=VC�G٨�2�3��g_��4�k�#o�D�+#X��M���B�Y��`�7��Uڊ����M|_(���=E�ڇp��;�1����~rn 6693�j-�o���Մ��~��\Q$!�t�z�15���Me������3��䫑I��lx���9�{��8���=V�JS��R�I�<D����5@QV��HQ�=+�6�`�����g�1=�lOe˯�R�Iu���_��qs}ĎH)�����!��%թ_��h���U���#�J�LQ�a�DP��7 Ɓ��}�B��,�'�߄��/�)P�)˲f�t�qE-�W��!���H,�oƌ��e=�׊�͊.@>�jeR楇��zbrd�"vKu�R��h��㬋��A�,ǲ��/�����d�;/��F�1��F�ƚ�6�6��E�ޑ<�\dmT3].�5;���o�
��]� ���/b�Ip&b~��	eV��]�-�:S���x���H-_[�I���4J8wZ\2Z^\�#��W/�7��h����W��;d��4 yY9G��o����Cn
�[��T vD.�0?��?pr����6M4��"�u�
��bo'5�@�zh��>���*4JY>a�񕿒�V���H��,�#����HƦj�!�ؗ����Q��rII�d*0��Im�=����6@�.�
pq9!�5.:l�yT��1҅�8��7���E��
.ҶjF`��U�l�X����X�K�N;��V��:x8�gQ���_������K�1n�L���#��ʍ{Q��5)�n����8qY���/ׄx�0q�d�p�x�u_��s+F`�iZUWbѲa`n��T���UI3���1��oA������X�1��F�\����3t���OT<�T-�8����@`�H�~��g�w�\���-UG�z[�4�ޮ������ߟ�y���OP@^�<*�(� ��O��K�y|A���b�Ŷ����I�6���b�$�qjp$9��X1ܒ@���߭��ȗ��g
��kAH�]y$���%�Vd�?�GF���Yo�U�#eU����I�7}s"����"�y�k�3�l�Q���ޱ:�&8���i���
��x
������:�8W���+o*>�Rd����| ѾO�y<����`�H�������g&oR�|T�U�+V�+,�\H��'�+��P�˲J>��G1�H%;��hi>xVl�m"5�I3\B����y�vSʗ%�5v�e4�<*Z���<lY$Ձ;��ل���ѓE`��V<�5�x2\���+���$0�R�8
�Ď`���:�!�� ~��H����T��`yctqN�bI�Е!˛�"���a�hz\-�R
�׸ޕ��W�#:4���6�b2P�C�႙�2U�A��!�
�O�T����Zao�zy��˺�2r���M��*1�K�c��m��l'I�ʯ=V���I�n:�ο6Ǣ��7~�xM�ʶk`W[�]�w36������7LQ�(�l�\�=	���Q�l�J���QNџ7N;��}?��N0����L��t���m�[�F-
VA> �s5P1&c���A�4Xf��\C�<��pɑ�Œ��5�ҼR�h�j�3�W���c��C��@�CZ��B�uQ�#�OOUY:��_h�d�T�C,�`°�}�n��x��60I�i����&2�9/��\��_�Qq����h�s��)q��'�ڣ4��GA@EGm���1@s[�	�؉��2���A{OD�l��B��m*�cӬP��*I[�l��1Ė��֗;[��=\��b�j�J���+��\�'Q����>e�bzoe���/��-RwĿ��Ü�;r�d0�, �LJ�M�򕯫�����oH�����u�I�Bm���9����Tg���������R���\E��ā��k�J�&^ ګ�V���҄]9�ִ�sS}9/�Ne��8�6�ǟ��V��Wu���0�A|n��t��I8fr����8(��}�ײ�OX�%�<��5t� ��M:R��oIxb����(Y.��at0�~�A>���[i��Hr�k���0	�E�c����+�F6�\Gr��Շ��Ϙޱ�￟V����H�~�����HUg!�Ƌ���e���qy}�B���K��Q�Q�i���_��/�k����������|���r�ԙ��}O7r3o���}e���88����Թ�v�����R��
��=��f�Z���Z�_Up�-�c��=%��֡��ޭ|r>-��83n��׀�fe�ڍh�[�[�s�+�?q[i����l����	���b�U�ċ��j�U`{Y�Mc&���4?����e�����7?Pٓ2��ͻy.�g�?Z{�e��No�[f!j.?Z(Wz4�r}O��.��P=!�=DA�.�v�h��7�oP_�ދ�m�:���pn���B�/�;��>�e?B���e�.n�I��.Н�����N~:���l�~�������d���M]�c�����j���9N��ѩ�gc?��5�z�If�)0�-��{�/��q�j�������n����w�{1��9�.�&Q&O��0�����X0e��
���B)Sҳ$.q�/N�]V$[�RM��2\{��(����l��v��J4�20+Z�A6���u�c�KF�X��r/c�-�u�o��	A�F��h�p�90u�F��"�N�9���%3e;������k��T�Ѵ1�s)������0���f%,.�..�g����F�|������Y��BW�K�?<2 ��°kWX�DϱMR�Z��>QO�U,������/�Ev�$y�ЭЂ��GMV��8U���L�b�{��9A��µ�	`�~W�@�%�-��5�0�<#簿\a�>�oh.�Ԓ���W�@� �a�&4�����T �b(�+�\"0�����Y�tQ����2L���M_����i[�B &�v�FeԐ���WzN?3���������e�y?Z��c�<K���q|l�2÷��š5�i��̸���`#a`=ڋ��>�U@�Ϳz����[0���;t�e"��w���VIV�ĥ��\i���-�_NUL�<��u?Q���>|�<#��Nq7y�xc�3px|?��'_!�%ѿI4�됼�3k����z�i�7"Y�����a:�u|;vIT}��uly>iI�Ybt�~0�Ҹ
�f���Vd ��/Q�fF>S5�#?�@��|��~�Ù���m�+�0���$����1 ��+��W�E������@v]"��Z�4���_P ���AC���>+5C��ɿ/<��A�%0��-��l6�\���7.��^�<ۂ+���V3��s?�K'���	��3mR���X4�5�{����H�Ç� �mV?�B�{/�',��� ��9-;��3 �_����fj�r�@�s�����J����C�i2>vv{ ���Z��w�Gt/@35}1�3�����˰η�hT��gȆ]��^�'~�|~�cAY��'��,1�A��G��:,��0��
�	��Y�����۳��y����DR]�P���<.�b��м�����r���M�@xK�sH�}�g¢���	í��ǀ<�{�ʕy�2m3Ib��>ju��̖�a�E�C�̙�eB=��c�6MQ�r��~�R���z#vS�#c�ռ�I�h����A���6��>��ޒ�c1��������yw��e����YC��I��>#��=a�w|b٨/�u����ӇD�j�7��`��{�V���/+��(W(#�i�����+s0�Gz��س��۴�|���jw��r�B��oN�.K��Z^����|:�ۂf�T��pt:���Z��߅k���y�޴nyҎ��B(���?�� (�T��V+�z�}a
H������l�t���	x��5���o��6�5q���H��5�{��O���
��G��7��r4;��5���CF����3�VKyծ����=�y}��W����0&��#�屩w��/.�[n�ה��,��SQ��UN�F2�1��I_92ܶh�թ�m�V��|X��WM��Jp+Y>��r����S�g��C�.(#{��+OXm�(��4��,�<��z��H�N1�ɳbS��
�N�l�9!vWn�_�wc'�@�Z��豫PG��#����JZ�5_Q7�]	�@��---����\�����)����a��aA�ƖOv���6�6r�i3<t ��u�"�f�T���WӦb3��Gᒱ�l�������>�F���L���#�'G���!R�?�������mC�L��hP�M��Gl�����_w��v��Q�5�4� �앪�J=� PK   �n�X�{��  B     jsons/user_defined.json�[ێ���� 	2������b	�[�C��e\r͋C��g�M95�%�;��uSȓ�AZ.gN�Tש:���i���f�������~�/VC?�f��v�^���"�e�o�������>|�\˽������۬��j�Y/qu�����/�z�@_���~W�=��}����CL�ڶN6P���%��,8���jX���D�h�ދ�f?�{5l���fw0�d�����h���y�[�c�!���P��\���kG�f��-�(���ֽmnj׮�ۺ飮�>����n�n�_�����u�c�t?��f�z���g/>�V��W��Ͳ���z	��LR��?���n�Q��FQr� �߯?��T�������c���v!��X�>6�c�HB���m������;�-�v�f�Vyl�b{���l+椼��bϛ��9�&��K�b�T0��Rp;�Ny+���W?���M�}���at�w�?����)�(�B�*ZcB)���`�z�/EO���(��)�՘A��;�.����Ltl���@�1CS��\�Q: ��O��9*�0RIW��r�3+���d0e�mqHҔ��R#Ex��I����൉*��!O��U�%Ud8(K:��g�~t8k�Q�s1���H�J������}���O)�Ⱦ���9HT�S�J�
V"ǃ�ޕ�J�+�G�uҊ�.��d�+j7ۤA+M	Ӑʫ��T��%'8S%�U$�S1z���71x�*���-S1���P�SH�
Ȗ�$Sn���'ۃ!�D����3�<�M�b��K��3���#�l������dJ,�Y�15A��Xn{�Ğ�CT3P�kl��J��S�0�q�<�Y#��u	�ґGG����
��NJ�KN�0��&��$�OҼPKtH����k1�Hb�d_�b��_�nBJA$1��/��)a9"�;��A;��k3%��FA� �W?�l�Qyɿ��1�����N9��MȘ��D����tS�F���|��LO>��uS֞��A�e��S�FBB�6A�*"+O������.c���Vn�Zq�`,�G�lϱ~��3�0�s3�S;e-W�vT9d4�}y�㦤��Li���<XP���,����Rf]�g2�=�b�T_�X�0���X�h��,g{�{D�L]x1�����Q&��U��O6��$O�
x�
�a�ү��rN��q����*X{���2�	�ce<A[R,�Ŝ!,���d�X�l���;<elB~���g��R6Ũ"����{G�8<�,
8:@+�0���]*��S֒1H�э�c!����2�OyK�1�|H����5.&E&��?I%fW�,:�.��������t9���ƀ��*c1�� ���O�k�	J��8�n�Pyn�S��\�7VQ���O�k��1ш�x���gJ_��I�%�t(���S���N&�_1�f�|�1L�Pق	��2�������=�'<
�/N�!�_4���Ȧ��?�kِ�/%��RzD� >��?�B��ucYE�/�-�O���z��-+Q�슕O�𗵴�H��ʯ\ί�᯳�38/���P�����I���I�Pj矐��[��IVHЈj[��b��g���������:#�09#����e��9�B9#%�*����l�r��Z!�Y�עU�.Xʏ�:% eŉT��+�?1�_)�6�������ֲ�@/߃�9�JQ'�(�h�`q~���ͯa�R�T���U&J��?e�{�'t�A{*�)�_��|�9�s�=�B)%T������2���)WO��F#��y���,��qc�S�~H�:�z�Hw��a,o�R��w�<�c��X=�{��p�*o.R��'�`����t��g��n]|q�Β�:`���єo��Β����Qi}Ao��:^TH?n��h�� �Ί�;|���]by�N:[|�4�UQ�l������{��W!]�6@:�^&ddv>V�C��1^���G�e�(����hS����%+��{��9;e�����Hd�|כ2ǧ���6����E<�5��@���!y���A����e�Pa ���\�ʛB{W��O�ST�0H��N�eHl�
>PЎ�v���� �b &-���e�6)s�
.Jr�Q��+��. ��u��6��a�[�:��Y��邃�9&�h�y�ոY�P��SE�L�xF�$�̉-�Ӥ̡��0C'���	Ɩ����:×�5���L�9X@�w�9Hh�l�e�V��߃(9���9\5����qc�9��y�9^u�B�xS9Y�O�;x�*9�������f�1��f��6���>�;1��+߯�����|��aPۡf�L�R��)�T�$E9ts���ߛh��GG�k����M���������wz��_7�
�їЙY��Ĝ�� eoQ�
^r�q�#xL��		*{"`�_s0����C/����N�5�ﻶvܷu�t}�"���up����^<�#�����_l}X/w��j;����U�]='Ɔ�u�a[sh絋=����ϝ�"�7�X�>��`����3u��n��	}SC�5C���f�ܥ��6��%B�R\����[�{4k����Oȅ�,s����dO����`4���W���v�~�,G4�F��Fx�����O�?����,��'������W��z���}��T<���}��o���D��_Y��.�^��wG�hji���=J���m��Sjڶ���Y���Iw��vȝu��P�mt����;��	���]��}� E+-?�>����U��5�\r,p��~?���v�d��� 9���'�8^��!�`�	z�#SFaG��'L9]�\S�pWe�]U(d�c&]Y���(�^hڥԎ���v�{��������1�!¯oV��Y������Y-v������7��(Gd��b������~ޏ�#@�؀�j?o:���l�7ÿ����.�_�0m?���w��t����I�nP�an|k#w&�@��P�����n�y�'�h�0�(MMh�6����a��@v���b�ͳ󄷍�F�m�xM�u�-�]2�&?���n/,�厚�-E*~�+���eO��B�;�<˔߶�ka���V�K�Q5O�~���,9�O��G��������'�x���Y���?�*�s�;#gc����i�7�%
޽qg�'|X��'Fϴ2㟴����w#�>�?I�g��h��Z�������f~�E��'��� Wq�5ֽ�m�����A��7�q��2� gcqFx��� PK
   �n�X���e"  ��                  cirkitFile.jsonPK
   �m�X�l����	 ��	 /             D"  images/50cc3d53-9c96-4f8d-a7da-648aea826718.pngPK
   �m�XK숤u  �x  /             �	 images/598b2a10-ddcb-45db-aacd-6c87816d7084.jpgPK
   Jm�Xl� t� /             ^
 images/700d3a7f-db95-4bf3-ad80-33d56978804d.pngPK
   �m�X��
��� � /             �I images/728f499b-3713-4da6-8795-3b437d35f612.pngPK
   �n�Xd��  �   /             �� images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   �n�Xj	hY� {� /             � images/a580090c-3dfd-4391-b47e-11bb84c3f632.pngPK
   �n�X	��#u } /             � images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   �m�X�,͓�u  sx  /             �R images/aced3900-1e1c-42d2-9dab-094da686c0f5.jpgPK
   �n�X�jߩ    /             t� images/d572cae8-d176-4294-a2fa-ef26b385cc14.pngPK
   Jm�XrQ$0 ?4 /             �� images/d821bf6f-d33d-4ee8-8367-12c4d0b7d041.pngPK
   �n�X�{��  B               >	$ jsons/user_defined.jsonPK      $  D$   